VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2223.700 BY 2027.600 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.330 1981.720 1156.610 1984.120 ;
    END
  END address[0]
  PIN address[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1687.630 1981.720 1687.910 1984.120 ;
    END
  END address[10]
  PIN address[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1775.950 1981.720 1776.230 1984.120 ;
    END
  END address[11]
  PIN address[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1682.960 51.880 1683.560 ;
    END
  END address[12]
  PIN address[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.170 44.120 1756.450 46.520 ;
    END
  END address[13]
  PIN address[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1820.570 44.120 1820.850 46.520 ;
    END
  END address[14]
  PIN address[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1702.000 2174.480 1702.600 ;
    END
  END address[15]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1576.880 2174.480 1577.480 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1627.370 44.120 1627.650 46.520 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1244.650 1981.720 1244.930 1984.120 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1691.770 44.120 1692.050 46.520 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1333.430 1981.720 1333.710 1984.120 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1421.750 1981.720 1422.030 1984.120 ;
    END
  END address[6]
  PIN address[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1510.530 1981.720 1510.810 1984.120 ;
    END
  END address[7]
  PIN address[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1639.440 2174.480 1640.040 ;
    END
  END address[8]
  PIN address[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1598.850 1981.720 1599.130 1984.120 ;
    END
  END address[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1764.560 2174.480 1765.160 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1884.970 44.120 1885.250 46.520 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1949.370 44.120 1949.650 46.520 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 93.730 1981.720 94.010 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 447.930 1981.720 448.210 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[10]
  PIN gfpga_pad_GPIO_PAD[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 536.250 1981.720 536.530 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[11]
  PIN gfpga_pad_GPIO_PAD[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 625.030 1981.720 625.310 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[12]
  PIN gfpga_pad_GPIO_PAD[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 713.350 1981.720 713.630 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[13]
  PIN gfpga_pad_GPIO_PAD[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2013.770 44.120 2014.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[14]
  PIN gfpga_pad_GPIO_PAD[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2078.170 44.120 2078.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[15]
  PIN gfpga_pad_GPIO_PAD[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1952.240 2174.480 1952.840 ;
    END
  END gfpga_pad_GPIO_PAD[16]
  PIN gfpga_pad_GPIO_PAD[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1883.560 51.880 1884.160 ;
    END
  END gfpga_pad_GPIO_PAD[17]
  PIN gfpga_pad_GPIO_PAD[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2041.830 1981.720 2042.110 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[18]
  PIN gfpga_pad_GPIO_PAD[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2130.150 1981.720 2130.430 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[19]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 182.050 1981.720 182.330 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 802.130 1981.720 802.410 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[20]
  PIN gfpga_pad_GPIO_PAD[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 890.450 1981.720 890.730 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[21]
  PIN gfpga_pad_GPIO_PAD[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 979.230 1981.720 979.510 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[22]
  PIN gfpga_pad_GPIO_PAD[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1067.550 1981.720 1067.830 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[23]
  PIN gfpga_pad_GPIO_PAD[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 75.440 2174.480 76.040 ;
    END
  END gfpga_pad_GPIO_PAD[24]
  PIN gfpga_pad_GPIO_PAD[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 138.000 2174.480 138.600 ;
    END
  END gfpga_pad_GPIO_PAD[25]
  PIN gfpga_pad_GPIO_PAD[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 200.560 2174.480 201.160 ;
    END
  END gfpga_pad_GPIO_PAD[26]
  PIN gfpga_pad_GPIO_PAD[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 263.120 2174.480 263.720 ;
    END
  END gfpga_pad_GPIO_PAD[27]
  PIN gfpga_pad_GPIO_PAD[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 325.680 2174.480 326.280 ;
    END
  END gfpga_pad_GPIO_PAD[28]
  PIN gfpga_pad_GPIO_PAD[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 388.240 2174.480 388.840 ;
    END
  END gfpga_pad_GPIO_PAD[29]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 270.830 1981.720 271.110 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 450.800 2174.480 451.400 ;
    END
  END gfpga_pad_GPIO_PAD[30]
  PIN gfpga_pad_GPIO_PAD[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 513.360 2174.480 513.960 ;
    END
  END gfpga_pad_GPIO_PAD[31]
  PIN gfpga_pad_GPIO_PAD[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 575.920 2174.480 576.520 ;
    END
  END gfpga_pad_GPIO_PAD[32]
  PIN gfpga_pad_GPIO_PAD[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 638.480 2174.480 639.080 ;
    END
  END gfpga_pad_GPIO_PAD[33]
  PIN gfpga_pad_GPIO_PAD[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 701.040 2174.480 701.640 ;
    END
  END gfpga_pad_GPIO_PAD[34]
  PIN gfpga_pad_GPIO_PAD[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 763.600 2174.480 764.200 ;
    END
  END gfpga_pad_GPIO_PAD[35]
  PIN gfpga_pad_GPIO_PAD[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 826.160 2174.480 826.760 ;
    END
  END gfpga_pad_GPIO_PAD[36]
  PIN gfpga_pad_GPIO_PAD[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 888.720 2174.480 889.320 ;
    END
  END gfpga_pad_GPIO_PAD[37]
  PIN gfpga_pad_GPIO_PAD[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 951.280 2174.480 951.880 ;
    END
  END gfpga_pad_GPIO_PAD[38]
  PIN gfpga_pad_GPIO_PAD[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1013.840 2174.480 1014.440 ;
    END
  END gfpga_pad_GPIO_PAD[39]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 359.150 1981.720 359.430 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1076.400 2174.480 1077.000 ;
    END
  END gfpga_pad_GPIO_PAD[40]
  PIN gfpga_pad_GPIO_PAD[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1138.960 2174.480 1139.560 ;
    END
  END gfpga_pad_GPIO_PAD[41]
  PIN gfpga_pad_GPIO_PAD[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1201.520 2174.480 1202.120 ;
    END
  END gfpga_pad_GPIO_PAD[42]
  PIN gfpga_pad_GPIO_PAD[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1264.080 2174.480 1264.680 ;
    END
  END gfpga_pad_GPIO_PAD[43]
  PIN gfpga_pad_GPIO_PAD[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1326.640 2174.480 1327.240 ;
    END
  END gfpga_pad_GPIO_PAD[44]
  PIN gfpga_pad_GPIO_PAD[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1389.200 2174.480 1389.800 ;
    END
  END gfpga_pad_GPIO_PAD[45]
  PIN gfpga_pad_GPIO_PAD[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1451.760 2174.480 1452.360 ;
    END
  END gfpga_pad_GPIO_PAD[46]
  PIN gfpga_pad_GPIO_PAD[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1514.320 2174.480 1514.920 ;
    END
  END gfpga_pad_GPIO_PAD[47]
  PIN gfpga_pad_GPIO_PAD[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.770 44.120 82.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[48]
  PIN gfpga_pad_GPIO_PAD[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 146.170 44.120 146.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[49]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1864.730 1981.720 1865.010 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 210.570 44.120 210.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[50]
  PIN gfpga_pad_GPIO_PAD[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 274.970 44.120 275.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[51]
  PIN gfpga_pad_GPIO_PAD[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 339.370 44.120 339.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[52]
  PIN gfpga_pad_GPIO_PAD[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 403.770 44.120 404.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[53]
  PIN gfpga_pad_GPIO_PAD[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 468.170 44.120 468.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[54]
  PIN gfpga_pad_GPIO_PAD[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 532.570 44.120 532.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[55]
  PIN gfpga_pad_GPIO_PAD[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 596.970 44.120 597.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[56]
  PIN gfpga_pad_GPIO_PAD[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 661.370 44.120 661.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[57]
  PIN gfpga_pad_GPIO_PAD[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 725.770 44.120 726.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[58]
  PIN gfpga_pad_GPIO_PAD[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 790.170 44.120 790.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[59]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1749.600 51.880 1750.200 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 854.570 44.120 854.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[60]
  PIN gfpga_pad_GPIO_PAD[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 918.970 44.120 919.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[61]
  PIN gfpga_pad_GPIO_PAD[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 983.370 44.120 983.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[62]
  PIN gfpga_pad_GPIO_PAD[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1047.770 44.120 1048.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[63]
  PIN gfpga_pad_GPIO_PAD[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1112.170 44.120 1112.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[64]
  PIN gfpga_pad_GPIO_PAD[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1176.570 44.120 1176.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[65]
  PIN gfpga_pad_GPIO_PAD[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1240.970 44.120 1241.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[66]
  PIN gfpga_pad_GPIO_PAD[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1305.370 44.120 1305.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[67]
  PIN gfpga_pad_GPIO_PAD[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1369.770 44.120 1370.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[68]
  PIN gfpga_pad_GPIO_PAD[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1434.170 44.120 1434.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[69]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1827.120 2174.480 1827.720 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1498.570 44.120 1498.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[70]
  PIN gfpga_pad_GPIO_PAD[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1562.970 44.120 1563.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[71]
  PIN gfpga_pad_GPIO_PAD[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 77.480 51.880 78.080 ;
    END
  END gfpga_pad_GPIO_PAD[72]
  PIN gfpga_pad_GPIO_PAD[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 144.120 51.880 144.720 ;
    END
  END gfpga_pad_GPIO_PAD[73]
  PIN gfpga_pad_GPIO_PAD[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 210.760 51.880 211.360 ;
    END
  END gfpga_pad_GPIO_PAD[74]
  PIN gfpga_pad_GPIO_PAD[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 278.080 51.880 278.680 ;
    END
  END gfpga_pad_GPIO_PAD[75]
  PIN gfpga_pad_GPIO_PAD[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 344.720 51.880 345.320 ;
    END
  END gfpga_pad_GPIO_PAD[76]
  PIN gfpga_pad_GPIO_PAD[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 411.360 51.880 411.960 ;
    END
  END gfpga_pad_GPIO_PAD[77]
  PIN gfpga_pad_GPIO_PAD[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 478.680 51.880 479.280 ;
    END
  END gfpga_pad_GPIO_PAD[78]
  PIN gfpga_pad_GPIO_PAD[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 545.320 51.880 545.920 ;
    END
  END gfpga_pad_GPIO_PAD[79]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1953.050 1981.720 1953.330 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN gfpga_pad_GPIO_PAD[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 612.640 51.880 613.240 ;
    END
  END gfpga_pad_GPIO_PAD[80]
  PIN gfpga_pad_GPIO_PAD[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 679.280 51.880 679.880 ;
    END
  END gfpga_pad_GPIO_PAD[81]
  PIN gfpga_pad_GPIO_PAD[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 745.920 51.880 746.520 ;
    END
  END gfpga_pad_GPIO_PAD[82]
  PIN gfpga_pad_GPIO_PAD[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 813.240 51.880 813.840 ;
    END
  END gfpga_pad_GPIO_PAD[83]
  PIN gfpga_pad_GPIO_PAD[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 879.880 51.880 880.480 ;
    END
  END gfpga_pad_GPIO_PAD[84]
  PIN gfpga_pad_GPIO_PAD[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 946.520 51.880 947.120 ;
    END
  END gfpga_pad_GPIO_PAD[85]
  PIN gfpga_pad_GPIO_PAD[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1013.840 51.880 1014.440 ;
    END
  END gfpga_pad_GPIO_PAD[86]
  PIN gfpga_pad_GPIO_PAD[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1080.480 51.880 1081.080 ;
    END
  END gfpga_pad_GPIO_PAD[87]
  PIN gfpga_pad_GPIO_PAD[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1147.800 51.880 1148.400 ;
    END
  END gfpga_pad_GPIO_PAD[88]
  PIN gfpga_pad_GPIO_PAD[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1214.440 51.880 1215.040 ;
    END
  END gfpga_pad_GPIO_PAD[89]
  PIN gfpga_pad_GPIO_PAD[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1889.680 2174.480 1890.280 ;
    END
  END gfpga_pad_GPIO_PAD[8]
  PIN gfpga_pad_GPIO_PAD[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1281.080 51.880 1281.680 ;
    END
  END gfpga_pad_GPIO_PAD[90]
  PIN gfpga_pad_GPIO_PAD[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1348.400 51.880 1349.000 ;
    END
  END gfpga_pad_GPIO_PAD[91]
  PIN gfpga_pad_GPIO_PAD[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1415.040 51.880 1415.640 ;
    END
  END gfpga_pad_GPIO_PAD[92]
  PIN gfpga_pad_GPIO_PAD[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1481.680 51.880 1482.280 ;
    END
  END gfpga_pad_GPIO_PAD[93]
  PIN gfpga_pad_GPIO_PAD[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1549.000 51.880 1549.600 ;
    END
  END gfpga_pad_GPIO_PAD[94]
  PIN gfpga_pad_GPIO_PAD[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1615.640 51.880 1616.240 ;
    END
  END gfpga_pad_GPIO_PAD[95]
  PIN gfpga_pad_GPIO_PAD[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1816.240 51.880 1816.840 ;
    END
  END gfpga_pad_GPIO_PAD[9]
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1950.200 51.880 1950.800 ;
    END
  END reset
  PIN set
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2142.570 44.120 2142.850 46.520 ;
    END
  END set
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 2198.700 45.000 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 2223.700 20.000 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 105.000 92.485 2118.540 1975.915 ;
      LAYER met1 ;
        RECT 63.350 46.880 2151.610 1975.960 ;
      LAYER met2 ;
        RECT 63.370 1981.440 93.450 1981.720 ;
        RECT 94.290 1981.440 181.770 1981.720 ;
        RECT 182.610 1981.440 270.550 1981.720 ;
        RECT 271.390 1981.440 358.870 1981.720 ;
        RECT 359.710 1981.440 447.650 1981.720 ;
        RECT 448.490 1981.440 535.970 1981.720 ;
        RECT 536.810 1981.440 624.750 1981.720 ;
        RECT 625.590 1981.440 713.070 1981.720 ;
        RECT 713.910 1981.440 801.850 1981.720 ;
        RECT 802.690 1981.440 890.170 1981.720 ;
        RECT 891.010 1981.440 978.950 1981.720 ;
        RECT 979.790 1981.440 1067.270 1981.720 ;
        RECT 1068.110 1981.440 1156.050 1981.720 ;
        RECT 1156.890 1981.440 1244.370 1981.720 ;
        RECT 1245.210 1981.440 1333.150 1981.720 ;
        RECT 1333.990 1981.440 1421.470 1981.720 ;
        RECT 1422.310 1981.440 1510.250 1981.720 ;
        RECT 1511.090 1981.440 1598.570 1981.720 ;
        RECT 1599.410 1981.440 1687.350 1981.720 ;
        RECT 1688.190 1981.440 1775.670 1981.720 ;
        RECT 1776.510 1981.440 1864.450 1981.720 ;
        RECT 1865.290 1981.440 1952.770 1981.720 ;
        RECT 1953.610 1981.440 2041.550 1981.720 ;
        RECT 2042.390 1981.440 2129.870 1981.720 ;
        RECT 2130.710 1981.440 2151.590 1981.720 ;
        RECT 63.370 46.800 2151.590 1981.440 ;
        RECT 63.370 46.520 81.490 46.800 ;
        RECT 82.330 46.520 145.890 46.800 ;
        RECT 146.730 46.520 210.290 46.800 ;
        RECT 211.130 46.520 274.690 46.800 ;
        RECT 275.530 46.520 339.090 46.800 ;
        RECT 339.930 46.520 403.490 46.800 ;
        RECT 404.330 46.520 467.890 46.800 ;
        RECT 468.730 46.520 532.290 46.800 ;
        RECT 533.130 46.520 596.690 46.800 ;
        RECT 597.530 46.520 661.090 46.800 ;
        RECT 661.930 46.520 725.490 46.800 ;
        RECT 726.330 46.520 789.890 46.800 ;
        RECT 790.730 46.520 854.290 46.800 ;
        RECT 855.130 46.520 918.690 46.800 ;
        RECT 919.530 46.520 983.090 46.800 ;
        RECT 983.930 46.520 1047.490 46.800 ;
        RECT 1048.330 46.520 1111.890 46.800 ;
        RECT 1112.730 46.520 1176.290 46.800 ;
        RECT 1177.130 46.520 1240.690 46.800 ;
        RECT 1241.530 46.520 1305.090 46.800 ;
        RECT 1305.930 46.520 1369.490 46.800 ;
        RECT 1370.330 46.520 1433.890 46.800 ;
        RECT 1434.730 46.520 1498.290 46.800 ;
        RECT 1499.130 46.520 1562.690 46.800 ;
        RECT 1563.530 46.520 1627.090 46.800 ;
        RECT 1627.930 46.520 1691.490 46.800 ;
        RECT 1692.330 46.520 1755.890 46.800 ;
        RECT 1756.730 46.520 1820.290 46.800 ;
        RECT 1821.130 46.520 1884.690 46.800 ;
        RECT 1885.530 46.520 1949.090 46.800 ;
        RECT 1949.930 46.520 2013.490 46.800 ;
        RECT 2014.330 46.520 2077.890 46.800 ;
        RECT 2078.730 46.520 2142.290 46.800 ;
        RECT 2143.130 46.520 2151.590 46.800 ;
      LAYER met3 ;
        RECT 51.880 1953.240 2172.080 1969.025 ;
        RECT 51.880 1951.840 2171.680 1953.240 ;
        RECT 51.880 1951.200 2172.080 1951.840 ;
        RECT 52.280 1949.800 2172.080 1951.200 ;
        RECT 51.880 1890.680 2172.080 1949.800 ;
        RECT 51.880 1889.280 2171.680 1890.680 ;
        RECT 51.880 1884.560 2172.080 1889.280 ;
        RECT 52.280 1883.160 2172.080 1884.560 ;
        RECT 51.880 1828.120 2172.080 1883.160 ;
        RECT 51.880 1826.720 2171.680 1828.120 ;
        RECT 51.880 1817.240 2172.080 1826.720 ;
        RECT 52.280 1815.840 2172.080 1817.240 ;
        RECT 51.880 1765.560 2172.080 1815.840 ;
        RECT 51.880 1764.160 2171.680 1765.560 ;
        RECT 51.880 1750.600 2172.080 1764.160 ;
        RECT 52.280 1749.200 2172.080 1750.600 ;
        RECT 51.880 1703.000 2172.080 1749.200 ;
        RECT 51.880 1701.600 2171.680 1703.000 ;
        RECT 51.880 1683.960 2172.080 1701.600 ;
        RECT 52.280 1682.560 2172.080 1683.960 ;
        RECT 51.880 1640.440 2172.080 1682.560 ;
        RECT 51.880 1639.040 2171.680 1640.440 ;
        RECT 51.880 1616.640 2172.080 1639.040 ;
        RECT 52.280 1615.240 2172.080 1616.640 ;
        RECT 51.880 1577.880 2172.080 1615.240 ;
        RECT 51.880 1576.480 2171.680 1577.880 ;
        RECT 51.880 1550.000 2172.080 1576.480 ;
        RECT 52.280 1548.600 2172.080 1550.000 ;
        RECT 51.880 1515.320 2172.080 1548.600 ;
        RECT 51.880 1513.920 2171.680 1515.320 ;
        RECT 51.880 1482.680 2172.080 1513.920 ;
        RECT 52.280 1481.280 2172.080 1482.680 ;
        RECT 51.880 1452.760 2172.080 1481.280 ;
        RECT 51.880 1451.360 2171.680 1452.760 ;
        RECT 51.880 1416.040 2172.080 1451.360 ;
        RECT 52.280 1414.640 2172.080 1416.040 ;
        RECT 51.880 1390.200 2172.080 1414.640 ;
        RECT 51.880 1388.800 2171.680 1390.200 ;
        RECT 51.880 1349.400 2172.080 1388.800 ;
        RECT 52.280 1348.000 2172.080 1349.400 ;
        RECT 51.880 1327.640 2172.080 1348.000 ;
        RECT 51.880 1326.240 2171.680 1327.640 ;
        RECT 51.880 1282.080 2172.080 1326.240 ;
        RECT 52.280 1280.680 2172.080 1282.080 ;
        RECT 51.880 1265.080 2172.080 1280.680 ;
        RECT 51.880 1263.680 2171.680 1265.080 ;
        RECT 51.880 1215.440 2172.080 1263.680 ;
        RECT 52.280 1214.040 2172.080 1215.440 ;
        RECT 51.880 1202.520 2172.080 1214.040 ;
        RECT 51.880 1201.120 2171.680 1202.520 ;
        RECT 51.880 1148.800 2172.080 1201.120 ;
        RECT 52.280 1147.400 2172.080 1148.800 ;
        RECT 51.880 1139.960 2172.080 1147.400 ;
        RECT 51.880 1138.560 2171.680 1139.960 ;
        RECT 51.880 1081.480 2172.080 1138.560 ;
        RECT 52.280 1080.080 2172.080 1081.480 ;
        RECT 51.880 1077.400 2172.080 1080.080 ;
        RECT 51.880 1076.000 2171.680 1077.400 ;
        RECT 51.880 1014.840 2172.080 1076.000 ;
        RECT 52.280 1013.440 2171.680 1014.840 ;
        RECT 51.880 952.280 2172.080 1013.440 ;
        RECT 51.880 950.880 2171.680 952.280 ;
        RECT 51.880 947.520 2172.080 950.880 ;
        RECT 52.280 946.120 2172.080 947.520 ;
        RECT 51.880 889.720 2172.080 946.120 ;
        RECT 51.880 888.320 2171.680 889.720 ;
        RECT 51.880 880.880 2172.080 888.320 ;
        RECT 52.280 879.480 2172.080 880.880 ;
        RECT 51.880 827.160 2172.080 879.480 ;
        RECT 51.880 825.760 2171.680 827.160 ;
        RECT 51.880 814.240 2172.080 825.760 ;
        RECT 52.280 812.840 2172.080 814.240 ;
        RECT 51.880 764.600 2172.080 812.840 ;
        RECT 51.880 763.200 2171.680 764.600 ;
        RECT 51.880 746.920 2172.080 763.200 ;
        RECT 52.280 745.520 2172.080 746.920 ;
        RECT 51.880 702.040 2172.080 745.520 ;
        RECT 51.880 700.640 2171.680 702.040 ;
        RECT 51.880 680.280 2172.080 700.640 ;
        RECT 52.280 678.880 2172.080 680.280 ;
        RECT 51.880 639.480 2172.080 678.880 ;
        RECT 51.880 638.080 2171.680 639.480 ;
        RECT 51.880 613.640 2172.080 638.080 ;
        RECT 52.280 612.240 2172.080 613.640 ;
        RECT 51.880 576.920 2172.080 612.240 ;
        RECT 51.880 575.520 2171.680 576.920 ;
        RECT 51.880 546.320 2172.080 575.520 ;
        RECT 52.280 544.920 2172.080 546.320 ;
        RECT 51.880 514.360 2172.080 544.920 ;
        RECT 51.880 512.960 2171.680 514.360 ;
        RECT 51.880 479.680 2172.080 512.960 ;
        RECT 52.280 478.280 2172.080 479.680 ;
        RECT 51.880 451.800 2172.080 478.280 ;
        RECT 51.880 450.400 2171.680 451.800 ;
        RECT 51.880 412.360 2172.080 450.400 ;
        RECT 52.280 410.960 2172.080 412.360 ;
        RECT 51.880 389.240 2172.080 410.960 ;
        RECT 51.880 387.840 2171.680 389.240 ;
        RECT 51.880 345.720 2172.080 387.840 ;
        RECT 52.280 344.320 2172.080 345.720 ;
        RECT 51.880 326.680 2172.080 344.320 ;
        RECT 51.880 325.280 2171.680 326.680 ;
        RECT 51.880 279.080 2172.080 325.280 ;
        RECT 52.280 277.680 2172.080 279.080 ;
        RECT 51.880 264.120 2172.080 277.680 ;
        RECT 51.880 262.720 2171.680 264.120 ;
        RECT 51.880 211.760 2172.080 262.720 ;
        RECT 52.280 210.360 2172.080 211.760 ;
        RECT 51.880 201.560 2172.080 210.360 ;
        RECT 51.880 200.160 2171.680 201.560 ;
        RECT 51.880 145.120 2172.080 200.160 ;
        RECT 52.280 143.720 2172.080 145.120 ;
        RECT 51.880 139.000 2172.080 143.720 ;
        RECT 51.880 137.600 2171.680 139.000 ;
        RECT 51.880 78.480 2172.080 137.600 ;
        RECT 52.280 77.080 2172.080 78.480 ;
        RECT 51.880 76.440 2172.080 77.080 ;
        RECT 51.880 75.575 2171.680 76.440 ;
      LAYER met4 ;
        RECT 0.000 0.000 2223.700 2027.600 ;
      LAYER met5 ;
        RECT 0.000 119.200 2223.700 2027.600 ;
  END
END fpga_top
END LIBRARY

