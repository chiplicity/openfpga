magic
tech EFS8A
magscale 1 2
timestamp 1604344731
<< locali >>
rect 24501 3995 24535 4233
rect 20085 3383 20119 3485
rect 23305 2839 23339 2941
<< viali >>
rect 15485 23817 15519 23851
rect 25145 23817 25179 23851
rect 14841 23613 14875 23647
rect 24593 23613 24627 23647
rect 15025 23477 15059 23511
rect 24777 23477 24811 23511
rect 16129 22049 16163 22083
rect 16313 21845 16347 21879
rect 16129 21641 16163 21675
rect 17509 20961 17543 20995
rect 17693 20757 17727 20791
rect 17509 20553 17543 20587
rect 24593 19873 24627 19907
rect 24777 19669 24811 19703
rect 24593 19465 24627 19499
rect 18889 19261 18923 19295
rect 19533 19193 19567 19227
rect 19073 19125 19107 19159
rect 19625 18785 19659 18819
rect 19809 18581 19843 18615
rect 19717 18377 19751 18411
rect 20913 18377 20947 18411
rect 20269 18173 20303 18207
rect 20453 18037 20487 18071
rect 20913 17697 20947 17731
rect 21097 17493 21131 17527
rect 21005 17289 21039 17323
rect 21833 16745 21867 16779
rect 21649 16609 21683 16643
rect 21649 16201 21683 16235
rect 23213 15521 23247 15555
rect 23397 15317 23431 15351
rect 23305 15113 23339 15147
rect 24501 15113 24535 15147
rect 23857 14909 23891 14943
rect 24041 14773 24075 14807
rect 25237 14025 25271 14059
rect 24777 13957 24811 13991
rect 24593 13821 24627 13855
rect 24593 13345 24627 13379
rect 24777 13141 24811 13175
rect 24501 12937 24535 12971
rect 25237 12937 25271 12971
rect 24777 12869 24811 12903
rect 24593 12733 24627 12767
rect 24593 12257 24627 12291
rect 24777 12053 24811 12087
rect 13829 11849 13863 11883
rect 24685 11849 24719 11883
rect 13645 11645 13679 11679
rect 14197 11509 14231 11543
rect 20361 11033 20395 11067
rect 20085 10693 20119 10727
rect 20361 10693 20395 10727
rect 20913 10625 20947 10659
rect 1409 10557 1443 10591
rect 1961 10557 1995 10591
rect 20637 10489 20671 10523
rect 20821 10489 20855 10523
rect 1593 10421 1627 10455
rect 19809 10217 19843 10251
rect 20361 10217 20395 10251
rect 22293 10217 22327 10251
rect 1409 10081 1443 10115
rect 20913 10081 20947 10115
rect 21180 10081 21214 10115
rect 1593 9945 1627 9979
rect 21833 9673 21867 9707
rect 2053 9469 2087 9503
rect 19809 9469 19843 9503
rect 19901 9469 19935 9503
rect 20146 9401 20180 9435
rect 22201 9401 22235 9435
rect 1593 9333 1627 9367
rect 2237 9333 2271 9367
rect 2605 9333 2639 9367
rect 18797 9333 18831 9367
rect 19441 9333 19475 9367
rect 21281 9333 21315 9367
rect 19809 9129 19843 9163
rect 21465 9129 21499 9163
rect 2697 8993 2731 9027
rect 19625 8993 19659 9027
rect 21281 8993 21315 9027
rect 22477 8993 22511 9027
rect 19901 8925 19935 8959
rect 21557 8925 21591 8959
rect 22661 8925 22695 8959
rect 2881 8857 2915 8891
rect 21005 8857 21039 8891
rect 19349 8789 19383 8823
rect 18889 8585 18923 8619
rect 20729 8585 20763 8619
rect 21649 8585 21683 8619
rect 22477 8585 22511 8619
rect 19349 8449 19383 8483
rect 19165 8381 19199 8415
rect 2789 8313 2823 8347
rect 18521 8313 18555 8347
rect 19594 8313 19628 8347
rect 21281 8313 21315 8347
rect 19257 8041 19291 8075
rect 20085 8041 20119 8075
rect 21189 8041 21223 8075
rect 19073 7973 19107 8007
rect 17417 7905 17451 7939
rect 17601 7837 17635 7871
rect 19349 7837 19383 7871
rect 18797 7769 18831 7803
rect 19717 7701 19751 7735
rect 17509 7497 17543 7531
rect 17877 7497 17911 7531
rect 18337 7497 18371 7531
rect 18705 7497 18739 7531
rect 20545 7497 20579 7531
rect 4077 7293 4111 7327
rect 19165 7293 19199 7327
rect 19432 7225 19466 7259
rect 4261 7157 4295 7191
rect 4629 7157 4663 7191
rect 19073 7157 19107 7191
rect 19809 6953 19843 6987
rect 24777 6953 24811 6987
rect 18245 6885 18279 6919
rect 21465 6885 21499 6919
rect 16589 6817 16623 6851
rect 18061 6817 18095 6851
rect 19625 6817 19659 6851
rect 21281 6817 21315 6851
rect 24593 6817 24627 6851
rect 18337 6749 18371 6783
rect 18797 6749 18831 6783
rect 19901 6749 19935 6783
rect 21557 6749 21591 6783
rect 23121 6749 23155 6783
rect 19349 6681 19383 6715
rect 16773 6613 16807 6647
rect 17785 6613 17819 6647
rect 19073 6613 19107 6647
rect 21005 6613 21039 6647
rect 16681 6409 16715 6443
rect 17417 6409 17451 6443
rect 18613 6409 18647 6443
rect 20453 6409 20487 6443
rect 21465 6409 21499 6443
rect 24685 6409 24719 6443
rect 17785 6273 17819 6307
rect 18061 6273 18095 6307
rect 23949 6273 23983 6307
rect 19073 6205 19107 6239
rect 23489 6205 23523 6239
rect 23673 6205 23707 6239
rect 24961 6205 24995 6239
rect 25513 6205 25547 6239
rect 19340 6137 19374 6171
rect 18889 6069 18923 6103
rect 21005 6069 21039 6103
rect 21741 6069 21775 6103
rect 25145 6069 25179 6103
rect 17785 5865 17819 5899
rect 18245 5865 18279 5899
rect 23581 5865 23615 5899
rect 22446 5797 22480 5831
rect 24961 5797 24995 5831
rect 16957 5729 16991 5763
rect 18604 5729 18638 5763
rect 22201 5729 22235 5763
rect 24685 5729 24719 5763
rect 17141 5661 17175 5695
rect 18337 5661 18371 5695
rect 20913 5661 20947 5695
rect 19717 5525 19751 5559
rect 20361 5525 20395 5559
rect 24133 5525 24167 5559
rect 16589 5321 16623 5355
rect 17049 5321 17083 5355
rect 18705 5321 18739 5355
rect 19533 5321 19567 5355
rect 21005 5321 21039 5355
rect 22201 5321 22235 5355
rect 23489 5321 23523 5355
rect 23765 5321 23799 5355
rect 18429 5253 18463 5287
rect 19625 5185 19659 5219
rect 24133 5185 24167 5219
rect 15945 5117 15979 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 19870 5049 19904 5083
rect 21925 5049 21959 5083
rect 23121 5049 23155 5083
rect 24317 5049 24351 5083
rect 16129 4981 16163 5015
rect 19165 4981 19199 5015
rect 22569 4981 22603 5015
rect 24225 4981 24259 5015
rect 24685 4981 24719 5015
rect 25421 4981 25455 5015
rect 18245 4777 18279 4811
rect 19165 4777 19199 4811
rect 19809 4777 19843 4811
rect 22385 4777 22419 4811
rect 24685 4777 24719 4811
rect 6837 4641 6871 4675
rect 15301 4641 15335 4675
rect 19625 4641 19659 4675
rect 22201 4641 22235 4675
rect 23572 4641 23606 4675
rect 15485 4573 15519 4607
rect 19901 4573 19935 4607
rect 20913 4573 20947 4607
rect 23305 4573 23339 4607
rect 7021 4505 7055 4539
rect 19349 4505 19383 4539
rect 22109 4505 22143 4539
rect 21373 4437 21407 4471
rect 22845 4437 22879 4471
rect 7665 4233 7699 4267
rect 15301 4233 15335 4267
rect 20177 4233 20211 4267
rect 20821 4233 20855 4267
rect 23765 4233 23799 4267
rect 24501 4233 24535 4267
rect 24777 4233 24811 4267
rect 14841 4097 14875 4131
rect 17877 4097 17911 4131
rect 20637 4097 20671 4131
rect 21189 4097 21223 4131
rect 22569 4097 22603 4131
rect 7481 4029 7515 4063
rect 8033 4029 8067 4063
rect 14197 4029 14231 4063
rect 18153 4029 18187 4063
rect 18409 4029 18443 4063
rect 22293 4029 22327 4063
rect 24317 4029 24351 4063
rect 25421 4097 25455 4131
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 25973 4029 26007 4063
rect 21373 3961 21407 3995
rect 23489 3961 23523 3995
rect 24041 3961 24075 3995
rect 24225 3961 24259 3995
rect 24501 3961 24535 3995
rect 7113 3893 7147 3927
rect 14381 3893 14415 3927
rect 19533 3893 19567 3927
rect 21281 3893 21315 3927
rect 21833 3893 21867 3927
rect 22109 3893 22143 3927
rect 23121 3893 23155 3927
rect 18797 3689 18831 3723
rect 19165 3689 19199 3723
rect 23397 3689 23431 3723
rect 24869 3689 24903 3723
rect 18245 3621 18279 3655
rect 18337 3621 18371 3655
rect 19809 3621 19843 3655
rect 8125 3553 8159 3587
rect 18061 3553 18095 3587
rect 19625 3553 19659 3587
rect 21180 3553 21214 3587
rect 22937 3553 22971 3587
rect 23756 3553 23790 3587
rect 19901 3485 19935 3519
rect 20085 3485 20119 3519
rect 20913 3485 20947 3519
rect 23489 3485 23523 3519
rect 8309 3417 8343 3451
rect 19349 3417 19383 3451
rect 16497 3349 16531 3383
rect 17785 3349 17819 3383
rect 20085 3349 20119 3383
rect 20361 3349 20395 3383
rect 20729 3349 20763 3383
rect 22293 3349 22327 3383
rect 16497 3145 16531 3179
rect 18521 3145 18555 3179
rect 20913 3145 20947 3179
rect 22109 3145 22143 3179
rect 18797 3077 18831 3111
rect 18981 3009 19015 3043
rect 21925 3009 21959 3043
rect 22477 3009 22511 3043
rect 8861 2941 8895 2975
rect 9413 2941 9447 2975
rect 17049 2941 17083 2975
rect 23305 2941 23339 2975
rect 23673 2941 23707 2975
rect 16313 2873 16347 2907
rect 16773 2873 16807 2907
rect 16957 2873 16991 2907
rect 19226 2873 19260 2907
rect 22569 2873 22603 2907
rect 22661 2873 22695 2907
rect 23940 2873 23974 2907
rect 25605 2873 25639 2907
rect 8217 2805 8251 2839
rect 9045 2805 9079 2839
rect 17693 2805 17727 2839
rect 20361 2805 20395 2839
rect 21281 2805 21315 2839
rect 23121 2805 23155 2839
rect 23305 2805 23339 2839
rect 23489 2805 23523 2839
rect 25053 2805 25087 2839
rect 11069 2601 11103 2635
rect 16497 2601 16531 2635
rect 17233 2601 17267 2635
rect 17785 2601 17819 2635
rect 18981 2601 19015 2635
rect 20913 2601 20947 2635
rect 22569 2601 22603 2635
rect 23857 2601 23891 2635
rect 18153 2533 18187 2567
rect 20085 2533 20119 2567
rect 20545 2533 20579 2567
rect 21456 2533 21490 2567
rect 24286 2533 24320 2567
rect 25973 2533 26007 2567
rect 4077 2465 4111 2499
rect 4629 2465 4663 2499
rect 5457 2465 5491 2499
rect 6929 2465 6963 2499
rect 7481 2465 7515 2499
rect 9781 2465 9815 2499
rect 10333 2465 10367 2499
rect 10885 2465 10919 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 18429 2465 18463 2499
rect 20177 2465 20211 2499
rect 21189 2465 21223 2499
rect 24041 2465 24075 2499
rect 17141 2397 17175 2431
rect 19993 2397 20027 2431
rect 5641 2329 5675 2363
rect 19625 2329 19659 2363
rect 4261 2261 4295 2295
rect 6009 2261 6043 2295
rect 7113 2261 7147 2295
rect 9965 2261 9999 2295
rect 11437 2261 11471 2295
rect 12817 2261 12851 2295
rect 16129 2261 16163 2295
rect 18613 2261 18647 2295
rect 19441 2261 19475 2295
rect 23489 2261 23523 2295
rect 25421 2261 25455 2295
<< metal1 >>
rect 20898 26664 20904 26716
rect 20956 26704 20962 26716
rect 24118 26704 24124 26716
rect 20956 26676 24124 26704
rect 20956 26664 20962 26676
rect 24118 26664 24124 26676
rect 24176 26664 24182 26716
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 21726 24896 21732 24948
rect 21784 24936 21790 24948
rect 23750 24936 23756 24948
rect 21784 24908 23756 24936
rect 21784 24896 21790 24908
rect 23750 24896 23756 24908
rect 23808 24896 23814 24948
rect 15470 24828 15476 24880
rect 15528 24868 15534 24880
rect 24762 24868 24768 24880
rect 15528 24840 24768 24868
rect 15528 24828 15534 24840
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 15470 23848 15476 23860
rect 15431 23820 15476 23848
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 24670 23808 24676 23860
rect 24728 23848 24734 23860
rect 25133 23851 25191 23857
rect 25133 23848 25145 23851
rect 24728 23820 25145 23848
rect 24728 23808 24734 23820
rect 25133 23817 25145 23820
rect 25179 23817 25191 23851
rect 25133 23811 25191 23817
rect 14829 23647 14887 23653
rect 14829 23613 14841 23647
rect 14875 23644 14887 23647
rect 15470 23644 15476 23656
rect 14875 23616 15476 23644
rect 14875 23613 14887 23616
rect 14829 23607 14887 23613
rect 15470 23604 15476 23616
rect 15528 23604 15534 23656
rect 24581 23647 24639 23653
rect 24581 23613 24593 23647
rect 24627 23644 24639 23647
rect 24670 23644 24676 23656
rect 24627 23616 24676 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 24670 23604 24676 23616
rect 24728 23604 24734 23656
rect 14826 23468 14832 23520
rect 14884 23508 14890 23520
rect 15013 23511 15071 23517
rect 15013 23508 15025 23511
rect 14884 23480 15025 23508
rect 14884 23468 14890 23480
rect 15013 23477 15025 23480
rect 15059 23477 15071 23511
rect 15013 23471 15071 23477
rect 23658 23468 23664 23520
rect 23716 23508 23722 23520
rect 24765 23511 24823 23517
rect 24765 23508 24777 23511
rect 23716 23480 24777 23508
rect 23716 23468 23722 23480
rect 24765 23477 24777 23480
rect 24811 23477 24823 23511
rect 24765 23471 24823 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 16114 22080 16120 22092
rect 16075 22052 16120 22080
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 16298 21876 16304 21888
rect 16259 21848 16304 21876
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 16114 21672 16120 21684
rect 16075 21644 16120 21672
rect 16114 21632 16120 21644
rect 16172 21632 16178 21684
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 23566 21088 23572 21140
rect 23624 21128 23630 21140
rect 23934 21128 23940 21140
rect 23624 21100 23940 21128
rect 23624 21088 23630 21100
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 17494 20992 17500 21004
rect 17455 20964 17500 20992
rect 17494 20952 17500 20964
rect 17552 20952 17558 21004
rect 17678 20788 17684 20800
rect 17639 20760 17684 20788
rect 17678 20748 17684 20760
rect 17736 20748 17742 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 17494 20584 17500 20596
rect 17455 20556 17500 20584
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 24026 19864 24032 19916
rect 24084 19904 24090 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 24084 19876 24593 19904
rect 24084 19864 24090 19876
rect 24581 19873 24593 19876
rect 24627 19904 24639 19907
rect 24670 19904 24676 19916
rect 24627 19876 24676 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 24762 19700 24768 19712
rect 24723 19672 24768 19700
rect 24762 19660 24768 19672
rect 24820 19660 24826 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24581 19499 24639 19505
rect 24581 19496 24593 19499
rect 24084 19468 24593 19496
rect 24084 19456 24090 19468
rect 24581 19465 24593 19468
rect 24627 19465 24639 19499
rect 24581 19459 24639 19465
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 16298 19292 16304 19304
rect 16172 19264 16304 19292
rect 16172 19252 16178 19264
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 18892 19224 18920 19255
rect 19518 19224 19524 19236
rect 18892 19196 19524 19224
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 19061 19159 19119 19165
rect 19061 19156 19073 19159
rect 19024 19128 19073 19156
rect 19024 19116 19030 19128
rect 19061 19125 19073 19128
rect 19107 19125 19119 19159
rect 19061 19119 19119 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 19613 18819 19671 18825
rect 19613 18785 19625 18819
rect 19659 18816 19671 18819
rect 19978 18816 19984 18828
rect 19659 18788 19984 18816
rect 19659 18785 19671 18788
rect 19613 18779 19671 18785
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 19797 18615 19855 18621
rect 19797 18581 19809 18615
rect 19843 18612 19855 18615
rect 20070 18612 20076 18624
rect 19843 18584 20076 18612
rect 19843 18581 19855 18584
rect 19797 18575 19855 18581
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 19705 18411 19763 18417
rect 19705 18377 19717 18411
rect 19751 18408 19763 18411
rect 19978 18408 19984 18420
rect 19751 18380 19984 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20898 18408 20904 18420
rect 20859 18380 20904 18408
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 20257 18207 20315 18213
rect 20257 18173 20269 18207
rect 20303 18204 20315 18207
rect 20898 18204 20904 18216
rect 20303 18176 20904 18204
rect 20303 18173 20315 18176
rect 20257 18167 20315 18173
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 20438 18068 20444 18080
rect 20399 18040 20444 18068
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 20990 17728 20996 17740
rect 20947 17700 20996 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 20990 17688 20996 17700
rect 21048 17688 21054 17740
rect 21085 17527 21143 17533
rect 21085 17493 21097 17527
rect 21131 17524 21143 17527
rect 21174 17524 21180 17536
rect 21131 17496 21180 17524
rect 21131 17493 21143 17496
rect 21085 17487 21143 17493
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 20990 17320 20996 17332
rect 20951 17292 20996 17320
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 21821 16779 21879 16785
rect 21821 16745 21833 16779
rect 21867 16776 21879 16779
rect 21910 16776 21916 16788
rect 21867 16748 21916 16776
rect 21867 16745 21879 16748
rect 21821 16739 21879 16745
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 21634 16640 21640 16652
rect 21595 16612 21640 16640
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 21634 16232 21640 16244
rect 21595 16204 21640 16232
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 23201 15555 23259 15561
rect 23201 15521 23213 15555
rect 23247 15552 23259 15555
rect 23382 15552 23388 15564
rect 23247 15524 23388 15552
rect 23247 15521 23259 15524
rect 23201 15515 23259 15521
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 23382 15348 23388 15360
rect 23343 15320 23388 15348
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 23290 15144 23296 15156
rect 23251 15116 23296 15144
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 24489 15147 24547 15153
rect 24489 15113 24501 15147
rect 24535 15144 24547 15147
rect 24762 15144 24768 15156
rect 24535 15116 24768 15144
rect 24535 15113 24547 15116
rect 24489 15107 24547 15113
rect 23845 14943 23903 14949
rect 23845 14909 23857 14943
rect 23891 14940 23903 14943
rect 24504 14940 24532 15107
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 23891 14912 24532 14940
rect 23891 14909 23903 14912
rect 23845 14903 23903 14909
rect 24026 14804 24032 14816
rect 23987 14776 24032 14804
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 25222 14056 25228 14068
rect 25183 14028 25228 14056
rect 25222 14016 25228 14028
rect 25280 14016 25286 14068
rect 23842 13948 23848 14000
rect 23900 13988 23906 14000
rect 24765 13991 24823 13997
rect 24765 13988 24777 13991
rect 23900 13960 24777 13988
rect 23900 13948 23906 13960
rect 24765 13957 24777 13960
rect 24811 13957 24823 13991
rect 24765 13951 24823 13957
rect 24581 13855 24639 13861
rect 24581 13821 24593 13855
rect 24627 13852 24639 13855
rect 25222 13852 25228 13864
rect 24627 13824 25228 13852
rect 24627 13821 24639 13824
rect 24581 13815 24639 13821
rect 25222 13812 25228 13824
rect 25280 13812 25286 13864
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 24581 13379 24639 13385
rect 24581 13345 24593 13379
rect 24627 13376 24639 13379
rect 24854 13376 24860 13388
rect 24627 13348 24860 13376
rect 24627 13345 24639 13348
rect 24581 13339 24639 13345
rect 24854 13336 24860 13348
rect 24912 13336 24918 13388
rect 24210 13200 24216 13252
rect 24268 13240 24274 13252
rect 25038 13240 25044 13252
rect 24268 13212 25044 13240
rect 24268 13200 24274 13212
rect 25038 13200 25044 13212
rect 25096 13200 25102 13252
rect 24670 13132 24676 13184
rect 24728 13172 24734 13184
rect 24765 13175 24823 13181
rect 24765 13172 24777 13175
rect 24728 13144 24777 13172
rect 24728 13132 24734 13144
rect 24765 13141 24777 13144
rect 24811 13141 24823 13175
rect 24765 13135 24823 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 24489 12971 24547 12977
rect 24489 12937 24501 12971
rect 24535 12968 24547 12971
rect 24854 12968 24860 12980
rect 24535 12940 24860 12968
rect 24535 12937 24547 12940
rect 24489 12931 24547 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 25225 12971 25283 12977
rect 25225 12937 25237 12971
rect 25271 12968 25283 12971
rect 25314 12968 25320 12980
rect 25271 12940 25320 12968
rect 25271 12937 25283 12940
rect 25225 12931 25283 12937
rect 23934 12860 23940 12912
rect 23992 12900 23998 12912
rect 24765 12903 24823 12909
rect 24765 12900 24777 12903
rect 23992 12872 24777 12900
rect 23992 12860 23998 12872
rect 24765 12869 24777 12872
rect 24811 12869 24823 12903
rect 24765 12863 24823 12869
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 25240 12764 25268 12931
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 24627 12736 25268 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 24578 12588 24584 12640
rect 24636 12628 24642 12640
rect 24762 12628 24768 12640
rect 24636 12600 24768 12628
rect 24636 12588 24642 12600
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 23658 12424 23664 12436
rect 23532 12396 23664 12424
rect 23532 12384 23538 12396
rect 23658 12384 23664 12396
rect 23716 12384 23722 12436
rect 23750 12384 23756 12436
rect 23808 12424 23814 12436
rect 23934 12424 23940 12436
rect 23808 12396 23940 12424
rect 23808 12384 23814 12396
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 24026 12384 24032 12436
rect 24084 12384 24090 12436
rect 24670 12424 24676 12436
rect 24136 12396 24676 12424
rect 24044 12232 24072 12384
rect 24136 12232 24164 12396
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 24581 12291 24639 12297
rect 24581 12257 24593 12291
rect 24627 12288 24639 12291
rect 24670 12288 24676 12300
rect 24627 12260 24676 12288
rect 24627 12257 24639 12260
rect 24581 12251 24639 12257
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 24026 12180 24032 12232
rect 24084 12180 24090 12232
rect 24118 12180 24124 12232
rect 24176 12180 24182 12232
rect 24762 12084 24768 12096
rect 24723 12056 24768 12084
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 13633 11679 13691 11685
rect 13633 11645 13645 11679
rect 13679 11676 13691 11679
rect 13679 11648 14228 11676
rect 13679 11645 13691 11648
rect 13633 11639 13691 11645
rect 14200 11552 14228 11648
rect 14182 11540 14188 11552
rect 14143 11512 14188 11540
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 20349 11067 20407 11073
rect 20349 11033 20361 11067
rect 20395 11064 20407 11067
rect 20714 11064 20720 11076
rect 20395 11036 20720 11064
rect 20395 11033 20407 11036
rect 20349 11027 20407 11033
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 19978 10684 19984 10736
rect 20036 10724 20042 10736
rect 20073 10727 20131 10733
rect 20073 10724 20085 10727
rect 20036 10696 20085 10724
rect 20036 10684 20042 10696
rect 20073 10693 20085 10696
rect 20119 10693 20131 10727
rect 20346 10724 20352 10736
rect 20307 10696 20352 10724
rect 20073 10687 20131 10693
rect 20088 10656 20116 10687
rect 20346 10684 20352 10696
rect 20404 10684 20410 10736
rect 20901 10659 20959 10665
rect 20901 10656 20913 10659
rect 20088 10628 20913 10656
rect 20901 10625 20913 10628
rect 20947 10656 20959 10659
rect 22278 10656 22284 10668
rect 20947 10628 22284 10656
rect 20947 10625 20959 10628
rect 20901 10619 20959 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1670 10588 1676 10600
rect 1443 10560 1676 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1670 10548 1676 10560
rect 1728 10588 1734 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1728 10560 1961 10588
rect 1728 10548 1734 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 20622 10520 20628 10532
rect 20583 10492 20628 10520
rect 20622 10480 20628 10492
rect 20680 10480 20686 10532
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 20809 10523 20867 10529
rect 20809 10520 20821 10523
rect 20772 10492 20821 10520
rect 20772 10480 20778 10492
rect 20809 10489 20821 10492
rect 20855 10489 20867 10523
rect 20809 10483 20867 10489
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 19797 10251 19855 10257
rect 19797 10217 19809 10251
rect 19843 10248 19855 10251
rect 20349 10251 20407 10257
rect 20349 10248 20361 10251
rect 19843 10220 20361 10248
rect 19843 10217 19855 10220
rect 19797 10211 19855 10217
rect 20349 10217 20361 10220
rect 20395 10248 20407 10251
rect 20622 10248 20628 10260
rect 20395 10220 20628 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 22278 10248 22284 10260
rect 22239 10220 22284 10248
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1486 10112 1492 10124
rect 1443 10084 1492 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20864 10084 20913 10112
rect 20864 10072 20870 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 21168 10115 21226 10121
rect 21168 10081 21180 10115
rect 21214 10112 21226 10115
rect 21542 10112 21548 10124
rect 21214 10084 21548 10112
rect 21214 10081 21226 10084
rect 21168 10075 21226 10081
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 1578 9976 1584 9988
rect 1539 9948 1584 9976
rect 1578 9936 1584 9948
rect 1636 9936 1642 9988
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 16206 9704 16212 9716
rect 16172 9676 16212 9704
rect 16172 9664 16178 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 21818 9704 21824 9716
rect 20864 9676 21824 9704
rect 20864 9664 20870 9676
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9500 2099 9503
rect 19797 9503 19855 9509
rect 2087 9472 2360 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 2332 9376 2360 9472
rect 19797 9469 19809 9503
rect 19843 9500 19855 9503
rect 19889 9503 19947 9509
rect 19889 9500 19901 9503
rect 19843 9472 19901 9500
rect 19843 9469 19855 9472
rect 19797 9463 19855 9469
rect 19889 9469 19901 9472
rect 19935 9500 19947 9503
rect 20916 9500 20944 9676
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 19935 9472 20944 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 20134 9435 20192 9441
rect 20134 9432 20146 9435
rect 19444 9404 20146 9432
rect 19444 9376 19472 9404
rect 20134 9401 20146 9404
rect 20180 9401 20192 9435
rect 22189 9435 22247 9441
rect 22189 9432 22201 9435
rect 20134 9395 20192 9401
rect 21560 9404 22201 9432
rect 21560 9376 21588 9404
rect 22189 9401 22201 9404
rect 22235 9401 22247 9435
rect 22189 9395 22247 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2314 9324 2320 9376
rect 2372 9364 2378 9376
rect 2593 9367 2651 9373
rect 2593 9364 2605 9367
rect 2372 9336 2605 9364
rect 2372 9324 2378 9336
rect 2593 9333 2605 9336
rect 2639 9333 2651 9367
rect 18782 9364 18788 9376
rect 18743 9336 18788 9364
rect 2593 9327 2651 9333
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 21269 9367 21327 9373
rect 21269 9333 21281 9367
rect 21315 9364 21327 9367
rect 21542 9364 21548 9376
rect 21315 9336 21548 9364
rect 21315 9333 21327 9336
rect 21269 9327 21327 9333
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 18874 9120 18880 9172
rect 18932 9160 18938 9172
rect 19797 9163 19855 9169
rect 19797 9160 19809 9163
rect 18932 9132 19809 9160
rect 18932 9120 18938 9132
rect 19797 9129 19809 9132
rect 19843 9160 19855 9163
rect 20162 9160 20168 9172
rect 19843 9132 20168 9160
rect 19843 9129 19855 9132
rect 19797 9123 19855 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 21450 9160 21456 9172
rect 21411 9132 21456 9160
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 2958 9024 2964 9036
rect 2731 8996 2964 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19300 8996 19625 9024
rect 19300 8984 19306 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 21266 9024 21272 9036
rect 21227 8996 21272 9024
rect 19613 8987 19671 8993
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 22462 9024 22468 9036
rect 22423 8996 22468 9024
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 19886 8956 19892 8968
rect 19847 8928 19892 8956
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 21542 8956 21548 8968
rect 21503 8928 21548 8956
rect 21542 8916 21548 8928
rect 21600 8916 21606 8968
rect 22646 8956 22652 8968
rect 22607 8928 22652 8956
rect 22646 8916 22652 8928
rect 22704 8916 22710 8968
rect 2866 8888 2872 8900
rect 2827 8860 2872 8888
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 20714 8848 20720 8900
rect 20772 8888 20778 8900
rect 20993 8891 21051 8897
rect 20993 8888 21005 8891
rect 20772 8860 21005 8888
rect 20772 8848 20778 8860
rect 20993 8857 21005 8860
rect 21039 8857 21051 8891
rect 20993 8851 21051 8857
rect 19334 8820 19340 8832
rect 19295 8792 19340 8820
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 18874 8616 18880 8628
rect 18835 8588 18880 8616
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 19518 8576 19524 8628
rect 19576 8616 19582 8628
rect 20717 8619 20775 8625
rect 20717 8616 20729 8619
rect 19576 8588 20729 8616
rect 19576 8576 19582 8588
rect 20717 8585 20729 8588
rect 20763 8585 20775 8619
rect 20717 8579 20775 8585
rect 21450 8576 21456 8628
rect 21508 8616 21514 8628
rect 21637 8619 21695 8625
rect 21637 8616 21649 8619
rect 21508 8588 21649 8616
rect 21508 8576 21514 8588
rect 21637 8585 21649 8588
rect 21683 8585 21695 8619
rect 22462 8616 22468 8628
rect 22423 8588 22468 8616
rect 21637 8579 21695 8585
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 19058 8440 19064 8492
rect 19116 8480 19122 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19116 8452 19349 8480
rect 19116 8440 19122 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 18874 8372 18880 8424
rect 18932 8412 18938 8424
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18932 8384 19165 8412
rect 18932 8372 18938 8384
rect 19153 8381 19165 8384
rect 19199 8412 19211 8415
rect 19242 8412 19248 8424
rect 19199 8384 19248 8412
rect 19199 8381 19211 8384
rect 19153 8375 19211 8381
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 2958 8344 2964 8356
rect 2823 8316 2964 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 19582 8347 19640 8353
rect 19582 8344 19594 8347
rect 18555 8316 19594 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 19582 8313 19594 8316
rect 19628 8344 19640 8347
rect 19886 8344 19892 8356
rect 19628 8316 19892 8344
rect 19628 8313 19640 8316
rect 19582 8307 19640 8313
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 21266 8344 21272 8356
rect 21227 8316 21272 8344
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 21818 8304 21824 8356
rect 21876 8344 21882 8356
rect 22094 8344 22100 8356
rect 21876 8316 22100 8344
rect 21876 8304 21882 8316
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 17920 8044 19257 8072
rect 17920 8032 17926 8044
rect 19245 8041 19257 8044
rect 19291 8072 19303 8075
rect 19334 8072 19340 8084
rect 19291 8044 19340 8072
rect 19291 8041 19303 8044
rect 19245 8035 19303 8041
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 19978 8032 19984 8084
rect 20036 8072 20042 8084
rect 20073 8075 20131 8081
rect 20073 8072 20085 8075
rect 20036 8044 20085 8072
rect 20036 8032 20042 8044
rect 20073 8041 20085 8044
rect 20119 8072 20131 8075
rect 20530 8072 20536 8084
rect 20119 8044 20536 8072
rect 20119 8041 20131 8044
rect 20073 8035 20131 8041
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21177 8075 21235 8081
rect 21177 8041 21189 8075
rect 21223 8072 21235 8075
rect 21542 8072 21548 8084
rect 21223 8044 21548 8072
rect 21223 8041 21235 8044
rect 21177 8035 21235 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 18782 7964 18788 8016
rect 18840 8004 18846 8016
rect 19061 8007 19119 8013
rect 19061 8004 19073 8007
rect 18840 7976 19073 8004
rect 18840 7964 18846 7976
rect 19061 7973 19073 7976
rect 19107 7973 19119 8007
rect 19061 7967 19119 7973
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 17420 7800 17448 7899
rect 17586 7868 17592 7880
rect 17547 7840 17592 7868
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 18322 7828 18328 7880
rect 18380 7868 18386 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 18380 7840 19349 7868
rect 18380 7828 18386 7840
rect 19337 7837 19349 7840
rect 19383 7868 19395 7871
rect 19426 7868 19432 7880
rect 19383 7840 19432 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 17494 7800 17500 7812
rect 17407 7772 17500 7800
rect 17494 7760 17500 7772
rect 17552 7800 17558 7812
rect 18785 7803 18843 7809
rect 18785 7800 18797 7803
rect 17552 7772 18797 7800
rect 17552 7760 17558 7772
rect 18785 7769 18797 7772
rect 18831 7769 18843 7803
rect 18785 7763 18843 7769
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 19705 7735 19763 7741
rect 19705 7732 19717 7735
rect 19116 7704 19717 7732
rect 19116 7692 19122 7704
rect 19705 7701 19717 7704
rect 19751 7701 19763 7735
rect 19705 7695 19763 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17862 7528 17868 7540
rect 17823 7500 17868 7528
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18322 7528 18328 7540
rect 18283 7500 18328 7528
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 18693 7531 18751 7537
rect 18693 7497 18705 7531
rect 18739 7528 18751 7531
rect 18782 7528 18788 7540
rect 18739 7500 18788 7528
rect 18739 7497 18751 7500
rect 18693 7491 18751 7497
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 20530 7528 20536 7540
rect 20491 7500 20536 7528
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7324 4123 7327
rect 19153 7327 19211 7333
rect 19153 7324 19165 7327
rect 4111 7296 4384 7324
rect 4111 7293 4123 7296
rect 4065 7287 4123 7293
rect 4356 7200 4384 7296
rect 19076 7296 19165 7324
rect 19076 7200 19104 7296
rect 19153 7293 19165 7296
rect 19199 7293 19211 7327
rect 19153 7287 19211 7293
rect 19420 7259 19478 7265
rect 19420 7225 19432 7259
rect 19466 7256 19478 7259
rect 19978 7256 19984 7268
rect 19466 7228 19984 7256
rect 19466 7225 19478 7228
rect 19420 7219 19478 7225
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 4246 7188 4252 7200
rect 4207 7160 4252 7188
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4396 7160 4629 7188
rect 4396 7148 4402 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 19058 7188 19064 7200
rect 19019 7160 19064 7188
rect 4617 7151 4675 7157
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 19797 6987 19855 6993
rect 19797 6953 19809 6987
rect 19843 6953 19855 6987
rect 24762 6984 24768 6996
rect 24723 6956 24768 6984
rect 19797 6947 19855 6953
rect 934 6876 940 6928
rect 992 6916 998 6928
rect 1670 6916 1676 6928
rect 992 6888 1676 6916
rect 992 6876 998 6888
rect 1670 6876 1676 6888
rect 1728 6876 1734 6928
rect 18233 6919 18291 6925
rect 18233 6916 18245 6919
rect 18156 6888 18245 6916
rect 18156 6860 18184 6888
rect 18233 6885 18245 6888
rect 18279 6885 18291 6919
rect 18233 6879 18291 6885
rect 19812 6860 19840 6947
rect 24762 6944 24768 6956
rect 24820 6944 24826 6996
rect 21453 6919 21511 6925
rect 21453 6885 21465 6919
rect 21499 6885 21511 6919
rect 21453 6879 21511 6885
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6848 16635 6851
rect 16666 6848 16672 6860
rect 16623 6820 16672 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 16666 6808 16672 6820
rect 16724 6848 16730 6860
rect 17586 6848 17592 6860
rect 16724 6820 17592 6848
rect 16724 6808 16730 6820
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 18046 6848 18052 6860
rect 18007 6820 18052 6848
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 18138 6808 18144 6860
rect 18196 6808 18202 6860
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 19613 6851 19671 6857
rect 19613 6848 19625 6851
rect 18932 6820 19625 6848
rect 18932 6808 18938 6820
rect 19613 6817 19625 6820
rect 19659 6817 19671 6851
rect 19613 6811 19671 6817
rect 19794 6808 19800 6860
rect 19852 6808 19858 6860
rect 21266 6848 21272 6860
rect 21227 6820 21272 6848
rect 21266 6808 21272 6820
rect 21324 6808 21330 6860
rect 21468 6848 21496 6879
rect 21726 6848 21732 6860
rect 21468 6820 21732 6848
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 24581 6851 24639 6857
rect 24581 6817 24593 6851
rect 24627 6848 24639 6851
rect 24670 6848 24676 6860
rect 24627 6820 24676 6848
rect 24627 6817 24639 6820
rect 24581 6811 24639 6817
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 17402 6740 17408 6792
rect 17460 6780 17466 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 17460 6752 18337 6780
rect 17460 6740 17466 6752
rect 18325 6749 18337 6752
rect 18371 6780 18383 6783
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18371 6752 18797 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 18785 6749 18797 6752
rect 18831 6780 18843 6783
rect 19886 6780 19892 6792
rect 18831 6752 19472 6780
rect 19847 6752 19892 6780
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 18138 6672 18144 6724
rect 18196 6712 18202 6724
rect 19337 6715 19395 6721
rect 19337 6712 19349 6715
rect 18196 6684 19349 6712
rect 18196 6672 18202 6684
rect 19337 6681 19349 6684
rect 19383 6681 19395 6715
rect 19444 6712 19472 6752
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 21634 6780 21640 6792
rect 21591 6752 21640 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6780 23167 6783
rect 23474 6780 23480 6792
rect 23155 6752 23480 6780
rect 23155 6749 23167 6752
rect 23109 6743 23167 6749
rect 23474 6740 23480 6752
rect 23532 6740 23538 6792
rect 19978 6712 19984 6724
rect 19444 6684 19984 6712
rect 19337 6675 19395 6681
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6644 16819 6647
rect 17310 6644 17316 6656
rect 16807 6616 17316 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 17770 6644 17776 6656
rect 17731 6616 17776 6644
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 19058 6644 19064 6656
rect 19019 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 20993 6647 21051 6653
rect 20993 6644 21005 6647
rect 20864 6616 21005 6644
rect 20864 6604 20870 6616
rect 20993 6613 21005 6616
rect 21039 6613 21051 6647
rect 20993 6607 21051 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 16666 6440 16672 6452
rect 16627 6412 16672 6440
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 18601 6443 18659 6449
rect 18601 6409 18613 6443
rect 18647 6440 18659 6443
rect 19794 6440 19800 6452
rect 18647 6412 19800 6440
rect 18647 6409 18659 6412
rect 18601 6403 18659 6409
rect 19794 6400 19800 6412
rect 19852 6400 19858 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20441 6443 20499 6449
rect 20441 6440 20453 6443
rect 20036 6412 20453 6440
rect 20036 6400 20042 6412
rect 20441 6409 20453 6412
rect 20487 6409 20499 6443
rect 20441 6403 20499 6409
rect 21453 6443 21511 6449
rect 21453 6409 21465 6443
rect 21499 6440 21511 6443
rect 21726 6440 21732 6452
rect 21499 6412 21732 6440
rect 21499 6409 21511 6412
rect 21453 6403 21511 6409
rect 21726 6400 21732 6412
rect 21784 6400 21790 6452
rect 23842 6400 23848 6452
rect 23900 6400 23906 6452
rect 24670 6440 24676 6452
rect 23952 6412 24676 6440
rect 23860 6316 23888 6400
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6304 17831 6307
rect 18046 6304 18052 6316
rect 17819 6276 18052 6304
rect 17819 6273 17831 6276
rect 17773 6267 17831 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 23842 6264 23848 6316
rect 23900 6264 23906 6316
rect 23952 6313 23980 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 23937 6307 23995 6313
rect 23937 6273 23949 6307
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 18322 6196 18328 6248
rect 18380 6236 18386 6248
rect 19058 6236 19064 6248
rect 18380 6208 19064 6236
rect 18380 6196 18386 6208
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 23477 6239 23535 6245
rect 23477 6205 23489 6239
rect 23523 6236 23535 6239
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23523 6208 23673 6236
rect 23523 6205 23535 6208
rect 23477 6199 23535 6205
rect 23661 6205 23673 6208
rect 23707 6236 23719 6239
rect 23750 6236 23756 6248
rect 23707 6208 23756 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 23750 6196 23756 6208
rect 23808 6196 23814 6248
rect 24946 6236 24952 6248
rect 24859 6208 24952 6236
rect 24946 6196 24952 6208
rect 25004 6236 25010 6248
rect 25501 6239 25559 6245
rect 25501 6236 25513 6239
rect 25004 6208 25513 6236
rect 25004 6196 25010 6208
rect 25501 6205 25513 6208
rect 25547 6205 25559 6239
rect 25501 6199 25559 6205
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 19328 6171 19386 6177
rect 19328 6168 19340 6171
rect 18288 6140 19340 6168
rect 18288 6128 18294 6140
rect 19328 6137 19340 6140
rect 19374 6168 19386 6171
rect 19978 6168 19984 6180
rect 19374 6140 19984 6168
rect 19374 6137 19386 6140
rect 19328 6131 19386 6137
rect 19978 6128 19984 6140
rect 20036 6128 20042 6180
rect 18874 6100 18880 6112
rect 18835 6072 18880 6100
rect 18874 6060 18880 6072
rect 18932 6100 18938 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 18932 6072 21005 6100
rect 18932 6060 18938 6072
rect 20993 6069 21005 6072
rect 21039 6100 21051 6103
rect 21266 6100 21272 6112
rect 21039 6072 21272 6100
rect 21039 6069 21051 6072
rect 20993 6063 21051 6069
rect 21266 6060 21272 6072
rect 21324 6060 21330 6112
rect 21726 6100 21732 6112
rect 21687 6072 21732 6100
rect 21726 6060 21732 6072
rect 21784 6060 21790 6112
rect 24854 6060 24860 6112
rect 24912 6100 24918 6112
rect 25133 6103 25191 6109
rect 25133 6100 25145 6103
rect 24912 6072 25145 6100
rect 24912 6060 24918 6072
rect 25133 6069 25145 6072
rect 25179 6069 25191 6103
rect 25133 6063 25191 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 18138 5896 18144 5908
rect 17819 5868 18144 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 23566 5896 23572 5908
rect 18288 5868 18333 5896
rect 23527 5868 23572 5896
rect 18288 5856 18294 5868
rect 23566 5856 23572 5868
rect 23624 5856 23630 5908
rect 24210 5856 24216 5908
rect 24268 5856 24274 5908
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 19242 5828 19248 5840
rect 9732 5800 19248 5828
rect 9732 5788 9738 5800
rect 19242 5788 19248 5800
rect 19300 5788 19306 5840
rect 22370 5788 22376 5840
rect 22428 5837 22434 5840
rect 22428 5831 22492 5837
rect 22428 5797 22446 5831
rect 22480 5797 22492 5831
rect 22428 5791 22492 5797
rect 22428 5788 22434 5791
rect 16945 5763 17003 5769
rect 16945 5729 16957 5763
rect 16991 5760 17003 5763
rect 17034 5760 17040 5772
rect 16991 5732 17040 5760
rect 16991 5729 17003 5732
rect 16945 5723 17003 5729
rect 17034 5720 17040 5732
rect 17092 5760 17098 5772
rect 17770 5760 17776 5772
rect 17092 5732 17776 5760
rect 17092 5720 17098 5732
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 18598 5769 18604 5772
rect 18592 5760 18604 5769
rect 18559 5732 18604 5760
rect 18592 5723 18604 5732
rect 18598 5720 18604 5723
rect 18656 5720 18662 5772
rect 22094 5720 22100 5772
rect 22152 5760 22158 5772
rect 22189 5763 22247 5769
rect 22189 5760 22201 5763
rect 22152 5732 22201 5760
rect 22152 5720 22158 5732
rect 22189 5729 22201 5732
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 16574 5652 16580 5704
rect 16632 5692 16638 5704
rect 17129 5695 17187 5701
rect 17129 5692 17141 5695
rect 16632 5664 17141 5692
rect 16632 5652 16638 5664
rect 17129 5661 17141 5664
rect 17175 5661 17187 5695
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 17129 5655 17187 5661
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20404 5664 20913 5692
rect 20404 5652 20410 5664
rect 20901 5661 20913 5664
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 24228 5636 24256 5856
rect 24946 5828 24952 5840
rect 24907 5800 24952 5828
rect 24946 5788 24952 5800
rect 25004 5788 25010 5840
rect 24670 5760 24676 5772
rect 24631 5732 24676 5760
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 24210 5584 24216 5636
rect 24268 5584 24274 5636
rect 19702 5556 19708 5568
rect 19663 5528 19708 5556
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20349 5559 20407 5565
rect 20349 5556 20361 5559
rect 20036 5528 20361 5556
rect 20036 5516 20042 5528
rect 20349 5525 20361 5528
rect 20395 5556 20407 5559
rect 20898 5556 20904 5568
rect 20395 5528 20904 5556
rect 20395 5525 20407 5528
rect 20349 5519 20407 5525
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 24118 5556 24124 5568
rect 24079 5528 24124 5556
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 16574 5352 16580 5364
rect 16535 5324 16580 5352
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 17034 5352 17040 5364
rect 16995 5324 17040 5352
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 18598 5312 18604 5364
rect 18656 5352 18662 5364
rect 18693 5355 18751 5361
rect 18693 5352 18705 5355
rect 18656 5324 18705 5352
rect 18656 5312 18662 5324
rect 18693 5321 18705 5324
rect 18739 5321 18751 5355
rect 18693 5315 18751 5321
rect 19521 5355 19579 5361
rect 19521 5321 19533 5355
rect 19567 5352 19579 5355
rect 19610 5352 19616 5364
rect 19567 5324 19616 5352
rect 19567 5321 19579 5324
rect 19521 5315 19579 5321
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20956 5324 21005 5352
rect 20956 5312 20962 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 20993 5315 21051 5321
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22189 5355 22247 5361
rect 22189 5352 22201 5355
rect 22152 5324 22201 5352
rect 22152 5312 22158 5324
rect 22189 5321 22201 5324
rect 22235 5321 22247 5355
rect 23474 5352 23480 5364
rect 23435 5324 23480 5352
rect 22189 5315 22247 5321
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 23750 5352 23756 5364
rect 23711 5324 23756 5352
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 24118 5312 24124 5364
rect 24176 5352 24182 5364
rect 24176 5324 24440 5352
rect 24176 5312 24182 5324
rect 18322 5244 18328 5296
rect 18380 5284 18386 5296
rect 18417 5287 18475 5293
rect 18417 5284 18429 5287
rect 18380 5256 18429 5284
rect 18380 5244 18386 5256
rect 18417 5253 18429 5256
rect 18463 5284 18475 5287
rect 19628 5284 19656 5312
rect 18463 5256 19656 5284
rect 18463 5253 18475 5256
rect 18417 5247 18475 5253
rect 19628 5225 19656 5256
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5185 19671 5219
rect 23492 5216 23520 5312
rect 24121 5219 24179 5225
rect 24121 5216 24133 5219
rect 23492 5188 24133 5216
rect 19613 5179 19671 5185
rect 24121 5185 24133 5188
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5148 15991 5151
rect 16574 5148 16580 5160
rect 15979 5120 16580 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 19702 5080 19708 5092
rect 19168 5052 19708 5080
rect 19168 5024 19196 5052
rect 19702 5040 19708 5052
rect 19760 5080 19766 5092
rect 19858 5083 19916 5089
rect 19858 5080 19870 5083
rect 19760 5052 19870 5080
rect 19760 5040 19766 5052
rect 19858 5049 19870 5052
rect 19904 5049 19916 5083
rect 19858 5043 19916 5049
rect 21913 5083 21971 5089
rect 21913 5049 21925 5083
rect 21959 5080 21971 5083
rect 22370 5080 22376 5092
rect 21959 5052 22376 5080
rect 21959 5049 21971 5052
rect 21913 5043 21971 5049
rect 22370 5040 22376 5052
rect 22428 5080 22434 5092
rect 23109 5083 23167 5089
rect 23109 5080 23121 5083
rect 22428 5052 23121 5080
rect 22428 5040 22434 5052
rect 23109 5049 23121 5052
rect 23155 5080 23167 5083
rect 24302 5080 24308 5092
rect 23155 5052 24308 5080
rect 23155 5049 23167 5052
rect 23109 5043 23167 5049
rect 24302 5040 24308 5052
rect 24360 5040 24366 5092
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 16117 5015 16175 5021
rect 16117 5012 16129 5015
rect 15988 4984 16129 5012
rect 15988 4972 15994 4984
rect 16117 4981 16129 4984
rect 16163 4981 16175 5015
rect 19150 5012 19156 5024
rect 19111 4984 19156 5012
rect 16117 4975 16175 4981
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 22462 4972 22468 5024
rect 22520 5012 22526 5024
rect 22557 5015 22615 5021
rect 22557 5012 22569 5015
rect 22520 4984 22569 5012
rect 22520 4972 22526 4984
rect 22557 4981 22569 4984
rect 22603 4981 22615 5015
rect 22557 4975 22615 4981
rect 23750 4972 23756 5024
rect 23808 5012 23814 5024
rect 24213 5015 24271 5021
rect 24213 5012 24225 5015
rect 23808 4984 24225 5012
rect 23808 4972 23814 4984
rect 24213 4981 24225 4984
rect 24259 5012 24271 5015
rect 24412 5012 24440 5324
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 25222 5108 25228 5120
rect 25280 5148 25286 5160
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25280 5120 25789 5148
rect 25280 5108 25286 5120
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 25777 5111 25835 5117
rect 24670 5012 24676 5024
rect 24259 4984 24440 5012
rect 24631 4984 24676 5012
rect 24259 4981 24271 4984
rect 24213 4975 24271 4981
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 25409 5015 25467 5021
rect 25409 4981 25421 5015
rect 25455 5012 25467 5015
rect 25682 5012 25688 5024
rect 25455 4984 25688 5012
rect 25455 4981 25467 4984
rect 25409 4975 25467 4981
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 18138 4768 18144 4820
rect 18196 4808 18202 4820
rect 18233 4811 18291 4817
rect 18233 4808 18245 4811
rect 18196 4780 18245 4808
rect 18196 4768 18202 4780
rect 18233 4777 18245 4780
rect 18279 4808 18291 4811
rect 18322 4808 18328 4820
rect 18279 4780 18328 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 19153 4811 19211 4817
rect 19153 4777 19165 4811
rect 19199 4808 19211 4811
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19199 4780 19809 4808
rect 19199 4777 19211 4780
rect 19153 4771 19211 4777
rect 19797 4777 19809 4780
rect 19843 4808 19855 4811
rect 20806 4808 20812 4820
rect 19843 4780 20812 4808
rect 19843 4777 19855 4780
rect 19797 4771 19855 4777
rect 20806 4768 20812 4780
rect 20864 4768 20870 4820
rect 22373 4811 22431 4817
rect 22373 4777 22385 4811
rect 22419 4808 22431 4811
rect 23658 4808 23664 4820
rect 22419 4780 23664 4808
rect 22419 4777 22431 4780
rect 22373 4771 22431 4777
rect 23658 4768 23664 4780
rect 23716 4768 23722 4820
rect 24302 4768 24308 4820
rect 24360 4808 24366 4820
rect 24673 4811 24731 4817
rect 24673 4808 24685 4811
rect 24360 4780 24685 4808
rect 24360 4768 24366 4780
rect 24673 4777 24685 4780
rect 24719 4777 24731 4811
rect 24673 4771 24731 4777
rect 6822 4672 6828 4684
rect 6783 4644 6828 4672
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 20346 4672 20352 4684
rect 19659 4644 20352 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 20346 4632 20352 4644
rect 20404 4632 20410 4684
rect 22189 4675 22247 4681
rect 22189 4641 22201 4675
rect 22235 4672 22247 4675
rect 22830 4672 22836 4684
rect 22235 4644 22836 4672
rect 22235 4641 22247 4644
rect 22189 4635 22247 4641
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 23566 4681 23572 4684
rect 23560 4635 23572 4681
rect 23624 4672 23630 4684
rect 23624 4644 23660 4672
rect 23566 4632 23572 4635
rect 23624 4632 23630 4644
rect 15470 4604 15476 4616
rect 15431 4576 15476 4604
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 19889 4607 19947 4613
rect 19889 4604 19901 4607
rect 19208 4576 19901 4604
rect 19208 4564 19214 4576
rect 19889 4573 19901 4576
rect 19935 4573 19947 4607
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 19889 4567 19947 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 23198 4564 23204 4616
rect 23256 4604 23262 4616
rect 23293 4607 23351 4613
rect 23293 4604 23305 4607
rect 23256 4576 23305 4604
rect 23256 4564 23262 4576
rect 23293 4573 23305 4576
rect 23339 4573 23351 4607
rect 23293 4567 23351 4573
rect 7006 4536 7012 4548
rect 6967 4508 7012 4536
rect 7006 4496 7012 4508
rect 7064 4496 7070 4548
rect 19334 4536 19340 4548
rect 19295 4508 19340 4536
rect 19334 4496 19340 4508
rect 19392 4496 19398 4548
rect 22097 4539 22155 4545
rect 22097 4505 22109 4539
rect 22143 4536 22155 4539
rect 22554 4536 22560 4548
rect 22143 4508 22560 4536
rect 22143 4505 22155 4508
rect 22097 4499 22155 4505
rect 22554 4496 22560 4508
rect 22612 4496 22618 4548
rect 21266 4428 21272 4480
rect 21324 4468 21330 4480
rect 21361 4471 21419 4477
rect 21361 4468 21373 4471
rect 21324 4440 21373 4468
rect 21324 4428 21330 4440
rect 21361 4437 21373 4440
rect 21407 4437 21419 4471
rect 22830 4468 22836 4480
rect 22791 4440 22836 4468
rect 21361 4431 21419 4437
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 7650 4264 7656 4276
rect 7611 4236 7656 4264
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 15286 4264 15292 4276
rect 15247 4236 15292 4264
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 20165 4267 20223 4273
rect 20165 4233 20177 4267
rect 20211 4264 20223 4267
rect 20346 4264 20352 4276
rect 20211 4236 20352 4264
rect 20211 4233 20223 4236
rect 20165 4227 20223 4233
rect 20346 4224 20352 4236
rect 20404 4224 20410 4276
rect 20806 4264 20812 4276
rect 20767 4236 20812 4264
rect 20806 4224 20812 4236
rect 20864 4224 20870 4276
rect 23750 4264 23756 4276
rect 23711 4236 23756 4264
rect 23750 4224 23756 4236
rect 23808 4224 23814 4276
rect 24489 4267 24547 4273
rect 24489 4233 24501 4267
rect 24535 4264 24547 4267
rect 24765 4267 24823 4273
rect 24765 4264 24777 4267
rect 24535 4236 24777 4264
rect 24535 4233 24547 4236
rect 24489 4227 24547 4233
rect 24765 4233 24777 4236
rect 24811 4264 24823 4267
rect 25038 4264 25044 4276
rect 24811 4236 25044 4264
rect 24811 4233 24823 4236
rect 24765 4227 24823 4233
rect 25038 4224 25044 4236
rect 25096 4224 25102 4276
rect 15470 4196 15476 4208
rect 15120 4168 15476 4196
rect 14829 4131 14887 4137
rect 14829 4128 14841 4131
rect 14200 4100 14841 4128
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 7742 4060 7748 4072
rect 7515 4032 7748 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 7742 4020 7748 4032
rect 7800 4060 7806 4072
rect 14200 4069 14228 4100
rect 14829 4097 14841 4100
rect 14875 4128 14887 4131
rect 15120 4128 15148 4168
rect 15470 4156 15476 4168
rect 15528 4156 15534 4208
rect 17862 4128 17868 4140
rect 14875 4100 15148 4128
rect 17823 4100 17868 4128
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 17862 4088 17868 4100
rect 17920 4128 17926 4140
rect 20625 4131 20683 4137
rect 17920 4100 18276 4128
rect 17920 4088 17926 4100
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7800 4032 8033 4060
rect 7800 4020 7806 4032
rect 8021 4029 8033 4032
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4029 14243 4063
rect 18138 4060 18144 4072
rect 18099 4032 18144 4060
rect 14185 4023 14243 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 18248 4060 18276 4100
rect 20625 4097 20637 4131
rect 20671 4128 20683 4131
rect 20898 4128 20904 4140
rect 20671 4100 20904 4128
rect 20671 4097 20683 4100
rect 20625 4091 20683 4097
rect 20898 4088 20904 4100
rect 20956 4128 20962 4140
rect 21177 4131 21235 4137
rect 21177 4128 21189 4131
rect 20956 4100 21189 4128
rect 20956 4088 20962 4100
rect 21177 4097 21189 4100
rect 21223 4097 21235 4131
rect 21177 4091 21235 4097
rect 22557 4131 22615 4137
rect 22557 4097 22569 4131
rect 22603 4128 22615 4131
rect 23290 4128 23296 4140
rect 22603 4100 23296 4128
rect 22603 4097 22615 4100
rect 22557 4091 22615 4097
rect 23290 4088 23296 4100
rect 23348 4088 23354 4140
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23750 4128 23756 4140
rect 23532 4100 23756 4128
rect 23532 4088 23538 4100
rect 23750 4088 23756 4100
rect 23808 4088 23814 4140
rect 25406 4128 25412 4140
rect 25367 4100 25412 4128
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 18397 4063 18455 4069
rect 18397 4060 18409 4063
rect 18248 4032 18409 4060
rect 18397 4029 18409 4032
rect 18443 4029 18455 4063
rect 22281 4063 22339 4069
rect 22281 4060 22293 4063
rect 18397 4023 18455 4029
rect 22112 4032 22293 4060
rect 21361 3995 21419 4001
rect 21361 3961 21373 3995
rect 21407 3961 21419 3995
rect 21361 3955 21419 3961
rect 7098 3924 7104 3936
rect 7059 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 14369 3927 14427 3933
rect 14369 3893 14381 3927
rect 14415 3924 14427 3927
rect 14550 3924 14556 3936
rect 14415 3896 14556 3924
rect 14415 3893 14427 3896
rect 14369 3887 14427 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19521 3927 19579 3933
rect 19521 3924 19533 3927
rect 18840 3896 19533 3924
rect 18840 3884 18846 3896
rect 19521 3893 19533 3896
rect 19567 3893 19579 3927
rect 19521 3887 19579 3893
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 21266 3924 21272 3936
rect 20864 3896 21272 3924
rect 20864 3884 20870 3896
rect 21266 3884 21272 3896
rect 21324 3884 21330 3936
rect 21376 3924 21404 3955
rect 22112 3936 22140 4032
rect 22281 4029 22293 4032
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 23566 4020 23572 4072
rect 23624 4060 23630 4072
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 23624 4032 24317 4060
rect 23624 4020 23630 4032
rect 24305 4029 24317 4032
rect 24351 4060 24363 4063
rect 24854 4060 24860 4072
rect 24351 4032 24860 4060
rect 24351 4029 24363 4032
rect 24305 4023 24363 4029
rect 24854 4020 24860 4032
rect 24912 4060 24918 4072
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 24912 4032 25053 4060
rect 24912 4020 24918 4032
rect 25041 4029 25053 4032
rect 25087 4029 25099 4063
rect 25222 4060 25228 4072
rect 25183 4032 25228 4060
rect 25041 4023 25099 4029
rect 25222 4020 25228 4032
rect 25280 4060 25286 4072
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 25280 4032 25973 4060
rect 25280 4020 25286 4032
rect 25961 4029 25973 4032
rect 26007 4029 26019 4063
rect 25961 4023 26019 4029
rect 23474 3992 23480 4004
rect 23435 3964 23480 3992
rect 23474 3952 23480 3964
rect 23532 3992 23538 4004
rect 24029 3995 24087 4001
rect 24029 3992 24041 3995
rect 23532 3964 24041 3992
rect 23532 3952 23538 3964
rect 24029 3961 24041 3964
rect 24075 3961 24087 3995
rect 24029 3955 24087 3961
rect 24213 3995 24271 4001
rect 24213 3961 24225 3995
rect 24259 3992 24271 3995
rect 24489 3995 24547 4001
rect 24489 3992 24501 3995
rect 24259 3964 24501 3992
rect 24259 3961 24271 3964
rect 24213 3955 24271 3961
rect 24489 3961 24501 3964
rect 24535 3961 24547 3995
rect 24489 3955 24547 3961
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 21376 3896 21833 3924
rect 21821 3893 21833 3896
rect 21867 3924 21879 3927
rect 22002 3924 22008 3936
rect 21867 3896 22008 3924
rect 21867 3893 21879 3896
rect 21821 3887 21879 3893
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 23109 3927 23167 3933
rect 22152 3896 22197 3924
rect 22152 3884 22158 3896
rect 23109 3893 23121 3927
rect 23155 3924 23167 3927
rect 23198 3924 23204 3936
rect 23155 3896 23204 3924
rect 23155 3893 23167 3896
rect 23109 3887 23167 3893
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 23934 3884 23940 3936
rect 23992 3924 23998 3936
rect 24228 3924 24256 3955
rect 23992 3896 24256 3924
rect 23992 3884 23998 3896
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 18782 3720 18788 3732
rect 18340 3692 18788 3720
rect 18230 3652 18236 3664
rect 18191 3624 18236 3652
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 18340 3661 18368 3692
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 19150 3720 19156 3732
rect 19111 3692 19156 3720
rect 19150 3680 19156 3692
rect 19208 3680 19214 3732
rect 23385 3723 23443 3729
rect 23385 3689 23397 3723
rect 23431 3720 23443 3723
rect 23566 3720 23572 3732
rect 23431 3692 23572 3720
rect 23431 3689 23443 3692
rect 23385 3683 23443 3689
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 24854 3720 24860 3732
rect 24815 3692 24860 3720
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 18325 3655 18383 3661
rect 18325 3621 18337 3655
rect 18371 3621 18383 3655
rect 18325 3615 18383 3621
rect 19702 3612 19708 3664
rect 19760 3652 19766 3664
rect 19797 3655 19855 3661
rect 19797 3652 19809 3655
rect 19760 3624 19809 3652
rect 19760 3612 19766 3624
rect 19797 3621 19809 3624
rect 19843 3652 19855 3655
rect 20254 3652 20260 3664
rect 19843 3624 20260 3652
rect 19843 3621 19855 3624
rect 19797 3615 19855 3621
rect 20254 3612 20260 3624
rect 20312 3652 20318 3664
rect 23934 3652 23940 3664
rect 20312 3624 23940 3652
rect 20312 3612 20318 3624
rect 23934 3612 23940 3624
rect 23992 3612 23998 3664
rect 8110 3584 8116 3596
rect 8071 3556 8116 3584
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 17586 3544 17592 3596
rect 17644 3584 17650 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17644 3556 18061 3584
rect 17644 3544 17650 3556
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 21174 3593 21180 3596
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 18748 3556 19625 3584
rect 18748 3544 18754 3556
rect 19613 3553 19625 3556
rect 19659 3553 19671 3587
rect 21168 3584 21180 3593
rect 21135 3556 21180 3584
rect 19613 3547 19671 3553
rect 21168 3547 21180 3556
rect 21174 3544 21180 3547
rect 21232 3544 21238 3596
rect 23750 3593 23756 3596
rect 22925 3587 22983 3593
rect 22925 3553 22937 3587
rect 22971 3584 22983 3587
rect 23744 3584 23756 3593
rect 22971 3556 23756 3584
rect 22971 3553 22983 3556
rect 22925 3547 22983 3553
rect 23744 3547 23756 3556
rect 23750 3544 23756 3547
rect 23808 3544 23814 3596
rect 19889 3519 19947 3525
rect 19889 3485 19901 3519
rect 19935 3516 19947 3519
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 19935 3488 20085 3516
rect 19935 3485 19947 3488
rect 19889 3479 19947 3485
rect 20073 3485 20085 3488
rect 20119 3485 20131 3519
rect 20898 3516 20904 3528
rect 20859 3488 20904 3516
rect 20073 3479 20131 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 23477 3519 23535 3525
rect 23477 3516 23489 3519
rect 23256 3488 23489 3516
rect 23256 3476 23262 3488
rect 23477 3485 23489 3488
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 8294 3448 8300 3460
rect 8255 3420 8300 3448
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 19337 3451 19395 3457
rect 19337 3417 19349 3451
rect 19383 3448 19395 3451
rect 20806 3448 20812 3460
rect 19383 3420 20812 3448
rect 19383 3417 19395 3420
rect 19337 3411 19395 3417
rect 20806 3408 20812 3420
rect 20864 3408 20870 3460
rect 16485 3383 16543 3389
rect 16485 3349 16497 3383
rect 16531 3380 16543 3383
rect 16942 3380 16948 3392
rect 16531 3352 16948 3380
rect 16531 3349 16543 3352
rect 16485 3343 16543 3349
rect 16942 3340 16948 3352
rect 17000 3380 17006 3392
rect 17773 3383 17831 3389
rect 17773 3380 17785 3383
rect 17000 3352 17785 3380
rect 17000 3340 17006 3352
rect 17773 3349 17785 3352
rect 17819 3349 17831 3383
rect 17773 3343 17831 3349
rect 20073 3383 20131 3389
rect 20073 3349 20085 3383
rect 20119 3380 20131 3383
rect 20349 3383 20407 3389
rect 20349 3380 20361 3383
rect 20119 3352 20361 3380
rect 20119 3349 20131 3352
rect 20073 3343 20131 3349
rect 20349 3349 20361 3352
rect 20395 3380 20407 3383
rect 20717 3383 20775 3389
rect 20717 3380 20729 3383
rect 20395 3352 20729 3380
rect 20395 3349 20407 3352
rect 20349 3343 20407 3349
rect 20717 3349 20729 3352
rect 20763 3380 20775 3383
rect 21542 3380 21548 3392
rect 20763 3352 21548 3380
rect 20763 3349 20775 3352
rect 20717 3343 20775 3349
rect 21542 3340 21548 3352
rect 21600 3380 21606 3392
rect 22281 3383 22339 3389
rect 22281 3380 22293 3383
rect 21600 3352 22293 3380
rect 21600 3340 21606 3352
rect 22281 3349 22293 3352
rect 22327 3349 22339 3383
rect 22281 3343 22339 3349
rect 23842 3340 23848 3392
rect 23900 3380 23906 3392
rect 24854 3380 24860 3392
rect 23900 3352 24860 3380
rect 23900 3340 23906 3352
rect 24854 3340 24860 3352
rect 24912 3340 24918 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 16482 3176 16488 3188
rect 16443 3148 16488 3176
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 18509 3179 18567 3185
rect 18509 3176 18521 3179
rect 18288 3148 18521 3176
rect 18288 3136 18294 3148
rect 18509 3145 18521 3148
rect 18555 3176 18567 3179
rect 19702 3176 19708 3188
rect 18555 3148 19708 3176
rect 18555 3145 18567 3148
rect 18509 3139 18567 3145
rect 19702 3136 19708 3148
rect 19760 3136 19766 3188
rect 20898 3176 20904 3188
rect 20859 3148 20904 3176
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 22097 3179 22155 3185
rect 22097 3145 22109 3179
rect 22143 3176 22155 3179
rect 23290 3176 23296 3188
rect 22143 3148 23296 3176
rect 22143 3145 22155 3148
rect 22097 3139 22155 3145
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 18690 3068 18696 3120
rect 18748 3108 18754 3120
rect 18785 3111 18843 3117
rect 18785 3108 18797 3111
rect 18748 3080 18797 3108
rect 18748 3068 18754 3080
rect 18785 3077 18797 3080
rect 18831 3077 18843 3111
rect 20916 3108 20944 3136
rect 23198 3108 23204 3120
rect 20916 3080 23204 3108
rect 18785 3071 18843 3077
rect 23198 3068 23204 3080
rect 23256 3068 23262 3120
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18966 3040 18972 3052
rect 18196 3012 18972 3040
rect 18196 3000 18202 3012
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 21913 3043 21971 3049
rect 21913 3009 21925 3043
rect 21959 3040 21971 3043
rect 22462 3040 22468 3052
rect 21959 3012 22468 3040
rect 21959 3009 21971 3012
rect 21913 3003 21971 3009
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 23382 3000 23388 3052
rect 23440 3040 23446 3052
rect 23440 3012 23796 3040
rect 23440 3000 23446 3012
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 9122 2972 9128 2984
rect 8895 2944 9128 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 9122 2932 9128 2944
rect 9180 2972 9186 2984
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 9180 2944 9413 2972
rect 9180 2932 9186 2944
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9401 2935 9459 2941
rect 16666 2932 16672 2984
rect 16724 2972 16730 2984
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 16724 2944 17049 2972
rect 16724 2932 16730 2944
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2904 16359 2907
rect 16758 2904 16764 2916
rect 16347 2876 16764 2904
rect 16347 2873 16359 2876
rect 16301 2867 16359 2873
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 16942 2904 16948 2916
rect 16903 2876 16948 2904
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 17052 2904 17080 2935
rect 18782 2932 18788 2984
rect 18840 2932 18846 2984
rect 23198 2932 23204 2984
rect 23256 2972 23262 2984
rect 23293 2975 23351 2981
rect 23293 2972 23305 2975
rect 23256 2944 23305 2972
rect 23256 2932 23262 2944
rect 23293 2941 23305 2944
rect 23339 2972 23351 2975
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23339 2944 23673 2972
rect 23339 2941 23351 2944
rect 23293 2935 23351 2941
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23768 2972 23796 3012
rect 23768 2944 23888 2972
rect 23661 2935 23719 2941
rect 18800 2904 18828 2932
rect 19214 2907 19272 2913
rect 19214 2904 19226 2907
rect 17052 2876 18552 2904
rect 18800 2876 19226 2904
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 8168 2808 8217 2836
rect 8168 2796 8174 2808
rect 8205 2805 8217 2808
rect 8251 2836 8263 2839
rect 8386 2836 8392 2848
rect 8251 2808 8392 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 9030 2836 9036 2848
rect 8991 2808 9036 2836
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 17586 2796 17592 2848
rect 17644 2836 17650 2848
rect 17681 2839 17739 2845
rect 17681 2836 17693 2839
rect 17644 2808 17693 2836
rect 17644 2796 17650 2808
rect 17681 2805 17693 2808
rect 17727 2805 17739 2839
rect 18524 2836 18552 2876
rect 19214 2873 19226 2876
rect 19260 2873 19272 2907
rect 22554 2904 22560 2916
rect 22515 2876 22560 2904
rect 19214 2867 19272 2873
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 22649 2907 22707 2913
rect 22649 2873 22661 2907
rect 22695 2904 22707 2907
rect 23750 2904 23756 2916
rect 22695 2876 23756 2904
rect 22695 2873 22707 2876
rect 22649 2867 22707 2873
rect 23750 2864 23756 2876
rect 23808 2864 23814 2916
rect 23860 2904 23888 2944
rect 23928 2907 23986 2913
rect 23928 2904 23940 2907
rect 23860 2876 23940 2904
rect 23928 2873 23940 2876
rect 23974 2904 23986 2907
rect 25593 2907 25651 2913
rect 25593 2904 25605 2907
rect 23974 2876 25605 2904
rect 23974 2873 23986 2876
rect 23928 2867 23986 2873
rect 25593 2873 25605 2876
rect 25639 2873 25651 2907
rect 25593 2867 25651 2873
rect 20349 2839 20407 2845
rect 20349 2836 20361 2839
rect 18524 2808 20361 2836
rect 17681 2799 17739 2805
rect 20349 2805 20361 2808
rect 20395 2836 20407 2839
rect 21174 2836 21180 2848
rect 20395 2808 21180 2836
rect 20395 2805 20407 2808
rect 20349 2799 20407 2805
rect 21174 2796 21180 2808
rect 21232 2836 21238 2848
rect 21269 2839 21327 2845
rect 21269 2836 21281 2839
rect 21232 2808 21281 2836
rect 21232 2796 21238 2808
rect 21269 2805 21281 2808
rect 21315 2805 21327 2839
rect 21269 2799 21327 2805
rect 23109 2839 23167 2845
rect 23109 2805 23121 2839
rect 23155 2836 23167 2839
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 23155 2808 23305 2836
rect 23155 2805 23167 2808
rect 23109 2799 23167 2805
rect 23293 2805 23305 2808
rect 23339 2836 23351 2839
rect 23477 2839 23535 2845
rect 23477 2836 23489 2839
rect 23339 2808 23489 2836
rect 23339 2805 23351 2808
rect 23293 2799 23351 2805
rect 23477 2805 23489 2808
rect 23523 2836 23535 2839
rect 23842 2836 23848 2848
rect 23523 2808 23848 2836
rect 23523 2805 23535 2808
rect 23477 2799 23535 2805
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 25038 2836 25044 2848
rect 24999 2808 25044 2836
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 11054 2632 11060 2644
rect 11015 2604 11060 2632
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 16485 2635 16543 2641
rect 16485 2601 16497 2635
rect 16531 2632 16543 2635
rect 16666 2632 16672 2644
rect 16531 2604 16672 2632
rect 16531 2601 16543 2604
rect 16485 2595 16543 2601
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 17221 2635 17279 2641
rect 17221 2632 17233 2635
rect 16816 2604 17233 2632
rect 16816 2592 16822 2604
rect 17221 2601 17233 2604
rect 17267 2601 17279 2635
rect 17221 2595 17279 2601
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 18230 2632 18236 2644
rect 17819 2604 18236 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 18230 2592 18236 2604
rect 18288 2592 18294 2644
rect 18966 2632 18972 2644
rect 18927 2604 18972 2632
rect 18966 2592 18972 2604
rect 19024 2632 19030 2644
rect 20898 2632 20904 2644
rect 19024 2604 20904 2632
rect 19024 2592 19030 2604
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 22002 2592 22008 2644
rect 22060 2632 22066 2644
rect 22557 2635 22615 2641
rect 22557 2632 22569 2635
rect 22060 2604 22569 2632
rect 22060 2592 22066 2604
rect 22557 2601 22569 2604
rect 22603 2632 22615 2635
rect 23382 2632 23388 2644
rect 22603 2604 23388 2632
rect 22603 2601 22615 2604
rect 22557 2595 22615 2601
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 23842 2632 23848 2644
rect 23803 2604 23848 2632
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 18782 2564 18788 2576
rect 18187 2536 18788 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 18782 2524 18788 2536
rect 18840 2524 18846 2576
rect 20073 2567 20131 2573
rect 20073 2533 20085 2567
rect 20119 2564 20131 2567
rect 20254 2564 20260 2576
rect 20119 2536 20260 2564
rect 20119 2533 20131 2536
rect 20073 2527 20131 2533
rect 20254 2524 20260 2536
rect 20312 2564 20318 2576
rect 20533 2567 20591 2573
rect 20533 2564 20545 2567
rect 20312 2536 20545 2564
rect 20312 2524 20318 2536
rect 20533 2533 20545 2536
rect 20579 2533 20591 2567
rect 20533 2527 20591 2533
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3752 2468 4077 2496
rect 3752 2456 3758 2468
rect 4065 2465 4077 2468
rect 4111 2496 4123 2499
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4111 2468 4629 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 5445 2499 5503 2505
rect 5445 2465 5457 2499
rect 5491 2496 5503 2499
rect 5994 2496 6000 2508
rect 5491 2468 6000 2496
rect 5491 2465 5503 2468
rect 5445 2459 5503 2465
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6362 2456 6368 2508
rect 6420 2496 6426 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6420 2468 6929 2496
rect 6420 2456 6426 2468
rect 6917 2465 6929 2468
rect 6963 2496 6975 2499
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 6963 2468 7481 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7469 2465 7481 2468
rect 7515 2465 7527 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 7469 2459 7527 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9824 2468 10333 2496
rect 9824 2456 9830 2468
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 10873 2499 10931 2505
rect 10873 2465 10885 2499
rect 10919 2496 10931 2499
rect 11146 2496 11152 2508
rect 10919 2468 11152 2496
rect 10919 2465 10931 2468
rect 10873 2459 10931 2465
rect 11146 2456 11152 2468
rect 11204 2456 11210 2508
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2496 12679 2499
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12667 2468 13185 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 18414 2496 18420 2508
rect 18375 2468 18420 2496
rect 13173 2459 13231 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 20162 2496 20168 2508
rect 19352 2468 20168 2496
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 19352 2428 19380 2468
rect 20162 2456 20168 2468
rect 20220 2456 20226 2508
rect 20916 2496 20944 2592
rect 21444 2567 21502 2573
rect 21444 2533 21456 2567
rect 21490 2564 21502 2567
rect 21542 2564 21548 2576
rect 21490 2536 21548 2564
rect 21490 2533 21502 2536
rect 21444 2527 21502 2533
rect 21542 2524 21548 2536
rect 21600 2524 21606 2576
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20916 2468 21189 2496
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 23860 2496 23888 2592
rect 23934 2524 23940 2576
rect 23992 2564 23998 2576
rect 24274 2567 24332 2573
rect 24274 2564 24286 2567
rect 23992 2536 24286 2564
rect 23992 2524 23998 2536
rect 24274 2533 24286 2536
rect 24320 2564 24332 2567
rect 25038 2564 25044 2576
rect 24320 2536 25044 2564
rect 24320 2533 24332 2536
rect 24274 2527 24332 2533
rect 25038 2524 25044 2536
rect 25096 2564 25102 2576
rect 25961 2567 26019 2573
rect 25961 2564 25973 2567
rect 25096 2536 25973 2564
rect 25096 2524 25102 2536
rect 25961 2533 25973 2536
rect 26007 2533 26019 2567
rect 25961 2527 26019 2533
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23860 2468 24041 2496
rect 21177 2459 21235 2465
rect 24029 2465 24041 2468
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 19981 2431 20039 2437
rect 19981 2428 19993 2431
rect 17175 2400 19380 2428
rect 19444 2400 19993 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 5629 2363 5687 2369
rect 5629 2329 5641 2363
rect 5675 2360 5687 2363
rect 6822 2360 6828 2372
rect 5675 2332 6828 2360
rect 5675 2329 5687 2332
rect 5629 2323 5687 2329
rect 6822 2320 6828 2332
rect 6880 2320 6886 2372
rect 19444 2304 19472 2400
rect 19981 2397 19993 2400
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 19613 2363 19671 2369
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 20622 2360 20628 2372
rect 19659 2332 20628 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 4246 2292 4252 2304
rect 4207 2264 4252 2292
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 5994 2292 6000 2304
rect 5955 2264 6000 2292
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 7101 2295 7159 2301
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 8202 2292 8208 2304
rect 7147 2264 8208 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 9950 2292 9956 2304
rect 9911 2264 9956 2292
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11425 2295 11483 2301
rect 11425 2292 11437 2295
rect 11204 2264 11437 2292
rect 11204 2252 11210 2264
rect 11425 2261 11437 2264
rect 11471 2261 11483 2295
rect 12802 2292 12808 2304
rect 12763 2264 12808 2292
rect 11425 2255 11483 2261
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 16114 2292 16120 2304
rect 16075 2264 16120 2292
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 18598 2292 18604 2304
rect 18559 2264 18604 2292
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 19426 2292 19432 2304
rect 19387 2264 19432 2292
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 23477 2295 23535 2301
rect 23477 2261 23489 2295
rect 23523 2292 23535 2295
rect 23750 2292 23756 2304
rect 23523 2264 23756 2292
rect 23523 2261 23535 2264
rect 23477 2255 23535 2261
rect 23750 2252 23756 2264
rect 23808 2292 23814 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 23808 2264 25421 2292
rect 23808 2252 23814 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 13906 552 13912 604
rect 13964 592 13970 604
rect 14182 592 14188 604
rect 13964 564 14188 592
rect 13964 552 13970 564
rect 14182 552 14188 564
rect 14240 552 14246 604
rect 17678 552 17684 604
rect 17736 592 17742 604
rect 17954 592 17960 604
rect 17736 564 17960 592
rect 17736 552 17742 564
rect 17954 552 17960 564
rect 18012 552 18018 604
<< via1 >>
rect 20904 26664 20956 26716
rect 24124 26664 24176 26716
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 21732 24896 21784 24948
rect 23756 24896 23808 24948
rect 15476 24828 15528 24880
rect 24768 24828 24820 24880
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 15476 23851 15528 23860
rect 15476 23817 15485 23851
rect 15485 23817 15519 23851
rect 15519 23817 15528 23851
rect 15476 23808 15528 23817
rect 24676 23808 24728 23860
rect 15476 23604 15528 23656
rect 24676 23604 24728 23656
rect 14832 23468 14884 23520
rect 23664 23468 23716 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 16304 21879 16356 21888
rect 16304 21845 16313 21879
rect 16313 21845 16347 21879
rect 16347 21845 16356 21879
rect 16304 21836 16356 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 16120 21675 16172 21684
rect 16120 21641 16129 21675
rect 16129 21641 16163 21675
rect 16163 21641 16172 21675
rect 16120 21632 16172 21641
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 23572 21088 23624 21140
rect 23940 21088 23992 21140
rect 17500 20995 17552 21004
rect 17500 20961 17509 20995
rect 17509 20961 17543 20995
rect 17543 20961 17552 20995
rect 17500 20952 17552 20961
rect 17684 20791 17736 20800
rect 17684 20757 17693 20791
rect 17693 20757 17727 20791
rect 17727 20757 17736 20791
rect 17684 20748 17736 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 24032 19864 24084 19916
rect 24676 19864 24728 19916
rect 24768 19703 24820 19712
rect 24768 19669 24777 19703
rect 24777 19669 24811 19703
rect 24811 19669 24820 19703
rect 24768 19660 24820 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 24032 19456 24084 19508
rect 16120 19252 16172 19304
rect 16304 19252 16356 19304
rect 19524 19227 19576 19236
rect 19524 19193 19533 19227
rect 19533 19193 19567 19227
rect 19567 19193 19576 19227
rect 19524 19184 19576 19193
rect 18972 19116 19024 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 19984 18776 20036 18828
rect 20076 18572 20128 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 19984 18368 20036 18420
rect 20904 18411 20956 18420
rect 20904 18377 20913 18411
rect 20913 18377 20947 18411
rect 20947 18377 20956 18411
rect 20904 18368 20956 18377
rect 20904 18164 20956 18216
rect 20444 18071 20496 18080
rect 20444 18037 20453 18071
rect 20453 18037 20487 18071
rect 20487 18037 20496 18071
rect 20444 18028 20496 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 20996 17688 21048 17740
rect 21180 17484 21232 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 21916 16736 21968 16788
rect 21640 16643 21692 16652
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 21640 16235 21692 16244
rect 21640 16201 21649 16235
rect 21649 16201 21683 16235
rect 21683 16201 21692 16235
rect 21640 16192 21692 16201
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 23388 15512 23440 15564
rect 23388 15351 23440 15360
rect 23388 15317 23397 15351
rect 23397 15317 23431 15351
rect 23431 15317 23440 15351
rect 23388 15308 23440 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 24768 15104 24820 15156
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 25228 14059 25280 14068
rect 25228 14025 25237 14059
rect 25237 14025 25271 14059
rect 25271 14025 25280 14059
rect 25228 14016 25280 14025
rect 23848 13948 23900 14000
rect 25228 13812 25280 13864
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 24860 13336 24912 13388
rect 24216 13200 24268 13252
rect 25044 13200 25096 13252
rect 24676 13132 24728 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 24860 12928 24912 12980
rect 23940 12860 23992 12912
rect 25320 12928 25372 12980
rect 24584 12588 24636 12640
rect 24768 12588 24820 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 23480 12384 23532 12436
rect 23664 12384 23716 12436
rect 23756 12384 23808 12436
rect 23940 12384 23992 12436
rect 24032 12384 24084 12436
rect 24676 12384 24728 12436
rect 24676 12248 24728 12300
rect 24032 12180 24084 12232
rect 24124 12180 24176 12232
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 14188 11543 14240 11552
rect 14188 11509 14197 11543
rect 14197 11509 14231 11543
rect 14231 11509 14240 11543
rect 14188 11500 14240 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 20720 11024 20772 11076
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 19984 10684 20036 10736
rect 20352 10727 20404 10736
rect 20352 10693 20361 10727
rect 20361 10693 20395 10727
rect 20395 10693 20404 10727
rect 20352 10684 20404 10693
rect 22284 10616 22336 10668
rect 1676 10548 1728 10600
rect 20628 10523 20680 10532
rect 20628 10489 20637 10523
rect 20637 10489 20671 10523
rect 20671 10489 20680 10523
rect 20628 10480 20680 10489
rect 20720 10480 20772 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 20628 10208 20680 10260
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 1492 10072 1544 10124
rect 20812 10072 20864 10124
rect 21548 10072 21600 10124
rect 1584 9979 1636 9988
rect 1584 9945 1593 9979
rect 1593 9945 1627 9979
rect 1627 9945 1636 9979
rect 1584 9936 1636 9945
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 16120 9664 16172 9716
rect 16212 9664 16264 9716
rect 20812 9664 20864 9716
rect 21824 9707 21876 9716
rect 21824 9673 21833 9707
rect 21833 9673 21867 9707
rect 21867 9673 21876 9707
rect 21824 9664 21876 9673
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 2320 9324 2372 9376
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 21548 9324 21600 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 18880 9120 18932 9172
rect 20168 9120 20220 9172
rect 21456 9163 21508 9172
rect 21456 9129 21465 9163
rect 21465 9129 21499 9163
rect 21499 9129 21508 9163
rect 21456 9120 21508 9129
rect 2964 8984 3016 9036
rect 19248 8984 19300 9036
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 22468 9027 22520 9036
rect 22468 8993 22477 9027
rect 22477 8993 22511 9027
rect 22511 8993 22520 9027
rect 22468 8984 22520 8993
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 21548 8959 21600 8968
rect 21548 8925 21557 8959
rect 21557 8925 21591 8959
rect 21591 8925 21600 8959
rect 21548 8916 21600 8925
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 2872 8891 2924 8900
rect 2872 8857 2881 8891
rect 2881 8857 2915 8891
rect 2915 8857 2924 8891
rect 2872 8848 2924 8857
rect 20720 8848 20772 8900
rect 19340 8823 19392 8832
rect 19340 8789 19349 8823
rect 19349 8789 19383 8823
rect 19383 8789 19392 8823
rect 19340 8780 19392 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 18880 8619 18932 8628
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 19524 8576 19576 8628
rect 21456 8576 21508 8628
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 19064 8440 19116 8492
rect 18880 8372 18932 8424
rect 19248 8372 19300 8424
rect 2964 8304 3016 8356
rect 19892 8304 19944 8356
rect 21272 8347 21324 8356
rect 21272 8313 21281 8347
rect 21281 8313 21315 8347
rect 21315 8313 21324 8347
rect 21272 8304 21324 8313
rect 21824 8304 21876 8356
rect 22100 8304 22152 8356
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 17868 8032 17920 8084
rect 19340 8032 19392 8084
rect 19984 8032 20036 8084
rect 20536 8032 20588 8084
rect 21548 8032 21600 8084
rect 18788 7964 18840 8016
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 18328 7828 18380 7880
rect 19432 7828 19484 7880
rect 17500 7760 17552 7812
rect 19064 7692 19116 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 18788 7488 18840 7540
rect 20536 7531 20588 7540
rect 20536 7497 20545 7531
rect 20545 7497 20579 7531
rect 20579 7497 20588 7531
rect 20536 7488 20588 7497
rect 19984 7216 20036 7268
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 4344 7148 4396 7200
rect 19064 7191 19116 7200
rect 19064 7157 19073 7191
rect 19073 7157 19107 7191
rect 19107 7157 19116 7191
rect 19064 7148 19116 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 24768 6987 24820 6996
rect 940 6876 992 6928
rect 1676 6876 1728 6928
rect 24768 6953 24777 6987
rect 24777 6953 24811 6987
rect 24811 6953 24820 6987
rect 24768 6944 24820 6953
rect 16672 6808 16724 6860
rect 17592 6808 17644 6860
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 18144 6808 18196 6860
rect 18880 6808 18932 6860
rect 19800 6808 19852 6860
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 21732 6808 21784 6860
rect 24676 6808 24728 6860
rect 17408 6740 17460 6792
rect 19892 6783 19944 6792
rect 18144 6672 18196 6724
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 21640 6740 21692 6792
rect 23480 6740 23532 6792
rect 19984 6672 20036 6724
rect 17316 6604 17368 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 20812 6604 20864 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 19800 6400 19852 6452
rect 19984 6400 20036 6452
rect 21732 6400 21784 6452
rect 23848 6400 23900 6452
rect 24676 6443 24728 6452
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 23848 6264 23900 6316
rect 24676 6409 24685 6443
rect 24685 6409 24719 6443
rect 24719 6409 24728 6443
rect 24676 6400 24728 6409
rect 18328 6196 18380 6248
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 23756 6196 23808 6248
rect 24952 6239 25004 6248
rect 24952 6205 24961 6239
rect 24961 6205 24995 6239
rect 24995 6205 25004 6239
rect 24952 6196 25004 6205
rect 18236 6128 18288 6180
rect 19984 6128 20036 6180
rect 18880 6103 18932 6112
rect 18880 6069 18889 6103
rect 18889 6069 18923 6103
rect 18923 6069 18932 6103
rect 18880 6060 18932 6069
rect 21272 6060 21324 6112
rect 21732 6103 21784 6112
rect 21732 6069 21741 6103
rect 21741 6069 21775 6103
rect 21775 6069 21784 6103
rect 21732 6060 21784 6069
rect 24860 6060 24912 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 18144 5856 18196 5908
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 23572 5899 23624 5908
rect 18236 5856 18288 5865
rect 23572 5865 23581 5899
rect 23581 5865 23615 5899
rect 23615 5865 23624 5899
rect 23572 5856 23624 5865
rect 24216 5856 24268 5908
rect 9680 5788 9732 5840
rect 19248 5788 19300 5840
rect 22376 5788 22428 5840
rect 17040 5720 17092 5772
rect 17776 5720 17828 5772
rect 18604 5763 18656 5772
rect 18604 5729 18638 5763
rect 18638 5729 18656 5763
rect 18604 5720 18656 5729
rect 22100 5720 22152 5772
rect 16580 5652 16632 5704
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 20352 5652 20404 5704
rect 24952 5831 25004 5840
rect 24952 5797 24961 5831
rect 24961 5797 24995 5831
rect 24995 5797 25004 5831
rect 24952 5788 25004 5797
rect 24676 5763 24728 5772
rect 24676 5729 24685 5763
rect 24685 5729 24719 5763
rect 24719 5729 24728 5763
rect 24676 5720 24728 5729
rect 24216 5584 24268 5636
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 19984 5516 20036 5568
rect 20904 5516 20956 5568
rect 24124 5559 24176 5568
rect 24124 5525 24133 5559
rect 24133 5525 24167 5559
rect 24167 5525 24176 5559
rect 24124 5516 24176 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 16580 5355 16632 5364
rect 16580 5321 16589 5355
rect 16589 5321 16623 5355
rect 16623 5321 16632 5355
rect 16580 5312 16632 5321
rect 17040 5355 17092 5364
rect 17040 5321 17049 5355
rect 17049 5321 17083 5355
rect 17083 5321 17092 5355
rect 17040 5312 17092 5321
rect 18604 5312 18656 5364
rect 19616 5312 19668 5364
rect 20904 5312 20956 5364
rect 22100 5312 22152 5364
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 23756 5355 23808 5364
rect 23756 5321 23765 5355
rect 23765 5321 23799 5355
rect 23799 5321 23808 5355
rect 23756 5312 23808 5321
rect 24124 5312 24176 5364
rect 18328 5244 18380 5296
rect 16580 5108 16632 5160
rect 19708 5040 19760 5092
rect 22376 5040 22428 5092
rect 24308 5083 24360 5092
rect 24308 5049 24317 5083
rect 24317 5049 24351 5083
rect 24351 5049 24360 5083
rect 24308 5040 24360 5049
rect 15936 4972 15988 5024
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 22468 4972 22520 5024
rect 23756 4972 23808 5024
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 25688 4972 25740 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 18144 4768 18196 4820
rect 18328 4768 18380 4820
rect 20812 4768 20864 4820
rect 23664 4768 23716 4820
rect 24308 4768 24360 4820
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 20352 4632 20404 4684
rect 22836 4632 22888 4684
rect 23572 4675 23624 4684
rect 23572 4641 23606 4675
rect 23606 4641 23624 4675
rect 23572 4632 23624 4641
rect 15476 4607 15528 4616
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 19156 4564 19208 4616
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 23204 4564 23256 4616
rect 7012 4539 7064 4548
rect 7012 4505 7021 4539
rect 7021 4505 7055 4539
rect 7055 4505 7064 4539
rect 7012 4496 7064 4505
rect 19340 4539 19392 4548
rect 19340 4505 19349 4539
rect 19349 4505 19383 4539
rect 19383 4505 19392 4539
rect 19340 4496 19392 4505
rect 22560 4496 22612 4548
rect 21272 4428 21324 4480
rect 22836 4471 22888 4480
rect 22836 4437 22845 4471
rect 22845 4437 22879 4471
rect 22879 4437 22888 4471
rect 22836 4428 22888 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 7656 4267 7708 4276
rect 7656 4233 7665 4267
rect 7665 4233 7699 4267
rect 7699 4233 7708 4267
rect 7656 4224 7708 4233
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 20352 4224 20404 4276
rect 20812 4267 20864 4276
rect 20812 4233 20821 4267
rect 20821 4233 20855 4267
rect 20855 4233 20864 4267
rect 20812 4224 20864 4233
rect 23756 4267 23808 4276
rect 23756 4233 23765 4267
rect 23765 4233 23799 4267
rect 23799 4233 23808 4267
rect 23756 4224 23808 4233
rect 25044 4224 25096 4276
rect 7748 4020 7800 4072
rect 15476 4156 15528 4208
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 18144 4063 18196 4072
rect 18144 4029 18153 4063
rect 18153 4029 18187 4063
rect 18187 4029 18196 4063
rect 18144 4020 18196 4029
rect 20904 4088 20956 4140
rect 23296 4088 23348 4140
rect 23480 4088 23532 4140
rect 23756 4088 23808 4140
rect 25412 4131 25464 4140
rect 25412 4097 25421 4131
rect 25421 4097 25455 4131
rect 25455 4097 25464 4131
rect 25412 4088 25464 4097
rect 7104 3927 7156 3936
rect 7104 3893 7113 3927
rect 7113 3893 7147 3927
rect 7147 3893 7156 3927
rect 7104 3884 7156 3893
rect 14556 3884 14608 3936
rect 18788 3884 18840 3936
rect 20812 3884 20864 3936
rect 21272 3927 21324 3936
rect 21272 3893 21281 3927
rect 21281 3893 21315 3927
rect 21315 3893 21324 3927
rect 21272 3884 21324 3893
rect 23572 4020 23624 4072
rect 24860 4020 24912 4072
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 23480 3995 23532 4004
rect 23480 3961 23489 3995
rect 23489 3961 23523 3995
rect 23523 3961 23532 3995
rect 23480 3952 23532 3961
rect 22008 3884 22060 3936
rect 22100 3927 22152 3936
rect 22100 3893 22109 3927
rect 22109 3893 22143 3927
rect 22143 3893 22152 3927
rect 22100 3884 22152 3893
rect 23204 3884 23256 3936
rect 23940 3884 23992 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 18788 3723 18840 3732
rect 18236 3655 18288 3664
rect 18236 3621 18245 3655
rect 18245 3621 18279 3655
rect 18279 3621 18288 3655
rect 18236 3612 18288 3621
rect 18788 3689 18797 3723
rect 18797 3689 18831 3723
rect 18831 3689 18840 3723
rect 18788 3680 18840 3689
rect 19156 3723 19208 3732
rect 19156 3689 19165 3723
rect 19165 3689 19199 3723
rect 19199 3689 19208 3723
rect 19156 3680 19208 3689
rect 23572 3680 23624 3732
rect 24860 3723 24912 3732
rect 24860 3689 24869 3723
rect 24869 3689 24903 3723
rect 24903 3689 24912 3723
rect 24860 3680 24912 3689
rect 19708 3612 19760 3664
rect 20260 3612 20312 3664
rect 23940 3612 23992 3664
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 17592 3544 17644 3596
rect 18696 3544 18748 3596
rect 21180 3587 21232 3596
rect 21180 3553 21214 3587
rect 21214 3553 21232 3587
rect 21180 3544 21232 3553
rect 23756 3587 23808 3596
rect 23756 3553 23790 3587
rect 23790 3553 23808 3587
rect 23756 3544 23808 3553
rect 20904 3519 20956 3528
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 23204 3476 23256 3528
rect 8300 3451 8352 3460
rect 8300 3417 8309 3451
rect 8309 3417 8343 3451
rect 8343 3417 8352 3451
rect 8300 3408 8352 3417
rect 20812 3408 20864 3460
rect 16948 3340 17000 3392
rect 21548 3340 21600 3392
rect 23848 3340 23900 3392
rect 24860 3340 24912 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 18236 3136 18288 3188
rect 19708 3136 19760 3188
rect 20904 3179 20956 3188
rect 20904 3145 20913 3179
rect 20913 3145 20947 3179
rect 20947 3145 20956 3179
rect 20904 3136 20956 3145
rect 23296 3136 23348 3188
rect 18696 3068 18748 3120
rect 23204 3068 23256 3120
rect 18144 3000 18196 3052
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 22468 3043 22520 3052
rect 22468 3009 22477 3043
rect 22477 3009 22511 3043
rect 22511 3009 22520 3043
rect 22468 3000 22520 3009
rect 23388 3000 23440 3052
rect 9128 2932 9180 2984
rect 16672 2932 16724 2984
rect 16764 2907 16816 2916
rect 16764 2873 16773 2907
rect 16773 2873 16807 2907
rect 16807 2873 16816 2907
rect 16764 2864 16816 2873
rect 16948 2907 17000 2916
rect 16948 2873 16957 2907
rect 16957 2873 16991 2907
rect 16991 2873 17000 2907
rect 16948 2864 17000 2873
rect 18788 2932 18840 2984
rect 23204 2932 23256 2984
rect 8116 2796 8168 2848
rect 8392 2796 8444 2848
rect 9036 2839 9088 2848
rect 9036 2805 9045 2839
rect 9045 2805 9079 2839
rect 9079 2805 9088 2839
rect 9036 2796 9088 2805
rect 17592 2796 17644 2848
rect 22560 2907 22612 2916
rect 22560 2873 22569 2907
rect 22569 2873 22603 2907
rect 22603 2873 22612 2907
rect 22560 2864 22612 2873
rect 23756 2864 23808 2916
rect 21180 2796 21232 2848
rect 23848 2796 23900 2848
rect 25044 2839 25096 2848
rect 25044 2805 25053 2839
rect 25053 2805 25087 2839
rect 25087 2805 25096 2839
rect 25044 2796 25096 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 16672 2592 16724 2644
rect 16764 2592 16816 2644
rect 18236 2592 18288 2644
rect 18972 2635 19024 2644
rect 18972 2601 18981 2635
rect 18981 2601 19015 2635
rect 19015 2601 19024 2635
rect 20904 2635 20956 2644
rect 18972 2592 19024 2601
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 22008 2592 22060 2644
rect 23388 2592 23440 2644
rect 23848 2635 23900 2644
rect 23848 2601 23857 2635
rect 23857 2601 23891 2635
rect 23891 2601 23900 2635
rect 23848 2592 23900 2601
rect 18788 2524 18840 2576
rect 20260 2524 20312 2576
rect 3700 2456 3752 2508
rect 6000 2456 6052 2508
rect 6368 2456 6420 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 11152 2456 11204 2508
rect 12532 2456 12584 2508
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 20168 2499 20220 2508
rect 20168 2465 20177 2499
rect 20177 2465 20211 2499
rect 20211 2465 20220 2499
rect 20168 2456 20220 2465
rect 21548 2524 21600 2576
rect 23940 2524 23992 2576
rect 25044 2524 25096 2576
rect 6828 2320 6880 2372
rect 20628 2320 20680 2372
rect 4252 2295 4304 2304
rect 4252 2261 4261 2295
rect 4261 2261 4295 2295
rect 4295 2261 4304 2295
rect 4252 2252 4304 2261
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 8208 2252 8260 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 11152 2252 11204 2304
rect 12808 2295 12860 2304
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 12808 2252 12860 2261
rect 16120 2295 16172 2304
rect 16120 2261 16129 2295
rect 16129 2261 16163 2295
rect 16163 2261 16172 2295
rect 16120 2252 16172 2261
rect 18604 2295 18656 2304
rect 18604 2261 18613 2295
rect 18613 2261 18647 2295
rect 18647 2261 18656 2295
rect 18604 2252 18656 2261
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 23756 2252 23808 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 13912 552 13964 604
rect 14188 552 14240 604
rect 17684 552 17736 604
rect 17960 552 18012 604
<< metal2 >>
rect 14002 27520 14058 28000
rect 24122 27704 24178 27713
rect 24122 27639 24178 27648
rect 14016 27418 14044 27520
rect 14016 27390 14320 27418
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 13818 12744 13874 12753
rect 13818 12679 13874 12688
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 13832 11898 13860 12679
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 1676 10600 1728 10606
rect 1582 10568 1638 10577
rect 1676 10542 1728 10548
rect 1582 10503 1638 10512
rect 1596 10470 1624 10503
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 9874 1532 10066
rect 1582 10024 1638 10033
rect 1582 9959 1584 9968
rect 1636 9959 1638 9968
rect 1584 9930 1636 9936
rect 1504 9846 1624 9874
rect 1596 9382 1624 9846
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 940 6928 992 6934
rect 940 6870 992 6876
rect 294 3088 350 3097
rect 294 3023 350 3032
rect 308 480 336 3023
rect 952 480 980 6870
rect 1596 480 1624 9318
rect 1688 6934 1716 10542
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 2226 9480 2282 9489
rect 2226 9415 2282 9424
rect 2240 9382 2268 9415
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 1676 6928 1728 6934
rect 1676 6870 1728 6876
rect 2332 480 2360 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2870 8936 2926 8945
rect 2870 8871 2872 8880
rect 2924 8871 2926 8880
rect 2872 8842 2924 8848
rect 2976 8362 3004 8978
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2976 480 3004 8298
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4250 7304 4306 7313
rect 4250 7239 4306 7248
rect 4264 7206 4292 7239
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3712 480 3740 2450
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4264 1465 4292 2246
rect 4250 1456 4306 1465
rect 4250 1391 4306 1400
rect 4356 480 4384 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 9680 5840 9732 5846
rect 7654 5808 7710 5817
rect 7654 5743 7710 5752
rect 9678 5808 9680 5817
rect 9732 5808 9734 5817
rect 9678 5743 9734 5752
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6840 4162 6868 4626
rect 7010 4584 7066 4593
rect 7010 4519 7012 4528
rect 7064 4519 7066 4528
rect 7012 4490 7064 4496
rect 7668 4282 7696 5743
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 6840 4134 7144 4162
rect 4986 4040 5042 4049
rect 4986 3975 5042 3984
rect 5000 480 5028 3975
rect 7116 3942 7144 4134
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6012 2310 6040 2450
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 1578 6040 2246
rect 5736 1550 6040 1578
rect 5736 480 5764 1550
rect 6380 480 6408 2450
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6840 1601 6868 2314
rect 6826 1592 6882 1601
rect 6826 1527 6882 1536
rect 7116 480 7144 3878
rect 7760 480 7788 4014
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 2854 8156 3538
rect 8298 3496 8354 3505
rect 8298 3431 8300 3440
rect 8352 3431 8354 3440
rect 8300 3402 8352 3408
rect 11886 3088 11942 3097
rect 11886 3023 11942 3032
rect 9128 2984 9180 2990
rect 9034 2952 9090 2961
rect 9128 2926 9180 2932
rect 9034 2887 9090 2896
rect 9048 2854 9076 2887
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 1873 8248 2246
rect 8206 1864 8262 1873
rect 8206 1799 8262 1808
rect 8404 480 8432 2790
rect 9140 480 9168 2926
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11072 2553 11100 2586
rect 11058 2544 11114 2553
rect 9772 2508 9824 2514
rect 11058 2479 11114 2488
rect 11152 2508 11204 2514
rect 9772 2450 9824 2456
rect 11152 2450 11204 2456
rect 9784 480 9812 2450
rect 11164 2310 11192 2450
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 9968 2145 9996 2246
rect 9954 2136 10010 2145
rect 9954 2071 10010 2080
rect 10506 1728 10562 1737
rect 10506 1663 10562 1672
rect 10520 480 10548 1663
rect 11164 480 11192 2246
rect 11900 480 11928 3023
rect 13174 2816 13230 2825
rect 13174 2751 13230 2760
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12544 480 12572 2450
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12820 1057 12848 2246
rect 12806 1048 12862 1057
rect 12806 983 12862 992
rect 13188 480 13216 2751
rect 14200 610 14228 11494
rect 14292 10713 14320 27390
rect 24136 26722 24164 27639
rect 24214 27024 24270 27033
rect 24214 26959 24270 26968
rect 20904 26716 20956 26722
rect 20904 26658 20956 26664
rect 24124 26716 24176 26722
rect 24124 26658 24176 26664
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15476 24880 15528 24886
rect 15476 24822 15528 24828
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15488 23866 15516 24822
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15488 23662 15516 23802
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14278 10704 14334 10713
rect 14278 10639 14334 10648
rect 14844 4026 14872 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 16118 22672 16174 22681
rect 16118 22607 16174 22616
rect 16132 22098 16160 22607
rect 17498 22536 17554 22545
rect 17498 22471 17554 22480
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 16132 21690 16160 22034
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 16316 19310 16344 21830
rect 17512 21010 17540 22471
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17512 20602 17540 20946
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 16132 9722 16160 19246
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15290 4720 15346 4729
rect 15290 4655 15292 4664
rect 15344 4655 15346 4664
rect 15292 4626 15344 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4282 15332 4626
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15488 4214 15516 4558
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 14844 3998 15332 4026
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14462 2544 14518 2553
rect 14462 2479 14518 2488
rect 14476 2009 14504 2479
rect 14462 2000 14518 2009
rect 14462 1935 14518 1944
rect 13912 604 13964 610
rect 13912 546 13964 552
rect 14188 604 14240 610
rect 14188 546 14240 552
rect 13924 480 13952 546
rect 14568 480 14596 3878
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14738 2544 14794 2553
rect 14738 2479 14794 2488
rect 14752 2145 14780 2479
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14738 2136 14794 2145
rect 14956 2128 15252 2148
rect 14738 2071 14794 2080
rect 15304 480 15332 3998
rect 15948 480 15976 4966
rect 16120 2304 16172 2310
rect 16118 2272 16120 2281
rect 16224 2292 16252 9658
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17512 7546 17540 7754
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17604 6866 17632 7822
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 16684 6458 16712 6802
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5370 16620 5646
rect 17052 5370 17080 5714
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16592 5166 16620 5306
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16486 3224 16542 3233
rect 16486 3159 16488 3168
rect 16540 3159 16542 3168
rect 16488 3130 16540 3136
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16684 2650 16712 2926
rect 16960 2922 16988 3334
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16776 2650 16804 2858
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16172 2272 16174 2281
rect 16224 2264 16620 2292
rect 16118 2207 16174 2216
rect 16592 480 16620 2264
rect 17038 2136 17094 2145
rect 17038 2071 17094 2080
rect 17052 1737 17080 2071
rect 17038 1728 17094 1737
rect 17038 1663 17094 1672
rect 17222 1728 17278 1737
rect 17222 1663 17278 1672
rect 17236 1465 17264 1663
rect 17222 1456 17278 1465
rect 17222 1391 17278 1400
rect 17328 480 17356 6598
rect 17420 6458 17448 6734
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17604 2854 17632 3538
rect 17592 2848 17644 2854
rect 17590 2816 17592 2825
rect 17644 2816 17646 2825
rect 17590 2751 17646 2760
rect 17696 610 17724 20742
rect 19982 20360 20038 20369
rect 19982 20295 20038 20304
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19522 19272 19578 19281
rect 19522 19207 19524 19216
rect 19576 19207 19578 19216
rect 19524 19178 19576 19184
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 17774 13832 17830 13841
rect 17774 13767 17830 13776
rect 17788 6746 17816 13767
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17880 7546 17908 8026
rect 18800 8022 18828 9318
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18892 8634 18920 9114
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18340 7546 18368 7822
rect 18800 7546 18828 7958
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18892 6866 18920 8366
rect 18984 6905 19012 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19996 18834 20024 20295
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19996 18426 20024 18770
rect 20916 18714 20944 26658
rect 23754 25664 23810 25673
rect 23754 25599 23810 25608
rect 23768 24954 23796 25599
rect 21732 24948 21784 24954
rect 21732 24890 21784 24896
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 20994 19000 21050 19009
rect 20994 18935 21050 18944
rect 20824 18686 20944 18714
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19984 10736 20036 10742
rect 19982 10704 19984 10713
rect 20036 10704 20038 10713
rect 19982 10639 20038 10648
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 19076 7750 19104 8434
rect 19260 8430 19288 8978
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19352 8090 19380 8774
rect 19444 8650 19472 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19444 8634 19564 8650
rect 19444 8628 19576 8634
rect 19444 8622 19524 8628
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19444 7886 19472 8622
rect 19524 8570 19576 8576
rect 19904 8362 19932 8910
rect 19892 8356 19944 8362
rect 19944 8316 20024 8344
rect 19892 8298 19944 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 8090 20024 8316
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19076 7206 19104 7686
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18970 6896 19026 6905
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18880 6860 18932 6866
rect 18970 6831 19026 6840
rect 18880 6802 18932 6808
rect 17788 6718 17908 6746
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 5778 17816 6598
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17880 4146 17908 6718
rect 18064 6322 18092 6802
rect 18156 6730 18184 6802
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 18156 5914 18184 6666
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18248 5914 18276 6122
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18340 5710 18368 6190
rect 18892 6118 18920 6802
rect 19076 6662 19104 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19522 6896 19578 6905
rect 19522 6831 19578 6840
rect 19798 6896 19854 6905
rect 19798 6831 19800 6840
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19076 6254 19104 6598
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18602 5808 18658 5817
rect 18602 5743 18604 5752
rect 18656 5743 18658 5752
rect 18604 5714 18656 5720
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18340 5302 18368 5646
rect 18616 5370 18644 5714
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18340 4826 18368 5238
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18156 4078 18184 4762
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18156 3058 18184 4014
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3738 18828 3878
rect 18892 3777 18920 6054
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19260 5681 19288 5782
rect 19246 5672 19302 5681
rect 19246 5607 19302 5616
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19168 4622 19196 4966
rect 19338 4720 19394 4729
rect 19338 4655 19394 4664
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 18878 3768 18934 3777
rect 18788 3732 18840 3738
rect 19168 3738 19196 4558
rect 19352 4554 19380 4655
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 18878 3703 18934 3712
rect 19156 3732 19208 3738
rect 18788 3674 18840 3680
rect 19156 3674 19208 3680
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18602 3632 18658 3641
rect 18248 3194 18276 3606
rect 18602 3567 18658 3576
rect 18696 3596 18748 3602
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18248 2650 18276 3130
rect 18616 2938 18644 3567
rect 18696 3538 18748 3544
rect 18708 3126 18736 3538
rect 18696 3120 18748 3126
rect 18694 3088 18696 3097
rect 18748 3088 18750 3097
rect 18694 3023 18750 3032
rect 18800 2990 18828 3674
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18788 2984 18840 2990
rect 18616 2910 18736 2938
rect 18788 2926 18840 2932
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18432 2281 18460 2450
rect 18604 2304 18656 2310
rect 18418 2272 18474 2281
rect 18604 2246 18656 2252
rect 18418 2207 18474 2216
rect 18616 1465 18644 2246
rect 18602 1456 18658 1465
rect 18602 1391 18658 1400
rect 17684 604 17736 610
rect 17684 546 17736 552
rect 17960 604 18012 610
rect 17960 546 18012 552
rect 17972 480 18000 546
rect 18708 480 18736 2910
rect 18800 2582 18828 2926
rect 18984 2650 19012 2994
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19444 2145 19472 2246
rect 19430 2136 19486 2145
rect 19430 2071 19486 2080
rect 19536 626 19564 6831
rect 19852 6831 19854 6840
rect 19800 6802 19852 6808
rect 19812 6458 19840 6802
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19904 6202 19932 6734
rect 19996 6730 20024 7210
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19996 6458 20024 6666
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19904 6186 20024 6202
rect 19904 6180 20036 6186
rect 19904 6174 19984 6180
rect 19984 6122 20036 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5574 20024 6122
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19614 5400 19670 5409
rect 19614 5335 19616 5344
rect 19668 5335 19670 5344
rect 19616 5306 19668 5312
rect 19720 5098 19748 5510
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 19720 3194 19748 3606
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 20088 2802 20116 18566
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 10736 20404 10742
rect 20352 10678 20404 10684
rect 20166 9616 20222 9625
rect 20166 9551 20222 9560
rect 20180 9178 20208 9551
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20364 9081 20392 10678
rect 20350 9072 20406 9081
rect 20350 9007 20406 9016
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20364 4690 20392 5646
rect 20456 5522 20484 18022
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20732 10538 20760 11018
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20640 10266 20668 10474
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20732 8906 20760 10474
rect 20824 10130 20852 18686
rect 20902 18592 20958 18601
rect 20902 18527 20958 18536
rect 20916 18426 20944 18527
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20916 18222 20944 18362
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 21008 17746 21036 18935
rect 21638 17912 21694 17921
rect 21638 17847 21694 17856
rect 20996 17740 21048 17746
rect 20996 17682 21048 17688
rect 21008 17338 21036 17682
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 9722 20852 10066
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 21192 9194 21220 17478
rect 21652 16658 21680 17847
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21652 16250 21680 16594
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21454 15328 21510 15337
rect 21454 15263 21510 15272
rect 21192 9166 21404 9194
rect 21468 9178 21496 15263
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21560 9382 21588 10066
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 21284 8362 21312 8978
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20548 7546 20576 8026
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 21284 6866 21312 8298
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20456 5494 20760 5522
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 20364 4282 20392 4626
rect 20352 4276 20404 4282
rect 20352 4218 20404 4224
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 19996 2774 20116 2802
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19614 2544 19670 2553
rect 19614 2479 19670 2488
rect 19628 2145 19656 2479
rect 19614 2136 19670 2145
rect 19614 2071 19670 2080
rect 19352 598 19564 626
rect 19996 626 20024 2774
rect 20272 2582 20300 3606
rect 20626 2680 20682 2689
rect 20626 2615 20682 2624
rect 20260 2576 20312 2582
rect 20166 2544 20222 2553
rect 20260 2518 20312 2524
rect 20166 2479 20168 2488
rect 20220 2479 20222 2488
rect 20168 2450 20220 2456
rect 20640 2378 20668 2615
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 19996 598 20116 626
rect 19352 480 19380 598
rect 20088 480 20116 598
rect 20732 480 20760 5494
rect 20824 4826 20852 6598
rect 21284 6118 21312 6802
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20916 5370 20944 5510
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20810 4720 20866 4729
rect 20810 4655 20866 4664
rect 20824 4282 20852 4655
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20916 4146 20944 4558
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 21284 3942 21312 4422
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 21272 3936 21324 3942
rect 21272 3878 21324 3884
rect 20824 3466 20852 3878
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20916 3194 20944 3470
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20916 2650 20944 3130
rect 21192 2854 21220 3538
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21376 480 21404 9166
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21468 8634 21496 9114
rect 21560 8974 21588 9318
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21560 8090 21588 8910
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21744 6866 21772 24890
rect 24122 24304 24178 24313
rect 24122 24239 24178 24248
rect 23754 23624 23810 23633
rect 23754 23559 23810 23568
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23478 16960 23534 16969
rect 23478 16895 23534 16904
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21836 8362 21864 9658
rect 21824 8356 21876 8362
rect 21824 8298 21876 8304
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21652 6338 21680 6734
rect 21744 6458 21772 6802
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21652 6310 21772 6338
rect 21744 6118 21772 6310
rect 21732 6112 21784 6118
rect 21730 6080 21732 6089
rect 21784 6080 21786 6089
rect 21730 6015 21786 6024
rect 21744 5817 21772 6015
rect 21730 5808 21786 5817
rect 21730 5743 21786 5752
rect 21928 4162 21956 16730
rect 23492 15586 23520 16895
rect 23400 15570 23520 15586
rect 23388 15564 23520 15570
rect 23440 15558 23520 15564
rect 23388 15506 23440 15512
rect 23400 15450 23428 15506
rect 23308 15422 23428 15450
rect 23308 15162 23336 15422
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22296 10266 22324 10610
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22466 9072 22522 9081
rect 22466 9007 22468 9016
rect 22520 9007 22522 9016
rect 22468 8978 22520 8984
rect 22480 8634 22508 8978
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22112 5778 22140 8298
rect 22376 5840 22428 5846
rect 22376 5782 22428 5788
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 22112 5409 22140 5714
rect 22098 5400 22154 5409
rect 22098 5335 22100 5344
rect 22152 5335 22154 5344
rect 22100 5306 22152 5312
rect 22112 5275 22140 5306
rect 22388 5098 22416 5782
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 21928 4134 22232 4162
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21560 2582 21588 3334
rect 22020 2650 22048 3878
rect 22112 3233 22140 3878
rect 22098 3224 22154 3233
rect 22098 3159 22154 3168
rect 22204 3074 22232 4134
rect 22112 3046 22232 3074
rect 22480 3058 22508 4966
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22468 3052 22520 3058
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 21548 2576 21600 2582
rect 21548 2518 21600 2524
rect 22006 2408 22062 2417
rect 22006 2343 22062 2352
rect 22020 2009 22048 2343
rect 22006 2000 22062 2009
rect 22006 1935 22062 1944
rect 22112 480 22140 3046
rect 22468 2994 22520 3000
rect 22572 2922 22600 4490
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22572 2689 22600 2858
rect 22558 2680 22614 2689
rect 22558 2615 22614 2624
rect 22664 2281 22692 8910
rect 23110 7032 23166 7041
rect 23110 6967 23166 6976
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22848 4486 22876 4626
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22848 4185 22876 4422
rect 22834 4176 22890 4185
rect 22834 4111 22890 4120
rect 23124 2802 23152 6967
rect 23294 5128 23350 5137
rect 23294 5063 23350 5072
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23216 3942 23244 4558
rect 23308 4146 23336 5063
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23294 3904 23350 3913
rect 23216 3534 23244 3878
rect 23400 3890 23428 15302
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23492 7698 23520 12378
rect 23584 9625 23612 21082
rect 23676 12442 23704 23462
rect 23768 22681 23796 23559
rect 23754 22672 23810 22681
rect 23754 22607 23810 22616
rect 23938 22672 23994 22681
rect 23938 22607 23994 22616
rect 23952 21146 23980 22607
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23938 21040 23994 21049
rect 23938 20975 23994 20984
rect 23846 19816 23902 19825
rect 23846 19751 23902 19760
rect 23860 18601 23888 19751
rect 23952 19281 23980 20975
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 24044 19514 24072 19858
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 23938 19272 23994 19281
rect 23938 19207 23994 19216
rect 23846 18592 23902 18601
rect 23846 18527 23902 18536
rect 24030 17640 24086 17649
rect 24030 17575 24086 17584
rect 24044 15337 24072 17575
rect 24030 15328 24086 15337
rect 24030 15263 24086 15272
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23768 12322 23796 12378
rect 23676 12294 23796 12322
rect 23570 9616 23626 9625
rect 23570 9551 23626 9560
rect 23676 7857 23704 12294
rect 23662 7848 23718 7857
rect 23662 7783 23718 7792
rect 23492 7670 23704 7698
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23492 5370 23520 6734
rect 23570 6080 23626 6089
rect 23570 6015 23626 6024
rect 23584 5914 23612 6015
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23676 5250 23704 7670
rect 23860 6458 23888 13942
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 23952 12442 23980 12854
rect 24044 12442 24072 14758
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24136 12322 24164 24239
rect 24228 13258 24256 26959
rect 24674 26344 24730 26353
rect 24674 26279 24730 26288
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23866 24716 26279
rect 24766 24984 24822 24993
rect 24766 24919 24822 24928
rect 24780 24886 24808 24919
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24688 23662 24716 23802
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24674 21584 24730 21593
rect 24674 21519 24730 21528
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 19922 24716 21519
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24780 19417 24808 19654
rect 24766 19408 24822 19417
rect 24766 19343 24822 19352
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24766 16280 24822 16289
rect 24766 16215 24822 16224
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24780 15162 24808 16215
rect 25226 15192 25282 15201
rect 24768 15156 24820 15162
rect 25226 15127 25282 15136
rect 24768 15098 24820 15104
rect 24858 14920 24914 14929
rect 24858 14855 24914 14864
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24766 13696 24822 13705
rect 24766 13631 24822 13640
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 23952 12294 24164 12322
rect 24214 12336 24270 12345
rect 23952 6905 23980 12294
rect 24596 12322 24624 12582
rect 24688 12442 24716 13126
rect 24780 12646 24808 13631
rect 24872 13394 24900 14855
rect 25240 14074 25268 15127
rect 25318 14376 25374 14385
rect 25318 14311 25374 14320
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25240 13870 25268 14010
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24872 12986 24900 13330
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24596 12306 24716 12322
rect 24596 12300 24728 12306
rect 24596 12294 24676 12300
rect 24214 12271 24270 12280
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 23938 6896 23994 6905
rect 23938 6831 23994 6840
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23768 5370 23796 6190
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23492 5222 23704 5250
rect 23492 4146 23520 5222
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23584 4078 23612 4626
rect 23572 4072 23624 4078
rect 23478 4040 23534 4049
rect 23572 4014 23624 4020
rect 23478 3975 23480 3984
rect 23532 3975 23534 3984
rect 23480 3946 23532 3952
rect 23400 3862 23520 3890
rect 23294 3839 23350 3848
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23216 3126 23244 3470
rect 23308 3194 23336 3839
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23204 3120 23256 3126
rect 23204 3062 23256 3068
rect 23216 2990 23244 3062
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23204 2984 23256 2990
rect 23204 2926 23256 2932
rect 23124 2774 23244 2802
rect 22650 2272 22706 2281
rect 22650 2207 22706 2216
rect 23216 1873 23244 2774
rect 23400 2650 23428 2994
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23202 1864 23258 1873
rect 23202 1799 23258 1808
rect 22742 1456 22798 1465
rect 22742 1391 22798 1400
rect 22756 480 22784 1391
rect 23492 480 23520 3862
rect 23584 3738 23612 4014
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23570 3632 23626 3641
rect 23570 3567 23626 3576
rect 23584 2145 23612 3567
rect 23676 2961 23704 4762
rect 23768 4282 23796 4966
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23768 4049 23796 4082
rect 23754 4040 23810 4049
rect 23754 3975 23810 3984
rect 23756 3596 23808 3602
rect 23756 3538 23808 3544
rect 23662 2952 23718 2961
rect 23768 2922 23796 3538
rect 23860 3398 23888 6258
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23952 3670 23980 3878
rect 23940 3664 23992 3670
rect 23940 3606 23992 3612
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 24044 2972 24072 12174
rect 24136 7449 24164 12174
rect 24228 10577 24256 12271
rect 24676 12242 24728 12248
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12242
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24780 11778 24808 12038
rect 24780 11750 24900 11778
rect 24766 11656 24822 11665
rect 24766 11591 24822 11600
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24214 10568 24270 10577
rect 24214 10503 24270 10512
rect 24214 10296 24270 10305
rect 24214 10231 24270 10240
rect 24228 8945 24256 10231
rect 24780 10033 24808 11591
rect 24872 10849 24900 11750
rect 24950 10976 25006 10985
rect 24950 10911 25006 10920
rect 24858 10840 24914 10849
rect 24858 10775 24914 10784
rect 24766 10024 24822 10033
rect 24766 9959 24822 9968
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24964 9738 24992 10911
rect 24780 9710 24992 9738
rect 24780 9704 24808 9710
rect 24688 9676 24808 9704
rect 24688 9489 24716 9676
rect 24674 9480 24730 9489
rect 24674 9415 24730 9424
rect 24214 8936 24270 8945
rect 24214 8871 24270 8880
rect 24674 8936 24730 8945
rect 24674 8871 24730 8880
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24122 7440 24178 7449
rect 24122 7375 24178 7384
rect 24688 7313 24716 8871
rect 24766 8256 24822 8265
rect 24766 8191 24822 8200
rect 24674 7304 24730 7313
rect 24674 7239 24730 7248
rect 24214 7168 24270 7177
rect 24214 7103 24270 7112
rect 24228 5914 24256 7103
rect 24780 7002 24808 8191
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6458 24716 6802
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24766 6352 24822 6361
rect 24766 6287 24822 6296
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24216 5636 24268 5642
rect 24216 5578 24268 5584
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24136 5370 24164 5510
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 24228 4978 24256 5578
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24308 5092 24360 5098
rect 24308 5034 24360 5040
rect 24136 4950 24256 4978
rect 24136 3074 24164 4950
rect 24214 4856 24270 4865
rect 24320 4826 24348 5034
rect 24688 5030 24716 5714
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24214 4791 24270 4800
rect 24308 4820 24360 4826
rect 24228 3505 24256 4791
rect 24308 4762 24360 4768
rect 24688 4729 24716 4966
rect 24674 4720 24730 4729
rect 24674 4655 24730 4664
rect 24780 4593 24808 6287
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24766 4584 24822 4593
rect 24766 4519 24822 4528
rect 24872 4434 24900 6054
rect 24964 5846 24992 6190
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24688 4406 24900 4434
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24214 3496 24270 3505
rect 24214 3431 24270 3440
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24136 3046 24532 3074
rect 24044 2944 24164 2972
rect 23662 2887 23718 2896
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 23662 2544 23718 2553
rect 23662 2479 23718 2488
rect 23570 2136 23626 2145
rect 23570 2071 23626 2080
rect 23676 1601 23704 2479
rect 23768 2310 23796 2858
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23860 2650 23888 2790
rect 23938 2680 23994 2689
rect 23848 2644 23900 2650
rect 23938 2615 23994 2624
rect 23848 2586 23900 2592
rect 23952 2582 23980 2615
rect 23940 2576 23992 2582
rect 23940 2518 23992 2524
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 23662 1592 23718 1601
rect 23662 1527 23718 1536
rect 24136 480 24164 2944
rect 24504 2553 24532 3046
rect 24490 2544 24546 2553
rect 24490 2479 24546 2488
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1601 24716 4406
rect 24766 4312 24822 4321
rect 25056 4282 25084 13194
rect 25332 12986 25360 14311
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 26882 10840 26938 10849
rect 26882 10775 26938 10784
rect 25134 9616 25190 9625
rect 25134 9551 25190 9560
rect 24766 4247 24822 4256
rect 25044 4276 25096 4282
rect 24780 3097 24808 4247
rect 25044 4218 25096 4224
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24872 3738 24900 4014
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24766 3088 24822 3097
rect 24766 3023 24822 3032
rect 24872 2972 24900 3334
rect 24780 2944 24900 2972
rect 24674 1592 24730 1601
rect 24674 1527 24730 1536
rect 24780 480 24808 2944
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25056 2582 25084 2790
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 25148 1737 25176 9551
rect 26146 7848 26202 7857
rect 26146 7783 26202 7792
rect 25502 7440 25558 7449
rect 25502 7375 25558 7384
rect 25228 5160 25280 5166
rect 25226 5128 25228 5137
rect 25280 5128 25282 5137
rect 25226 5063 25282 5072
rect 25410 4176 25466 4185
rect 25410 4111 25412 4120
rect 25464 4111 25466 4120
rect 25412 4082 25464 4088
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25240 3913 25268 4014
rect 25226 3904 25282 3913
rect 25226 3839 25282 3848
rect 25134 1728 25190 1737
rect 25134 1663 25190 1672
rect 25516 480 25544 7375
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2318 0 2374 480
rect 2962 0 3018 480
rect 3698 0 3754 480
rect 4342 0 4398 480
rect 4986 0 5042 480
rect 5722 0 5778 480
rect 6366 0 6422 480
rect 7102 0 7158 480
rect 7746 0 7802 480
rect 8390 0 8446 480
rect 9126 0 9182 480
rect 9770 0 9826 480
rect 10506 0 10562 480
rect 11150 0 11206 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13174 0 13230 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15290 0 15346 480
rect 15934 0 15990 480
rect 16578 0 16634 480
rect 17314 0 17370 480
rect 17958 0 18014 480
rect 18694 0 18750 480
rect 19338 0 19394 480
rect 20074 0 20130 480
rect 20718 0 20774 480
rect 21362 0 21418 480
rect 22098 0 22154 480
rect 22742 0 22798 480
rect 23478 0 23534 480
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25502 0 25558 480
rect 25700 377 25728 4966
rect 26160 480 26188 7783
rect 26896 480 26924 10775
rect 27526 4040 27582 4049
rect 27526 3975 27582 3984
rect 27540 480 27568 3975
rect 25686 368 25742 377
rect 25686 303 25742 312
rect 26146 0 26202 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 24122 27648 24178 27704
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 13818 12688 13874 12744
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 1582 10512 1638 10568
rect 1582 9988 1638 10024
rect 1582 9968 1584 9988
rect 1584 9968 1636 9988
rect 1636 9968 1638 9988
rect 294 3032 350 3088
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 2226 9424 2282 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 2870 8900 2926 8936
rect 2870 8880 2872 8900
rect 2872 8880 2924 8900
rect 2924 8880 2926 8900
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 4250 7248 4306 7304
rect 4250 1400 4306 1456
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 7654 5752 7710 5808
rect 9678 5788 9680 5808
rect 9680 5788 9732 5808
rect 9732 5788 9734 5808
rect 9678 5752 9734 5788
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 7010 4548 7066 4584
rect 7010 4528 7012 4548
rect 7012 4528 7064 4548
rect 7064 4528 7066 4548
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 4986 3984 5042 4040
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6826 1536 6882 1592
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 8298 3460 8354 3496
rect 8298 3440 8300 3460
rect 8300 3440 8352 3460
rect 8352 3440 8354 3460
rect 11886 3032 11942 3088
rect 9034 2896 9090 2952
rect 8206 1808 8262 1864
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11058 2488 11114 2544
rect 9954 2080 10010 2136
rect 10506 1672 10562 1728
rect 13174 2760 13230 2816
rect 12806 992 12862 1048
rect 24214 26968 24270 27024
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 14278 10648 14334 10704
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 16118 22616 16174 22672
rect 17498 22480 17554 22536
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15290 4684 15346 4720
rect 15290 4664 15292 4684
rect 15292 4664 15344 4684
rect 15344 4664 15346 4684
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14462 2488 14518 2544
rect 14462 1944 14518 2000
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14738 2488 14794 2544
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14738 2080 14794 2136
rect 16486 3188 16542 3224
rect 16486 3168 16488 3188
rect 16488 3168 16540 3188
rect 16540 3168 16542 3188
rect 16118 2252 16120 2272
rect 16120 2252 16172 2272
rect 16172 2252 16174 2272
rect 16118 2216 16174 2252
rect 17038 2080 17094 2136
rect 17038 1672 17094 1728
rect 17222 1672 17278 1728
rect 17222 1400 17278 1456
rect 17590 2796 17592 2816
rect 17592 2796 17644 2816
rect 17644 2796 17646 2816
rect 17590 2760 17646 2796
rect 19982 20304 20038 20360
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19522 19236 19578 19272
rect 19522 19216 19524 19236
rect 19524 19216 19576 19236
rect 19576 19216 19578 19236
rect 17774 13776 17830 13832
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 23754 25608 23810 25664
rect 20994 18944 21050 19000
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19982 10684 19984 10704
rect 19984 10684 20036 10704
rect 20036 10684 20038 10704
rect 19982 10648 20038 10684
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 18970 6840 19026 6896
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19522 6840 19578 6896
rect 19798 6860 19854 6896
rect 19798 6840 19800 6860
rect 19800 6840 19852 6860
rect 19852 6840 19854 6860
rect 18602 5772 18658 5808
rect 18602 5752 18604 5772
rect 18604 5752 18656 5772
rect 18656 5752 18658 5772
rect 19246 5616 19302 5672
rect 19338 4664 19394 4720
rect 18878 3712 18934 3768
rect 18602 3576 18658 3632
rect 18694 3068 18696 3088
rect 18696 3068 18748 3088
rect 18748 3068 18750 3088
rect 18694 3032 18750 3068
rect 18418 2216 18474 2272
rect 18602 1400 18658 1456
rect 19430 2080 19486 2136
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19614 5364 19670 5400
rect 19614 5344 19616 5364
rect 19616 5344 19668 5364
rect 19668 5344 19670 5364
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20166 9560 20222 9616
rect 20350 9016 20406 9072
rect 20902 18536 20958 18592
rect 21638 17856 21694 17912
rect 21454 15272 21510 15328
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19614 2488 19670 2544
rect 19614 2080 19670 2136
rect 20626 2624 20682 2680
rect 20166 2508 20222 2544
rect 20166 2488 20168 2508
rect 20168 2488 20220 2508
rect 20220 2488 20222 2508
rect 20810 4664 20866 4720
rect 24122 24248 24178 24304
rect 23754 23568 23810 23624
rect 23478 16904 23534 16960
rect 21730 6060 21732 6080
rect 21732 6060 21784 6080
rect 21784 6060 21786 6080
rect 21730 6024 21786 6060
rect 21730 5752 21786 5808
rect 22466 9036 22522 9072
rect 22466 9016 22468 9036
rect 22468 9016 22520 9036
rect 22520 9016 22522 9036
rect 22098 5364 22154 5400
rect 22098 5344 22100 5364
rect 22100 5344 22152 5364
rect 22152 5344 22154 5364
rect 22098 3168 22154 3224
rect 22006 2352 22062 2408
rect 22006 1944 22062 2000
rect 22558 2624 22614 2680
rect 23110 6976 23166 7032
rect 22834 4120 22890 4176
rect 23294 5072 23350 5128
rect 23294 3848 23350 3904
rect 23754 22616 23810 22672
rect 23938 22616 23994 22672
rect 23938 20984 23994 21040
rect 23846 19760 23902 19816
rect 23938 19216 23994 19272
rect 23846 18536 23902 18592
rect 24030 17584 24086 17640
rect 24030 15272 24086 15328
rect 23570 9560 23626 9616
rect 23662 7792 23718 7848
rect 23570 6024 23626 6080
rect 24674 26288 24730 26344
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 24928 24822 24984
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24674 21528 24730 21584
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 19352 24822 19408
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24766 16224 24822 16280
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 25226 15136 25282 15192
rect 24858 14864 24914 14920
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13640 24822 13696
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24214 12280 24270 12336
rect 25318 14320 25374 14376
rect 23938 6840 23994 6896
rect 23478 4004 23534 4040
rect 23478 3984 23480 4004
rect 23480 3984 23532 4004
rect 23532 3984 23534 4004
rect 22650 2216 22706 2272
rect 23202 1808 23258 1864
rect 22742 1400 22798 1456
rect 23570 3576 23626 3632
rect 23754 3984 23810 4040
rect 23662 2896 23718 2952
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11600 24822 11656
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24214 10512 24270 10568
rect 24214 10240 24270 10296
rect 24950 10920 25006 10976
rect 24858 10784 24914 10840
rect 24766 9968 24822 10024
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 9424 24730 9480
rect 24214 8880 24270 8936
rect 24674 8880 24730 8936
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24122 7384 24178 7440
rect 24766 8200 24822 8256
rect 24674 7248 24730 7304
rect 24214 7112 24270 7168
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24766 6296 24822 6352
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24214 4800 24270 4856
rect 24674 4664 24730 4720
rect 24766 4528 24822 4584
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24214 3440 24270 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23662 2488 23718 2544
rect 23570 2080 23626 2136
rect 23938 2624 23994 2680
rect 23662 1536 23718 1592
rect 24490 2488 24546 2544
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24766 4256 24822 4312
rect 26882 10784 26938 10840
rect 25134 9560 25190 9616
rect 24766 3032 24822 3088
rect 24674 1536 24730 1592
rect 26146 7792 26202 7848
rect 25502 7384 25558 7440
rect 25226 5108 25228 5128
rect 25228 5108 25280 5128
rect 25280 5108 25282 5128
rect 25226 5072 25282 5108
rect 25410 4140 25466 4176
rect 25410 4120 25412 4140
rect 25412 4120 25464 4140
rect 25464 4120 25466 4140
rect 25226 3848 25282 3904
rect 25134 1672 25190 1728
rect 27526 3984 27582 4040
rect 25686 312 25742 368
<< metal3 >>
rect 24117 27706 24183 27709
rect 27520 27706 28000 27736
rect 24117 27704 28000 27706
rect 24117 27648 24122 27704
rect 24178 27648 28000 27704
rect 24117 27646 28000 27648
rect 24117 27643 24183 27646
rect 27520 27616 28000 27646
rect 24209 27026 24275 27029
rect 27520 27026 28000 27056
rect 24209 27024 28000 27026
rect 24209 26968 24214 27024
rect 24270 26968 28000 27024
rect 24209 26966 28000 26968
rect 24209 26963 24275 26966
rect 27520 26936 28000 26966
rect 24669 26346 24735 26349
rect 27520 26346 28000 26376
rect 24669 26344 28000 26346
rect 24669 26288 24674 26344
rect 24730 26288 28000 26344
rect 24669 26286 28000 26288
rect 24669 26283 24735 26286
rect 27520 26256 28000 26286
rect 23749 25666 23815 25669
rect 27520 25666 28000 25696
rect 23749 25664 28000 25666
rect 23749 25608 23754 25664
rect 23810 25608 28000 25664
rect 23749 25606 28000 25608
rect 23749 25603 23815 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 27520 25576 28000 25606
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 24761 24986 24827 24989
rect 27520 24986 28000 25016
rect 24761 24984 28000 24986
rect 24761 24928 24766 24984
rect 24822 24928 28000 24984
rect 24761 24926 28000 24928
rect 24761 24923 24827 24926
rect 27520 24896 28000 24926
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 24117 24306 24183 24309
rect 27520 24306 28000 24336
rect 24117 24304 28000 24306
rect 24117 24248 24122 24304
rect 24178 24248 28000 24304
rect 24117 24246 28000 24248
rect 24117 24243 24183 24246
rect 27520 24216 28000 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 23749 23626 23815 23629
rect 27520 23626 28000 23656
rect 23749 23624 28000 23626
rect 23749 23568 23754 23624
rect 23810 23568 28000 23624
rect 23749 23566 28000 23568
rect 23749 23563 23815 23566
rect 27520 23536 28000 23566
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 27520 22946 28000 22976
rect 24718 22886 28000 22946
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 16113 22674 16179 22677
rect 23749 22674 23815 22677
rect 16113 22672 23815 22674
rect 16113 22616 16118 22672
rect 16174 22616 23754 22672
rect 23810 22616 23815 22672
rect 16113 22614 23815 22616
rect 16113 22611 16179 22614
rect 23749 22611 23815 22614
rect 23933 22674 23999 22677
rect 24718 22674 24778 22886
rect 27520 22856 28000 22886
rect 23933 22672 24778 22674
rect 23933 22616 23938 22672
rect 23994 22616 24778 22672
rect 23933 22614 24778 22616
rect 23933 22611 23999 22614
rect 17493 22538 17559 22541
rect 17493 22536 24962 22538
rect 17493 22480 17498 22536
rect 17554 22480 24962 22536
rect 17493 22478 24962 22480
rect 17493 22475 17559 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 24902 22266 24962 22478
rect 27520 22266 28000 22296
rect 24902 22206 28000 22266
rect 27520 22176 28000 22206
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 24669 21586 24735 21589
rect 27520 21586 28000 21616
rect 24669 21584 28000 21586
rect 24669 21528 24674 21584
rect 24730 21528 28000 21584
rect 24669 21526 28000 21528
rect 24669 21523 24735 21526
rect 27520 21496 28000 21526
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 23933 21042 23999 21045
rect 27520 21042 28000 21072
rect 23933 21040 28000 21042
rect 23933 20984 23938 21040
rect 23994 20984 28000 21040
rect 23933 20982 28000 20984
rect 23933 20979 23999 20982
rect 27520 20952 28000 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 19977 20362 20043 20365
rect 27520 20362 28000 20392
rect 19977 20360 28000 20362
rect 19977 20304 19982 20360
rect 20038 20304 28000 20360
rect 19977 20302 28000 20304
rect 19977 20299 20043 20302
rect 27520 20272 28000 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 23841 19818 23907 19821
rect 23841 19816 24778 19818
rect 23841 19760 23846 19816
rect 23902 19760 24778 19816
rect 23841 19758 24778 19760
rect 23841 19755 23907 19758
rect 24718 19682 24778 19758
rect 27520 19682 28000 19712
rect 24718 19622 28000 19682
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19622
rect 24277 19551 24597 19552
rect 24761 19412 24827 19413
rect 24710 19410 24716 19412
rect 24670 19350 24716 19410
rect 24780 19408 24827 19412
rect 24822 19352 24827 19408
rect 24710 19348 24716 19350
rect 24780 19348 24827 19352
rect 24761 19347 24827 19348
rect 19517 19274 19583 19277
rect 23933 19274 23999 19277
rect 19517 19272 23999 19274
rect 19517 19216 19522 19272
rect 19578 19216 23938 19272
rect 23994 19216 23999 19272
rect 19517 19214 23999 19216
rect 19517 19211 19583 19214
rect 23933 19211 23999 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 20989 19002 21055 19005
rect 27520 19002 28000 19032
rect 20989 19000 28000 19002
rect 20989 18944 20994 19000
rect 21050 18944 28000 19000
rect 20989 18942 28000 18944
rect 20989 18939 21055 18942
rect 27520 18912 28000 18942
rect 20897 18594 20963 18597
rect 23841 18594 23907 18597
rect 20897 18592 23907 18594
rect 20897 18536 20902 18592
rect 20958 18536 23846 18592
rect 23902 18536 23907 18592
rect 20897 18534 23907 18536
rect 20897 18531 20963 18534
rect 23841 18531 23907 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 27520 18322 28000 18352
rect 24718 18262 28000 18322
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 21633 17914 21699 17917
rect 24718 17914 24778 18262
rect 27520 18232 28000 18262
rect 21633 17912 24778 17914
rect 21633 17856 21638 17912
rect 21694 17856 24778 17912
rect 21633 17854 24778 17856
rect 21633 17851 21699 17854
rect 24025 17642 24091 17645
rect 27520 17642 28000 17672
rect 24025 17640 28000 17642
rect 24025 17584 24030 17640
rect 24086 17584 28000 17640
rect 24025 17582 28000 17584
rect 24025 17579 24091 17582
rect 27520 17552 28000 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 23473 16962 23539 16965
rect 27520 16962 28000 16992
rect 23473 16960 28000 16962
rect 23473 16904 23478 16960
rect 23534 16904 28000 16960
rect 23473 16902 28000 16904
rect 23473 16899 23539 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 27520 16872 28000 16902
rect 19610 16831 19930 16832
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 24761 16282 24827 16285
rect 27520 16282 28000 16312
rect 24761 16280 28000 16282
rect 24761 16224 24766 16280
rect 24822 16224 28000 16280
rect 24761 16222 28000 16224
rect 24761 16219 24827 16222
rect 27520 16192 28000 16222
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 27520 15602 28000 15632
rect 25270 15542 28000 15602
rect 21449 15330 21515 15333
rect 24025 15330 24091 15333
rect 21449 15328 24091 15330
rect 21449 15272 21454 15328
rect 21510 15272 24030 15328
rect 24086 15272 24091 15328
rect 21449 15270 24091 15272
rect 21449 15267 21515 15270
rect 24025 15267 24091 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 25270 15197 25330 15542
rect 27520 15512 28000 15542
rect 25221 15192 25330 15197
rect 25221 15136 25226 15192
rect 25282 15136 25330 15192
rect 25221 15134 25330 15136
rect 25221 15131 25287 15134
rect 24853 14922 24919 14925
rect 27520 14922 28000 14952
rect 24853 14920 28000 14922
rect 24853 14864 24858 14920
rect 24914 14864 28000 14920
rect 24853 14862 28000 14864
rect 24853 14859 24919 14862
rect 27520 14832 28000 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 25313 14378 25379 14381
rect 27520 14378 28000 14408
rect 25313 14376 28000 14378
rect 25313 14320 25318 14376
rect 25374 14320 28000 14376
rect 25313 14318 28000 14320
rect 25313 14315 25379 14318
rect 27520 14288 28000 14318
rect 5610 14176 5930 14177
rect 0 14106 480 14136
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 14046 3618 14106
rect 0 14016 480 14046
rect 3558 13834 3618 14046
rect 17769 13834 17835 13837
rect 3558 13832 17835 13834
rect 3558 13776 17774 13832
rect 17830 13776 17835 13832
rect 3558 13774 17835 13776
rect 17769 13771 17835 13774
rect 24761 13698 24827 13701
rect 27520 13698 28000 13728
rect 24761 13696 28000 13698
rect 24761 13640 24766 13696
rect 24822 13640 28000 13696
rect 24761 13638 28000 13640
rect 24761 13635 24827 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 27520 13018 28000 13048
rect 24902 12958 28000 13018
rect 13813 12746 13879 12749
rect 24902 12746 24962 12958
rect 27520 12928 28000 12958
rect 13813 12744 24962 12746
rect 13813 12688 13818 12744
rect 13874 12688 24962 12744
rect 13813 12686 24962 12688
rect 13813 12683 13879 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 24209 12338 24275 12341
rect 27520 12338 28000 12368
rect 24209 12336 28000 12338
rect 24209 12280 24214 12336
rect 24270 12280 28000 12336
rect 24209 12278 28000 12280
rect 24209 12275 24275 12278
rect 27520 12248 28000 12278
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 24761 11658 24827 11661
rect 27520 11658 28000 11688
rect 24761 11656 28000 11658
rect 24761 11600 24766 11656
rect 24822 11600 28000 11656
rect 24761 11598 28000 11600
rect 24761 11595 24827 11598
rect 27520 11568 28000 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 24945 10978 25011 10981
rect 27520 10978 28000 11008
rect 24945 10976 28000 10978
rect 24945 10920 24950 10976
rect 25006 10920 28000 10976
rect 24945 10918 28000 10920
rect 24945 10915 25011 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 27520 10888 28000 10918
rect 24277 10847 24597 10848
rect 24853 10842 24919 10845
rect 26877 10842 26943 10845
rect 24853 10840 26943 10842
rect 24853 10784 24858 10840
rect 24914 10784 26882 10840
rect 26938 10784 26943 10840
rect 24853 10782 26943 10784
rect 24853 10779 24919 10782
rect 26877 10779 26943 10782
rect 14273 10706 14339 10709
rect 19977 10706 20043 10709
rect 14273 10704 20043 10706
rect 14273 10648 14278 10704
rect 14334 10648 19982 10704
rect 20038 10648 20043 10704
rect 14273 10646 20043 10648
rect 14273 10643 14339 10646
rect 19977 10643 20043 10646
rect 1577 10570 1643 10573
rect 24209 10570 24275 10573
rect 1577 10568 24275 10570
rect 1577 10512 1582 10568
rect 1638 10512 24214 10568
rect 24270 10512 24275 10568
rect 1577 10510 24275 10512
rect 1577 10507 1643 10510
rect 24209 10507 24275 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 24209 10298 24275 10301
rect 27520 10298 28000 10328
rect 24209 10296 28000 10298
rect 24209 10240 24214 10296
rect 24270 10240 28000 10296
rect 24209 10238 28000 10240
rect 24209 10235 24275 10238
rect 27520 10208 28000 10238
rect 1577 10026 1643 10029
rect 24761 10026 24827 10029
rect 1577 10024 24827 10026
rect 1577 9968 1582 10024
rect 1638 9968 24766 10024
rect 24822 9968 24827 10024
rect 1577 9966 24827 9968
rect 1577 9963 1643 9966
rect 24761 9963 24827 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 20161 9618 20227 9621
rect 23565 9618 23631 9621
rect 20161 9616 23631 9618
rect 20161 9560 20166 9616
rect 20222 9560 23570 9616
rect 23626 9560 23631 9616
rect 20161 9558 23631 9560
rect 20161 9555 20227 9558
rect 23565 9555 23631 9558
rect 25129 9618 25195 9621
rect 27520 9618 28000 9648
rect 25129 9616 28000 9618
rect 25129 9560 25134 9616
rect 25190 9560 28000 9616
rect 25129 9558 28000 9560
rect 25129 9555 25195 9558
rect 27520 9528 28000 9558
rect 2221 9482 2287 9485
rect 24669 9482 24735 9485
rect 2221 9480 24735 9482
rect 2221 9424 2226 9480
rect 2282 9424 24674 9480
rect 24730 9424 24735 9480
rect 2221 9422 24735 9424
rect 2221 9419 2287 9422
rect 24669 9419 24735 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 20345 9074 20411 9077
rect 22461 9074 22527 9077
rect 20345 9072 22527 9074
rect 20345 9016 20350 9072
rect 20406 9016 22466 9072
rect 22522 9016 22527 9072
rect 20345 9014 22527 9016
rect 20345 9011 20411 9014
rect 22461 9011 22527 9014
rect 2865 8938 2931 8941
rect 24209 8938 24275 8941
rect 2865 8936 24275 8938
rect 2865 8880 2870 8936
rect 2926 8880 24214 8936
rect 24270 8880 24275 8936
rect 2865 8878 24275 8880
rect 2865 8875 2931 8878
rect 24209 8875 24275 8878
rect 24669 8938 24735 8941
rect 27520 8938 28000 8968
rect 24669 8936 28000 8938
rect 24669 8880 24674 8936
rect 24730 8880 28000 8936
rect 24669 8878 28000 8880
rect 24669 8875 24735 8878
rect 27520 8848 28000 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 24761 8258 24827 8261
rect 27520 8258 28000 8288
rect 24761 8256 28000 8258
rect 24761 8200 24766 8256
rect 24822 8200 28000 8256
rect 24761 8198 28000 8200
rect 24761 8195 24827 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 23657 7850 23723 7853
rect 26141 7850 26207 7853
rect 23657 7848 26207 7850
rect 23657 7792 23662 7848
rect 23718 7792 26146 7848
rect 26202 7792 26207 7848
rect 23657 7790 26207 7792
rect 23657 7787 23723 7790
rect 26141 7787 26207 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27520 7578 28000 7608
rect 25638 7518 28000 7578
rect 24117 7442 24183 7445
rect 25497 7442 25563 7445
rect 24117 7440 25563 7442
rect 24117 7384 24122 7440
rect 24178 7384 25502 7440
rect 25558 7384 25563 7440
rect 24117 7382 25563 7384
rect 24117 7379 24183 7382
rect 25497 7379 25563 7382
rect 4245 7306 4311 7309
rect 24669 7306 24735 7309
rect 4245 7304 24735 7306
rect 4245 7248 4250 7304
rect 4306 7248 24674 7304
rect 24730 7248 24735 7304
rect 4245 7246 24735 7248
rect 4245 7243 4311 7246
rect 24669 7243 24735 7246
rect 24209 7170 24275 7173
rect 25638 7170 25698 7518
rect 27520 7488 28000 7518
rect 24209 7168 25698 7170
rect 24209 7112 24214 7168
rect 24270 7112 25698 7168
rect 24209 7110 25698 7112
rect 24209 7107 24275 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 23105 7034 23171 7037
rect 27520 7034 28000 7064
rect 23105 7032 28000 7034
rect 23105 6976 23110 7032
rect 23166 6976 28000 7032
rect 23105 6974 28000 6976
rect 23105 6971 23171 6974
rect 27520 6944 28000 6974
rect 18965 6898 19031 6901
rect 19517 6898 19583 6901
rect 18965 6896 19583 6898
rect 18965 6840 18970 6896
rect 19026 6840 19522 6896
rect 19578 6840 19583 6896
rect 18965 6838 19583 6840
rect 18965 6835 19031 6838
rect 19517 6835 19583 6838
rect 19793 6898 19859 6901
rect 23933 6898 23999 6901
rect 19793 6896 23999 6898
rect 19793 6840 19798 6896
rect 19854 6840 23938 6896
rect 23994 6840 23999 6896
rect 19793 6838 23999 6840
rect 19793 6835 19859 6838
rect 23933 6835 23999 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 24761 6354 24827 6357
rect 27520 6354 28000 6384
rect 24761 6352 28000 6354
rect 24761 6296 24766 6352
rect 24822 6296 28000 6352
rect 24761 6294 28000 6296
rect 24761 6291 24827 6294
rect 27520 6264 28000 6294
rect 21725 6082 21791 6085
rect 23565 6082 23631 6085
rect 21725 6080 23631 6082
rect 21725 6024 21730 6080
rect 21786 6024 23570 6080
rect 23626 6024 23631 6080
rect 21725 6022 23631 6024
rect 21725 6019 21791 6022
rect 23565 6019 23631 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 7649 5810 7715 5813
rect 9673 5810 9739 5813
rect 7649 5808 9739 5810
rect 7649 5752 7654 5808
rect 7710 5752 9678 5808
rect 9734 5752 9739 5808
rect 7649 5750 9739 5752
rect 7649 5747 7715 5750
rect 9673 5747 9739 5750
rect 18597 5810 18663 5813
rect 21725 5810 21791 5813
rect 18597 5808 21791 5810
rect 18597 5752 18602 5808
rect 18658 5752 21730 5808
rect 21786 5752 21791 5808
rect 18597 5750 21791 5752
rect 18597 5747 18663 5750
rect 21725 5747 21791 5750
rect 19241 5674 19307 5677
rect 27520 5674 28000 5704
rect 19241 5672 28000 5674
rect 19241 5616 19246 5672
rect 19302 5616 28000 5672
rect 19241 5614 28000 5616
rect 19241 5611 19307 5614
rect 27520 5584 28000 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 19609 5402 19675 5405
rect 22093 5402 22159 5405
rect 19609 5400 22159 5402
rect 19609 5344 19614 5400
rect 19670 5344 22098 5400
rect 22154 5344 22159 5400
rect 19609 5342 22159 5344
rect 19609 5339 19675 5342
rect 22093 5339 22159 5342
rect 23289 5130 23355 5133
rect 25221 5130 25287 5133
rect 23289 5128 25287 5130
rect 23289 5072 23294 5128
rect 23350 5072 25226 5128
rect 25282 5072 25287 5128
rect 23289 5070 25287 5072
rect 23289 5067 23355 5070
rect 25221 5067 25287 5070
rect 27520 4994 28000 5024
rect 24350 4934 28000 4994
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 24209 4858 24275 4861
rect 24350 4858 24410 4934
rect 27520 4904 28000 4934
rect 24209 4856 24410 4858
rect 24209 4800 24214 4856
rect 24270 4800 24410 4856
rect 24209 4798 24410 4800
rect 24209 4795 24275 4798
rect 15285 4722 15351 4725
rect 19333 4722 19399 4725
rect 15285 4720 19399 4722
rect 15285 4664 15290 4720
rect 15346 4664 19338 4720
rect 19394 4664 19399 4720
rect 15285 4662 19399 4664
rect 15285 4659 15351 4662
rect 19333 4659 19399 4662
rect 20805 4722 20871 4725
rect 24669 4722 24735 4725
rect 20805 4720 24735 4722
rect 20805 4664 20810 4720
rect 20866 4664 24674 4720
rect 24730 4664 24735 4720
rect 20805 4662 24735 4664
rect 20805 4659 20871 4662
rect 24669 4659 24735 4662
rect 7005 4586 7071 4589
rect 24761 4586 24827 4589
rect 7005 4584 24827 4586
rect 7005 4528 7010 4584
rect 7066 4528 24766 4584
rect 24822 4528 24827 4584
rect 7005 4526 24827 4528
rect 7005 4523 7071 4526
rect 24761 4523 24827 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 24761 4314 24827 4317
rect 27520 4314 28000 4344
rect 24761 4312 28000 4314
rect 24761 4256 24766 4312
rect 24822 4256 28000 4312
rect 24761 4254 28000 4256
rect 24761 4251 24827 4254
rect 27520 4224 28000 4254
rect 22829 4178 22895 4181
rect 25405 4178 25471 4181
rect 22829 4176 25471 4178
rect 22829 4120 22834 4176
rect 22890 4120 25410 4176
rect 25466 4120 25471 4176
rect 22829 4118 25471 4120
rect 22829 4115 22895 4118
rect 25405 4115 25471 4118
rect 4981 4042 5047 4045
rect 23473 4042 23539 4045
rect 4981 4040 23539 4042
rect 4981 3984 4986 4040
rect 5042 3984 23478 4040
rect 23534 3984 23539 4040
rect 4981 3982 23539 3984
rect 4981 3979 5047 3982
rect 23473 3979 23539 3982
rect 23749 4042 23815 4045
rect 27521 4042 27587 4045
rect 23749 4040 27587 4042
rect 23749 3984 23754 4040
rect 23810 3984 27526 4040
rect 27582 3984 27587 4040
rect 23749 3982 27587 3984
rect 23749 3979 23815 3982
rect 27521 3979 27587 3982
rect 23289 3906 23355 3909
rect 25221 3906 25287 3909
rect 23289 3904 25287 3906
rect 23289 3848 23294 3904
rect 23350 3848 25226 3904
rect 25282 3848 25287 3904
rect 23289 3846 25287 3848
rect 23289 3843 23355 3846
rect 25221 3843 25287 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 18873 3770 18939 3773
rect 24710 3770 24716 3772
rect 10734 3768 18939 3770
rect 10734 3712 18878 3768
rect 18934 3712 18939 3768
rect 10734 3710 18939 3712
rect 10734 3634 10794 3710
rect 18873 3707 18939 3710
rect 20164 3710 24716 3770
rect 7606 3574 10794 3634
rect 18597 3634 18663 3637
rect 20164 3634 20224 3710
rect 24710 3708 24716 3710
rect 24780 3708 24786 3772
rect 18597 3632 20224 3634
rect 18597 3576 18602 3632
rect 18658 3576 20224 3632
rect 18597 3574 20224 3576
rect 23565 3634 23631 3637
rect 27520 3634 28000 3664
rect 23565 3632 28000 3634
rect 23565 3576 23570 3632
rect 23626 3576 28000 3632
rect 23565 3574 28000 3576
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 289 3090 355 3093
rect 7606 3090 7666 3574
rect 18597 3571 18663 3574
rect 23565 3571 23631 3574
rect 27520 3544 28000 3574
rect 8293 3498 8359 3501
rect 24209 3498 24275 3501
rect 8293 3496 24275 3498
rect 8293 3440 8298 3496
rect 8354 3440 24214 3496
rect 24270 3440 24275 3496
rect 8293 3438 24275 3440
rect 8293 3435 8359 3438
rect 24209 3435 24275 3438
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 16481 3226 16547 3229
rect 22093 3226 22159 3229
rect 16481 3224 22159 3226
rect 16481 3168 16486 3224
rect 16542 3168 22098 3224
rect 22154 3168 22159 3224
rect 16481 3166 22159 3168
rect 16481 3163 16547 3166
rect 22093 3163 22159 3166
rect 289 3088 7666 3090
rect 289 3032 294 3088
rect 350 3032 7666 3088
rect 289 3030 7666 3032
rect 11881 3090 11947 3093
rect 18689 3090 18755 3093
rect 24761 3090 24827 3093
rect 11881 3088 18755 3090
rect 11881 3032 11886 3088
rect 11942 3032 18694 3088
rect 18750 3032 18755 3088
rect 11881 3030 18755 3032
rect 289 3027 355 3030
rect 11881 3027 11947 3030
rect 18689 3027 18755 3030
rect 18830 3088 24827 3090
rect 18830 3032 24766 3088
rect 24822 3032 24827 3088
rect 18830 3030 24827 3032
rect 9029 2954 9095 2957
rect 18830 2954 18890 3030
rect 24761 3027 24827 3030
rect 9029 2952 18890 2954
rect 9029 2896 9034 2952
rect 9090 2896 18890 2952
rect 9029 2894 18890 2896
rect 23657 2954 23723 2957
rect 27520 2954 28000 2984
rect 23657 2952 28000 2954
rect 23657 2896 23662 2952
rect 23718 2896 28000 2952
rect 23657 2894 28000 2896
rect 9029 2891 9095 2894
rect 23657 2891 23723 2894
rect 27520 2864 28000 2894
rect 13169 2818 13235 2821
rect 17585 2818 17651 2821
rect 13169 2816 17651 2818
rect 13169 2760 13174 2816
rect 13230 2760 17590 2816
rect 17646 2760 17651 2816
rect 13169 2758 17651 2760
rect 13169 2755 13235 2758
rect 17585 2755 17651 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 20621 2682 20687 2685
rect 22553 2682 22619 2685
rect 23933 2682 23999 2685
rect 20621 2680 22619 2682
rect 20621 2624 20626 2680
rect 20682 2624 22558 2680
rect 22614 2624 22619 2680
rect 20621 2622 22619 2624
rect 20621 2619 20687 2622
rect 22553 2619 22619 2622
rect 23430 2680 23999 2682
rect 23430 2624 23938 2680
rect 23994 2624 23999 2680
rect 23430 2622 23999 2624
rect 11053 2546 11119 2549
rect 14457 2546 14523 2549
rect 11053 2544 14523 2546
rect 11053 2488 11058 2544
rect 11114 2488 14462 2544
rect 14518 2488 14523 2544
rect 11053 2486 14523 2488
rect 11053 2483 11119 2486
rect 14457 2483 14523 2486
rect 14733 2546 14799 2549
rect 19609 2546 19675 2549
rect 14733 2544 19675 2546
rect 14733 2488 14738 2544
rect 14794 2488 19614 2544
rect 19670 2488 19675 2544
rect 14733 2486 19675 2488
rect 14733 2483 14799 2486
rect 19609 2483 19675 2486
rect 20161 2546 20227 2549
rect 23430 2546 23490 2622
rect 23933 2619 23999 2622
rect 20161 2544 23490 2546
rect 20161 2488 20166 2544
rect 20222 2488 23490 2544
rect 20161 2486 23490 2488
rect 23657 2546 23723 2549
rect 24485 2546 24551 2549
rect 23657 2544 24551 2546
rect 23657 2488 23662 2544
rect 23718 2488 24490 2544
rect 24546 2488 24551 2544
rect 23657 2486 24551 2488
rect 20161 2483 20227 2486
rect 23657 2483 23723 2486
rect 24485 2483 24551 2486
rect 22001 2410 22067 2413
rect 22001 2408 24962 2410
rect 22001 2352 22006 2408
rect 22062 2352 24962 2408
rect 22001 2350 24962 2352
rect 22001 2347 22067 2350
rect 16113 2274 16179 2277
rect 18413 2274 18479 2277
rect 22645 2274 22711 2277
rect 16113 2272 22711 2274
rect 16113 2216 16118 2272
rect 16174 2216 18418 2272
rect 18474 2216 22650 2272
rect 22706 2216 22711 2272
rect 16113 2214 22711 2216
rect 24902 2274 24962 2350
rect 27520 2274 28000 2304
rect 24902 2214 28000 2274
rect 16113 2211 16179 2214
rect 18413 2211 18479 2214
rect 22645 2211 22711 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 27520 2184 28000 2214
rect 24277 2143 24597 2144
rect 9949 2138 10015 2141
rect 14733 2138 14799 2141
rect 9949 2136 14799 2138
rect 9949 2080 9954 2136
rect 10010 2080 14738 2136
rect 14794 2080 14799 2136
rect 9949 2078 14799 2080
rect 9949 2075 10015 2078
rect 14733 2075 14799 2078
rect 17033 2138 17099 2141
rect 19425 2138 19491 2141
rect 17033 2136 19491 2138
rect 17033 2080 17038 2136
rect 17094 2080 19430 2136
rect 19486 2080 19491 2136
rect 17033 2078 19491 2080
rect 17033 2075 17099 2078
rect 19425 2075 19491 2078
rect 19609 2138 19675 2141
rect 23565 2138 23631 2141
rect 19609 2136 23631 2138
rect 19609 2080 19614 2136
rect 19670 2080 23570 2136
rect 23626 2080 23631 2136
rect 19609 2078 23631 2080
rect 19609 2075 19675 2078
rect 23565 2075 23631 2078
rect 14457 2002 14523 2005
rect 22001 2002 22067 2005
rect 14457 2000 22067 2002
rect 14457 1944 14462 2000
rect 14518 1944 22006 2000
rect 22062 1944 22067 2000
rect 14457 1942 22067 1944
rect 14457 1939 14523 1942
rect 22001 1939 22067 1942
rect 8201 1866 8267 1869
rect 23197 1866 23263 1869
rect 8201 1864 23263 1866
rect 8201 1808 8206 1864
rect 8262 1808 23202 1864
rect 23258 1808 23263 1864
rect 8201 1806 23263 1808
rect 8201 1803 8267 1806
rect 23197 1803 23263 1806
rect 10501 1730 10567 1733
rect 17033 1730 17099 1733
rect 10501 1728 17099 1730
rect 10501 1672 10506 1728
rect 10562 1672 17038 1728
rect 17094 1672 17099 1728
rect 10501 1670 17099 1672
rect 10501 1667 10567 1670
rect 17033 1667 17099 1670
rect 17217 1730 17283 1733
rect 25129 1730 25195 1733
rect 17217 1728 25195 1730
rect 17217 1672 17222 1728
rect 17278 1672 25134 1728
rect 25190 1672 25195 1728
rect 17217 1670 25195 1672
rect 17217 1667 17283 1670
rect 25129 1667 25195 1670
rect 6821 1594 6887 1597
rect 23657 1594 23723 1597
rect 6821 1592 23723 1594
rect 6821 1536 6826 1592
rect 6882 1536 23662 1592
rect 23718 1536 23723 1592
rect 6821 1534 23723 1536
rect 6821 1531 6887 1534
rect 23657 1531 23723 1534
rect 24669 1594 24735 1597
rect 27520 1594 28000 1624
rect 24669 1592 28000 1594
rect 24669 1536 24674 1592
rect 24730 1536 28000 1592
rect 24669 1534 28000 1536
rect 24669 1531 24735 1534
rect 27520 1504 28000 1534
rect 4245 1458 4311 1461
rect 17217 1458 17283 1461
rect 4245 1456 17283 1458
rect 4245 1400 4250 1456
rect 4306 1400 17222 1456
rect 17278 1400 17283 1456
rect 4245 1398 17283 1400
rect 4245 1395 4311 1398
rect 17217 1395 17283 1398
rect 18597 1458 18663 1461
rect 22737 1458 22803 1461
rect 18597 1456 22803 1458
rect 18597 1400 18602 1456
rect 18658 1400 22742 1456
rect 22798 1400 22803 1456
rect 18597 1398 22803 1400
rect 18597 1395 18663 1398
rect 22737 1395 22803 1398
rect 12801 1050 12867 1053
rect 12801 1048 27538 1050
rect 12801 992 12806 1048
rect 12862 992 27538 1048
rect 12801 990 27538 992
rect 12801 987 12867 990
rect 27478 944 27538 990
rect 27478 854 28000 944
rect 27520 824 28000 854
rect 25681 370 25747 373
rect 27520 370 28000 400
rect 25681 368 28000 370
rect 25681 312 25686 368
rect 25742 312 28000 368
rect 25681 310 28000 312
rect 25681 307 25747 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 24716 19408 24780 19412
rect 24716 19352 24766 19408
rect 24766 19352 24780 19408
rect 24716 19348 24780 19352
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 24716 3708 24780 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24715 19412 24781 19413
rect 24715 19348 24716 19412
rect 24780 19348 24781 19412
rect 24715 19347 24781 19348
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24718 3773 24778 19347
rect 24715 3772 24781 3773
rect 24715 3708 24716 3772
rect 24780 3708 24781 3772
rect 24715 3707 24781 3708
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _50_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__50__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_36 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_40 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_46 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_51
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_55
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_61
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_78
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_91
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_110
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_104
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_122
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_153
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_163
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_172
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _12_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_190
timestamp 1586364061
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_192
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_213
timestamp 1586364061
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_241
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_264
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_0_272
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_268
timestamp 1586364061
transform 1 0 25760 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_276
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_189
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_234
timestamp 1586364061
transform 1 0 22632 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_238
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_262
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 590 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_141
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_150
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18124 0 1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 314 592
use scs8hd_buf_4  mux_right_track_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_268
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_272
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 590 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_66
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_172
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 774 592
use scs8hd_conb_1  _14_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 22724 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_233
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_237
timestamp 1586364061
transform 1 0 22908 0 -1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 1786 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_260
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_272
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_165
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_189
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _15_
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _24_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _10_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 1786 592
use scs8hd_conb_1  _08_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_218
timestamp 1586364061
transform 1 0 21160 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_218
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_226
timestamp 1586364061
transform 1 0 21896 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_238
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_251
timestamp 1586364061
transform 1 0 24196 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_248
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_252
timestamp 1586364061
transform 1 0 24288 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24656 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_8  FILLER_7_267
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_262
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_172
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_conb_1  _13_
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_242
timestamp 1586364061
transform 1 0 23368 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_183
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_219
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_231
timestamp 1586364061
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_255
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_43
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_190
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_242
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_21
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_196
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_238
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_250
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_262
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_conb_1  _11_
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_200
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _09_
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_223
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_234
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_246
timestamp 1586364061
transform 1 0 23736 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_258
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_270
timestamp 1586364061
transform 1 0 25944 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_253
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _26_
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _27_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _28_
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _29_
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_253
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_263
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _30_
timestamp 1586364061
transform 1 0 23828 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_242
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_251
timestamp 1586364061
transform 1 0 24196 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_255
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_267
timestamp 1586364061
transform 1 0 25668 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_2  _31_
timestamp 1586364061
transform 1 0 23184 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_244
timestamp 1586364061
transform 1 0 23552 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_256
timestamp 1586364061
transform 1 0 24656 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_268
timestamp 1586364061
transform 1 0 25760 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_237
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_6  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 21620 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_241
timestamp 1586364061
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_231
timestamp 1586364061
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_243
timestamp 1586364061
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_255
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_200
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_207
timestamp 1586364061
transform 1 0 20148 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_216
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_228
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_198
timestamp 1586364061
transform 1 0 19320 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_192
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_201
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_213
timestamp 1586364061
transform 1 0 20700 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_237
timestamp 1586364061
transform 1 0 22908 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_243
timestamp 1586364061
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_259
timestamp 1586364061
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_182
timestamp 1586364061
transform 1 0 17848 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_194
timestamp 1586364061
transform 1 0 18952 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_165
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 774 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_162
timestamp 1586364061
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_179
timestamp 1586364061
transform 1 0 17572 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_203
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_153
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_157
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_169
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_181
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _25_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 14016 480 14136 6 ccff_head
port 1 nsew default input
rlabel metal2 s 14002 27520 14058 28000 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27520 21496 28000 21616 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27520 22856 28000 22976 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27520 23536 28000 23656 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27520 24896 28000 25016 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27520 25576 28000 25696 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27520 26256 28000 26376 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27520 15512 28000 15632 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27520 16872 28000 16992 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27520 17552 28000 17672 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27520 18232 28000 18352 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27520 280 28000 400 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27520 10208 28000 10328 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27520 10888 28000 11008 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27520 11568 28000 11688 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27520 12928 28000 13048 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27520 824 28000 944 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 1504 28000 1624 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 2184 28000 2304 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27520 2864 28000 2984 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 3544 28000 3664 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 4224 28000 4344 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 5584 28000 5704 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26882 0 26938 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 prog_clk
port 83 nsew default input
rlabel metal3 s 27520 26936 28000 27056 6 right_top_grid_pin_1_
port 84 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 85 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 86 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
