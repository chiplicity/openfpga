VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__2_
  CLASS BLOCK ;
  FOREIGN sb_0__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 2.400 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 137.600 52.810 140.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 2.400 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.450 137.600 122.730 140.000 ;
    END
  END SC_OUT_TOP
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 137.600 87.770 140.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.840 140.000 24.440 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 52.400 140.000 53.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 55.120 140.000 55.720 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 58.520 140.000 59.120 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 61.240 140.000 61.840 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 63.960 140.000 64.560 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.680 140.000 67.280 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 72.800 140.000 73.400 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 75.520 140.000 76.120 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 78.240 140.000 78.840 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 26.560 140.000 27.160 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.960 140.000 30.560 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 32.680 140.000 33.280 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 35.400 140.000 36.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 40.840 140.000 41.440 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 46.960 140.000 47.560 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.680 140.000 50.280 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.960 140.000 81.560 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 109.520 140.000 110.120 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.640 140.000 116.240 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 118.360 140.000 118.960 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.080 140.000 121.680 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 123.800 140.000 124.400 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.920 140.000 130.520 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 132.640 140.000 133.240 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 135.360 140.000 135.960 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 83.680 140.000 84.280 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.080 140.000 87.680 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.800 140.000 90.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 92.520 140.000 93.120 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.240 140.000 95.840 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 97.960 140.000 98.560 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.080 140.000 104.680 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 106.800 140.000 107.400 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 2.400 ;
    END
  END chany_bottom_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 137.600 17.850 140.000 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 1.400 140.000 2.000 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.120 140.000 4.720 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 9.560 140.000 10.160 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 12.280 140.000 12.880 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.680 140.000 16.280 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 21.120 140.000 21.720 ;
    END
  END right_bottom_grid_pin_41_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 138.080 140.000 138.680 ;
    END
  END right_top_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 5.520 2.760 134.710 128.080 ;
      LAYER met2 ;
        RECT 1.470 137.320 17.290 138.565 ;
        RECT 18.130 137.320 52.250 138.565 ;
        RECT 53.090 137.320 87.210 138.565 ;
        RECT 88.050 137.320 122.170 138.565 ;
        RECT 123.010 137.320 137.910 138.565 ;
        RECT 1.470 2.680 137.910 137.320 ;
        RECT 2.030 1.515 4.410 2.680 ;
        RECT 5.250 1.515 7.630 2.680 ;
        RECT 8.470 1.515 10.850 2.680 ;
        RECT 11.690 1.515 14.070 2.680 ;
        RECT 14.910 1.515 17.290 2.680 ;
        RECT 18.130 1.515 20.510 2.680 ;
        RECT 21.350 1.515 23.730 2.680 ;
        RECT 24.570 1.515 26.950 2.680 ;
        RECT 27.790 1.515 30.170 2.680 ;
        RECT 31.010 1.515 33.390 2.680 ;
        RECT 34.230 1.515 36.610 2.680 ;
        RECT 37.450 1.515 39.830 2.680 ;
        RECT 40.670 1.515 43.050 2.680 ;
        RECT 43.890 1.515 46.270 2.680 ;
        RECT 47.110 1.515 49.950 2.680 ;
        RECT 50.790 1.515 53.170 2.680 ;
        RECT 54.010 1.515 56.390 2.680 ;
        RECT 57.230 1.515 59.610 2.680 ;
        RECT 60.450 1.515 62.830 2.680 ;
        RECT 63.670 1.515 66.050 2.680 ;
        RECT 66.890 1.515 69.270 2.680 ;
        RECT 70.110 1.515 72.490 2.680 ;
        RECT 73.330 1.515 75.710 2.680 ;
        RECT 76.550 1.515 78.930 2.680 ;
        RECT 79.770 1.515 82.150 2.680 ;
        RECT 82.990 1.515 85.370 2.680 ;
        RECT 86.210 1.515 88.590 2.680 ;
        RECT 89.430 1.515 91.810 2.680 ;
        RECT 92.650 1.515 95.490 2.680 ;
        RECT 96.330 1.515 98.710 2.680 ;
        RECT 99.550 1.515 101.930 2.680 ;
        RECT 102.770 1.515 105.150 2.680 ;
        RECT 105.990 1.515 108.370 2.680 ;
        RECT 109.210 1.515 111.590 2.680 ;
        RECT 112.430 1.515 114.810 2.680 ;
        RECT 115.650 1.515 118.030 2.680 ;
        RECT 118.870 1.515 121.250 2.680 ;
        RECT 122.090 1.515 124.470 2.680 ;
        RECT 125.310 1.515 127.690 2.680 ;
        RECT 128.530 1.515 130.910 2.680 ;
        RECT 131.750 1.515 134.130 2.680 ;
        RECT 134.970 1.515 137.350 2.680 ;
      LAYER met3 ;
        RECT 1.445 137.680 137.200 138.545 ;
        RECT 1.445 136.360 137.935 137.680 ;
        RECT 1.445 134.960 137.200 136.360 ;
        RECT 1.445 133.640 137.935 134.960 ;
        RECT 1.445 132.240 137.200 133.640 ;
        RECT 1.445 130.920 137.935 132.240 ;
        RECT 1.445 129.520 137.200 130.920 ;
        RECT 1.445 127.520 137.935 129.520 ;
        RECT 1.445 126.120 137.200 127.520 ;
        RECT 1.445 124.800 137.935 126.120 ;
        RECT 1.445 123.400 137.200 124.800 ;
        RECT 1.445 122.080 137.935 123.400 ;
        RECT 1.445 120.680 137.200 122.080 ;
        RECT 1.445 119.360 137.935 120.680 ;
        RECT 1.445 117.960 137.200 119.360 ;
        RECT 1.445 116.640 137.935 117.960 ;
        RECT 1.445 115.240 137.200 116.640 ;
        RECT 1.445 113.240 137.935 115.240 ;
        RECT 1.445 111.840 137.200 113.240 ;
        RECT 1.445 110.520 137.935 111.840 ;
        RECT 1.445 109.120 137.200 110.520 ;
        RECT 1.445 107.800 137.935 109.120 ;
        RECT 1.445 106.400 137.200 107.800 ;
        RECT 1.445 105.080 137.935 106.400 ;
        RECT 1.445 103.680 137.200 105.080 ;
        RECT 1.445 102.360 137.935 103.680 ;
        RECT 1.445 100.960 137.200 102.360 ;
        RECT 1.445 98.960 137.935 100.960 ;
        RECT 1.445 97.560 137.200 98.960 ;
        RECT 1.445 96.240 137.935 97.560 ;
        RECT 1.445 94.840 137.200 96.240 ;
        RECT 1.445 93.520 137.935 94.840 ;
        RECT 1.445 92.120 137.200 93.520 ;
        RECT 1.445 90.800 137.935 92.120 ;
        RECT 1.445 89.400 137.200 90.800 ;
        RECT 1.445 88.080 137.935 89.400 ;
        RECT 1.445 86.680 137.200 88.080 ;
        RECT 1.445 84.680 137.935 86.680 ;
        RECT 1.445 83.280 137.200 84.680 ;
        RECT 1.445 81.960 137.935 83.280 ;
        RECT 1.445 80.560 137.200 81.960 ;
        RECT 1.445 79.240 137.935 80.560 ;
        RECT 1.445 77.840 137.200 79.240 ;
        RECT 1.445 76.520 137.935 77.840 ;
        RECT 1.445 75.120 137.200 76.520 ;
        RECT 1.445 73.800 137.935 75.120 ;
        RECT 1.445 72.400 137.200 73.800 ;
        RECT 1.445 71.080 137.935 72.400 ;
        RECT 2.800 70.400 137.935 71.080 ;
        RECT 2.800 69.680 137.200 70.400 ;
        RECT 1.445 69.000 137.200 69.680 ;
        RECT 1.445 67.680 137.935 69.000 ;
        RECT 1.445 66.280 137.200 67.680 ;
        RECT 1.445 64.960 137.935 66.280 ;
        RECT 1.445 63.560 137.200 64.960 ;
        RECT 1.445 62.240 137.935 63.560 ;
        RECT 1.445 60.840 137.200 62.240 ;
        RECT 1.445 59.520 137.935 60.840 ;
        RECT 1.445 58.120 137.200 59.520 ;
        RECT 1.445 56.120 137.935 58.120 ;
        RECT 1.445 54.720 137.200 56.120 ;
        RECT 1.445 53.400 137.935 54.720 ;
        RECT 1.445 52.000 137.200 53.400 ;
        RECT 1.445 50.680 137.935 52.000 ;
        RECT 1.445 49.280 137.200 50.680 ;
        RECT 1.445 47.960 137.935 49.280 ;
        RECT 1.445 46.560 137.200 47.960 ;
        RECT 1.445 45.240 137.935 46.560 ;
        RECT 1.445 43.840 137.200 45.240 ;
        RECT 1.445 41.840 137.935 43.840 ;
        RECT 1.445 40.440 137.200 41.840 ;
        RECT 1.445 39.120 137.935 40.440 ;
        RECT 1.445 37.720 137.200 39.120 ;
        RECT 1.445 36.400 137.935 37.720 ;
        RECT 1.445 35.000 137.200 36.400 ;
        RECT 1.445 33.680 137.935 35.000 ;
        RECT 1.445 32.280 137.200 33.680 ;
        RECT 1.445 30.960 137.935 32.280 ;
        RECT 1.445 29.560 137.200 30.960 ;
        RECT 1.445 27.560 137.935 29.560 ;
        RECT 1.445 26.160 137.200 27.560 ;
        RECT 1.445 24.840 137.935 26.160 ;
        RECT 1.445 23.440 137.200 24.840 ;
        RECT 1.445 22.120 137.935 23.440 ;
        RECT 1.445 20.720 137.200 22.120 ;
        RECT 1.445 19.400 137.935 20.720 ;
        RECT 1.445 18.000 137.200 19.400 ;
        RECT 1.445 16.680 137.935 18.000 ;
        RECT 1.445 15.280 137.200 16.680 ;
        RECT 1.445 13.280 137.935 15.280 ;
        RECT 1.445 11.880 137.200 13.280 ;
        RECT 1.445 10.560 137.935 11.880 ;
        RECT 1.445 9.160 137.200 10.560 ;
        RECT 1.445 7.840 137.935 9.160 ;
        RECT 1.445 6.440 137.200 7.840 ;
        RECT 1.445 5.120 137.935 6.440 ;
        RECT 1.445 3.720 137.200 5.120 ;
        RECT 1.445 2.400 137.935 3.720 ;
        RECT 1.445 1.535 137.200 2.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_0__2_
END LIBRARY

