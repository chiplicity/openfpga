VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2223.700 BY 2027.600 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1314.570 1981.720 1314.850 1984.120 ;
    END
  END address[0]
  PIN address[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1589.120 51.880 1589.720 ;
    END
  END address[10]
  PIN address[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1780.090 44.120 1780.370 46.520 ;
    END
  END address[11]
  PIN address[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1650.320 51.880 1650.920 ;
    END
  END address[12]
  PIN address[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1710.840 51.880 1711.440 ;
    END
  END address[13]
  PIN address[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1816.240 2174.480 1816.840 ;
    END
  END address[14]
  PIN address[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1771.360 51.880 1771.960 ;
    END
  END address[15]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1682.960 2174.480 1683.560 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1537.210 44.120 1537.490 46.520 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.770 1981.720 1416.050 1984.120 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1528.600 51.880 1529.200 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1597.930 44.120 1598.210 46.520 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1658.650 44.120 1658.930 46.520 ;
    END
  END address[6]
  PIN address[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1749.600 2174.480 1750.200 ;
    END
  END address[7]
  PIN address[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1719.370 44.120 1719.650 46.520 ;
    END
  END address[8]
  PIN address[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1516.970 1981.720 1517.250 1984.120 ;
    END
  END address[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1840.810 44.120 1841.090 46.520 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1618.170 1981.720 1618.450 1984.120 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1901.530 44.120 1901.810 46.520 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 100.170 1981.720 100.450 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 504.970 1981.720 505.250 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[10]
  PIN gfpga_pad_GPIO_PAD[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 606.170 1981.720 606.450 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[11]
  PIN gfpga_pad_GPIO_PAD[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 707.370 1981.720 707.650 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[12]
  PIN gfpga_pad_GPIO_PAD[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 808.570 1981.720 808.850 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[13]
  PIN gfpga_pad_GPIO_PAD[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1831.880 51.880 1832.480 ;
    END
  END gfpga_pad_GPIO_PAD[14]
  PIN gfpga_pad_GPIO_PAD[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2144.410 44.120 2144.690 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[15]
  PIN gfpga_pad_GPIO_PAD[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1921.770 1981.720 1922.050 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[16]
  PIN gfpga_pad_GPIO_PAD[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2022.970 1981.720 2023.250 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[17]
  PIN gfpga_pad_GPIO_PAD[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2124.170 1981.720 2124.450 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[18]
  PIN gfpga_pad_GPIO_PAD[19]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1892.400 51.880 1893.000 ;
    END
  END gfpga_pad_GPIO_PAD[19]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 201.370 1981.720 201.650 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 909.770 1981.720 910.050 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[20]
  PIN gfpga_pad_GPIO_PAD[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1010.970 1981.720 1011.250 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[21]
  PIN gfpga_pad_GPIO_PAD[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1112.170 1981.720 1112.450 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[22]
  PIN gfpga_pad_GPIO_PAD[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1213.370 1981.720 1213.650 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[23]
  PIN gfpga_pad_GPIO_PAD[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 77.480 2174.480 78.080 ;
    END
  END gfpga_pad_GPIO_PAD[24]
  PIN gfpga_pad_GPIO_PAD[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 144.120 2174.480 144.720 ;
    END
  END gfpga_pad_GPIO_PAD[25]
  PIN gfpga_pad_GPIO_PAD[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 210.760 2174.480 211.360 ;
    END
  END gfpga_pad_GPIO_PAD[26]
  PIN gfpga_pad_GPIO_PAD[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 278.080 2174.480 278.680 ;
    END
  END gfpga_pad_GPIO_PAD[27]
  PIN gfpga_pad_GPIO_PAD[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 344.720 2174.480 345.320 ;
    END
  END gfpga_pad_GPIO_PAD[28]
  PIN gfpga_pad_GPIO_PAD[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 411.360 2174.480 411.960 ;
    END
  END gfpga_pad_GPIO_PAD[29]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 302.570 1981.720 302.850 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 478.680 2174.480 479.280 ;
    END
  END gfpga_pad_GPIO_PAD[30]
  PIN gfpga_pad_GPIO_PAD[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 545.320 2174.480 545.920 ;
    END
  END gfpga_pad_GPIO_PAD[31]
  PIN gfpga_pad_GPIO_PAD[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 612.640 2174.480 613.240 ;
    END
  END gfpga_pad_GPIO_PAD[32]
  PIN gfpga_pad_GPIO_PAD[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 679.280 2174.480 679.880 ;
    END
  END gfpga_pad_GPIO_PAD[33]
  PIN gfpga_pad_GPIO_PAD[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 745.920 2174.480 746.520 ;
    END
  END gfpga_pad_GPIO_PAD[34]
  PIN gfpga_pad_GPIO_PAD[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 813.240 2174.480 813.840 ;
    END
  END gfpga_pad_GPIO_PAD[35]
  PIN gfpga_pad_GPIO_PAD[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 879.880 2174.480 880.480 ;
    END
  END gfpga_pad_GPIO_PAD[36]
  PIN gfpga_pad_GPIO_PAD[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 946.520 2174.480 947.120 ;
    END
  END gfpga_pad_GPIO_PAD[37]
  PIN gfpga_pad_GPIO_PAD[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1013.840 2174.480 1014.440 ;
    END
  END gfpga_pad_GPIO_PAD[38]
  PIN gfpga_pad_GPIO_PAD[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1080.480 2174.480 1081.080 ;
    END
  END gfpga_pad_GPIO_PAD[39]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 403.770 1981.720 404.050 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1147.800 2174.480 1148.400 ;
    END
  END gfpga_pad_GPIO_PAD[40]
  PIN gfpga_pad_GPIO_PAD[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1214.440 2174.480 1215.040 ;
    END
  END gfpga_pad_GPIO_PAD[41]
  PIN gfpga_pad_GPIO_PAD[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1281.080 2174.480 1281.680 ;
    END
  END gfpga_pad_GPIO_PAD[42]
  PIN gfpga_pad_GPIO_PAD[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1348.400 2174.480 1349.000 ;
    END
  END gfpga_pad_GPIO_PAD[43]
  PIN gfpga_pad_GPIO_PAD[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1415.040 2174.480 1415.640 ;
    END
  END gfpga_pad_GPIO_PAD[44]
  PIN gfpga_pad_GPIO_PAD[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1481.680 2174.480 1482.280 ;
    END
  END gfpga_pad_GPIO_PAD[45]
  PIN gfpga_pad_GPIO_PAD[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1549.000 2174.480 1549.600 ;
    END
  END gfpga_pad_GPIO_PAD[46]
  PIN gfpga_pad_GPIO_PAD[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1615.640 2174.480 1616.240 ;
    END
  END gfpga_pad_GPIO_PAD[47]
  PIN gfpga_pad_GPIO_PAD[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 79.930 44.120 80.210 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[48]
  PIN gfpga_pad_GPIO_PAD[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 140.650 44.120 140.930 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[49]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1719.370 1981.720 1719.650 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 201.370 44.120 201.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[50]
  PIN gfpga_pad_GPIO_PAD[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 262.090 44.120 262.370 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[51]
  PIN gfpga_pad_GPIO_PAD[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 322.810 44.120 323.090 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[52]
  PIN gfpga_pad_GPIO_PAD[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 383.530 44.120 383.810 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[53]
  PIN gfpga_pad_GPIO_PAD[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 444.250 44.120 444.530 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[54]
  PIN gfpga_pad_GPIO_PAD[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 504.970 44.120 505.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[55]
  PIN gfpga_pad_GPIO_PAD[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 565.690 44.120 565.970 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[56]
  PIN gfpga_pad_GPIO_PAD[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 626.410 44.120 626.690 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[57]
  PIN gfpga_pad_GPIO_PAD[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 687.130 44.120 687.410 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[58]
  PIN gfpga_pad_GPIO_PAD[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 747.850 44.120 748.130 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[59]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1820.570 1981.720 1820.850 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 808.570 44.120 808.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[60]
  PIN gfpga_pad_GPIO_PAD[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 869.290 44.120 869.570 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[61]
  PIN gfpga_pad_GPIO_PAD[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 930.010 44.120 930.290 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[62]
  PIN gfpga_pad_GPIO_PAD[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 990.730 44.120 991.010 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[63]
  PIN gfpga_pad_GPIO_PAD[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1051.450 44.120 1051.730 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[64]
  PIN gfpga_pad_GPIO_PAD[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1112.170 44.120 1112.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[65]
  PIN gfpga_pad_GPIO_PAD[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1172.890 44.120 1173.170 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[66]
  PIN gfpga_pad_GPIO_PAD[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1233.610 44.120 1233.890 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[67]
  PIN gfpga_pad_GPIO_PAD[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1294.330 44.120 1294.610 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[68]
  PIN gfpga_pad_GPIO_PAD[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1355.050 44.120 1355.330 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[69]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1962.250 44.120 1962.530 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1415.770 44.120 1416.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[70]
  PIN gfpga_pad_GPIO_PAD[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1476.490 44.120 1476.770 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[71]
  PIN gfpga_pad_GPIO_PAD[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 74.080 51.880 74.680 ;
    END
  END gfpga_pad_GPIO_PAD[72]
  PIN gfpga_pad_GPIO_PAD[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 134.600 51.880 135.200 ;
    END
  END gfpga_pad_GPIO_PAD[73]
  PIN gfpga_pad_GPIO_PAD[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 195.120 51.880 195.720 ;
    END
  END gfpga_pad_GPIO_PAD[74]
  PIN gfpga_pad_GPIO_PAD[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 255.640 51.880 256.240 ;
    END
  END gfpga_pad_GPIO_PAD[75]
  PIN gfpga_pad_GPIO_PAD[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 316.160 51.880 316.760 ;
    END
  END gfpga_pad_GPIO_PAD[76]
  PIN gfpga_pad_GPIO_PAD[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 376.680 51.880 377.280 ;
    END
  END gfpga_pad_GPIO_PAD[77]
  PIN gfpga_pad_GPIO_PAD[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 437.200 51.880 437.800 ;
    END
  END gfpga_pad_GPIO_PAD[78]
  PIN gfpga_pad_GPIO_PAD[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 498.400 51.880 499.000 ;
    END
  END gfpga_pad_GPIO_PAD[79]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1883.560 2174.480 1884.160 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN gfpga_pad_GPIO_PAD[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 558.920 51.880 559.520 ;
    END
  END gfpga_pad_GPIO_PAD[80]
  PIN gfpga_pad_GPIO_PAD[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 619.440 51.880 620.040 ;
    END
  END gfpga_pad_GPIO_PAD[81]
  PIN gfpga_pad_GPIO_PAD[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 679.960 51.880 680.560 ;
    END
  END gfpga_pad_GPIO_PAD[82]
  PIN gfpga_pad_GPIO_PAD[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 740.480 51.880 741.080 ;
    END
  END gfpga_pad_GPIO_PAD[83]
  PIN gfpga_pad_GPIO_PAD[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 801.000 51.880 801.600 ;
    END
  END gfpga_pad_GPIO_PAD[84]
  PIN gfpga_pad_GPIO_PAD[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 862.200 51.880 862.800 ;
    END
  END gfpga_pad_GPIO_PAD[85]
  PIN gfpga_pad_GPIO_PAD[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 922.720 51.880 923.320 ;
    END
  END gfpga_pad_GPIO_PAD[86]
  PIN gfpga_pad_GPIO_PAD[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 983.240 51.880 983.840 ;
    END
  END gfpga_pad_GPIO_PAD[87]
  PIN gfpga_pad_GPIO_PAD[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1043.760 51.880 1044.360 ;
    END
  END gfpga_pad_GPIO_PAD[88]
  PIN gfpga_pad_GPIO_PAD[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1104.280 51.880 1104.880 ;
    END
  END gfpga_pad_GPIO_PAD[89]
  PIN gfpga_pad_GPIO_PAD[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2022.970 44.120 2023.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[8]
  PIN gfpga_pad_GPIO_PAD[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1164.800 51.880 1165.400 ;
    END
  END gfpga_pad_GPIO_PAD[90]
  PIN gfpga_pad_GPIO_PAD[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1225.320 51.880 1225.920 ;
    END
  END gfpga_pad_GPIO_PAD[91]
  PIN gfpga_pad_GPIO_PAD[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1286.520 51.880 1287.120 ;
    END
  END gfpga_pad_GPIO_PAD[92]
  PIN gfpga_pad_GPIO_PAD[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1347.040 51.880 1347.640 ;
    END
  END gfpga_pad_GPIO_PAD[93]
  PIN gfpga_pad_GPIO_PAD[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1407.560 51.880 1408.160 ;
    END
  END gfpga_pad_GPIO_PAD[94]
  PIN gfpga_pad_GPIO_PAD[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1468.080 51.880 1468.680 ;
    END
  END gfpga_pad_GPIO_PAD[95]
  PIN gfpga_pad_GPIO_PAD[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2083.690 44.120 2083.970 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[9]
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1950.200 2174.480 1950.800 ;
    END
  END reset
  PIN set
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1952.920 51.880 1953.520 ;
    END
  END set
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 2198.700 45.000 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 2223.700 20.000 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 105.000 104.915 2118.540 1922.205 ;
      LAYER met1 ;
        RECT 63.350 46.880 2151.610 1969.160 ;
      LAYER met2 ;
        RECT 63.370 1981.440 99.890 1981.720 ;
        RECT 100.730 1981.440 201.090 1981.720 ;
        RECT 201.930 1981.440 302.290 1981.720 ;
        RECT 303.130 1981.440 403.490 1981.720 ;
        RECT 404.330 1981.440 504.690 1981.720 ;
        RECT 505.530 1981.440 605.890 1981.720 ;
        RECT 606.730 1981.440 707.090 1981.720 ;
        RECT 707.930 1981.440 808.290 1981.720 ;
        RECT 809.130 1981.440 909.490 1981.720 ;
        RECT 910.330 1981.440 1010.690 1981.720 ;
        RECT 1011.530 1981.440 1111.890 1981.720 ;
        RECT 1112.730 1981.440 1213.090 1981.720 ;
        RECT 1213.930 1981.440 1314.290 1981.720 ;
        RECT 1315.130 1981.440 1415.490 1981.720 ;
        RECT 1416.330 1981.440 1516.690 1981.720 ;
        RECT 1517.530 1981.440 1617.890 1981.720 ;
        RECT 1618.730 1981.440 1719.090 1981.720 ;
        RECT 1719.930 1981.440 1820.290 1981.720 ;
        RECT 1821.130 1981.440 1921.490 1981.720 ;
        RECT 1922.330 1981.440 2022.690 1981.720 ;
        RECT 2023.530 1981.440 2123.890 1981.720 ;
        RECT 2124.730 1981.440 2151.590 1981.720 ;
        RECT 63.370 46.800 2151.590 1981.440 ;
        RECT 63.370 46.520 79.650 46.800 ;
        RECT 80.490 46.520 140.370 46.800 ;
        RECT 141.210 46.520 201.090 46.800 ;
        RECT 201.930 46.520 261.810 46.800 ;
        RECT 262.650 46.520 322.530 46.800 ;
        RECT 323.370 46.520 383.250 46.800 ;
        RECT 384.090 46.520 443.970 46.800 ;
        RECT 444.810 46.520 504.690 46.800 ;
        RECT 505.530 46.520 565.410 46.800 ;
        RECT 566.250 46.520 626.130 46.800 ;
        RECT 626.970 46.520 686.850 46.800 ;
        RECT 687.690 46.520 747.570 46.800 ;
        RECT 748.410 46.520 808.290 46.800 ;
        RECT 809.130 46.520 869.010 46.800 ;
        RECT 869.850 46.520 929.730 46.800 ;
        RECT 930.570 46.520 990.450 46.800 ;
        RECT 991.290 46.520 1051.170 46.800 ;
        RECT 1052.010 46.520 1111.890 46.800 ;
        RECT 1112.730 46.520 1172.610 46.800 ;
        RECT 1173.450 46.520 1233.330 46.800 ;
        RECT 1234.170 46.520 1294.050 46.800 ;
        RECT 1294.890 46.520 1354.770 46.800 ;
        RECT 1355.610 46.520 1415.490 46.800 ;
        RECT 1416.330 46.520 1476.210 46.800 ;
        RECT 1477.050 46.520 1536.930 46.800 ;
        RECT 1537.770 46.520 1597.650 46.800 ;
        RECT 1598.490 46.520 1658.370 46.800 ;
        RECT 1659.210 46.520 1719.090 46.800 ;
        RECT 1719.930 46.520 1779.810 46.800 ;
        RECT 1780.650 46.520 1840.530 46.800 ;
        RECT 1841.370 46.520 1901.250 46.800 ;
        RECT 1902.090 46.520 1961.970 46.800 ;
        RECT 1962.810 46.520 2022.690 46.800 ;
        RECT 2023.530 46.520 2083.410 46.800 ;
        RECT 2084.250 46.520 2144.130 46.800 ;
        RECT 2144.970 46.520 2151.590 46.800 ;
      LAYER met3 ;
        RECT 51.880 1953.920 2172.080 1969.025 ;
        RECT 52.280 1952.520 2172.080 1953.920 ;
        RECT 51.880 1951.200 2172.080 1952.520 ;
        RECT 51.880 1949.800 2171.680 1951.200 ;
        RECT 51.880 1893.400 2172.080 1949.800 ;
        RECT 52.280 1892.000 2172.080 1893.400 ;
        RECT 51.880 1884.560 2172.080 1892.000 ;
        RECT 51.880 1883.160 2171.680 1884.560 ;
        RECT 51.880 1832.880 2172.080 1883.160 ;
        RECT 52.280 1831.480 2172.080 1832.880 ;
        RECT 51.880 1817.240 2172.080 1831.480 ;
        RECT 51.880 1815.840 2171.680 1817.240 ;
        RECT 51.880 1772.360 2172.080 1815.840 ;
        RECT 52.280 1770.960 2172.080 1772.360 ;
        RECT 51.880 1750.600 2172.080 1770.960 ;
        RECT 51.880 1749.200 2171.680 1750.600 ;
        RECT 51.880 1711.840 2172.080 1749.200 ;
        RECT 52.280 1710.440 2172.080 1711.840 ;
        RECT 51.880 1683.960 2172.080 1710.440 ;
        RECT 51.880 1682.560 2171.680 1683.960 ;
        RECT 51.880 1651.320 2172.080 1682.560 ;
        RECT 52.280 1649.920 2172.080 1651.320 ;
        RECT 51.880 1616.640 2172.080 1649.920 ;
        RECT 51.880 1615.240 2171.680 1616.640 ;
        RECT 51.880 1590.120 2172.080 1615.240 ;
        RECT 52.280 1588.720 2172.080 1590.120 ;
        RECT 51.880 1550.000 2172.080 1588.720 ;
        RECT 51.880 1548.600 2171.680 1550.000 ;
        RECT 51.880 1529.600 2172.080 1548.600 ;
        RECT 52.280 1528.200 2172.080 1529.600 ;
        RECT 51.880 1482.680 2172.080 1528.200 ;
        RECT 51.880 1481.280 2171.680 1482.680 ;
        RECT 51.880 1469.080 2172.080 1481.280 ;
        RECT 52.280 1467.680 2172.080 1469.080 ;
        RECT 51.880 1416.040 2172.080 1467.680 ;
        RECT 51.880 1414.640 2171.680 1416.040 ;
        RECT 51.880 1408.560 2172.080 1414.640 ;
        RECT 52.280 1407.160 2172.080 1408.560 ;
        RECT 51.880 1349.400 2172.080 1407.160 ;
        RECT 51.880 1348.040 2171.680 1349.400 ;
        RECT 52.280 1348.000 2171.680 1348.040 ;
        RECT 52.280 1346.640 2172.080 1348.000 ;
        RECT 51.880 1287.520 2172.080 1346.640 ;
        RECT 52.280 1286.120 2172.080 1287.520 ;
        RECT 51.880 1282.080 2172.080 1286.120 ;
        RECT 51.880 1280.680 2171.680 1282.080 ;
        RECT 51.880 1226.320 2172.080 1280.680 ;
        RECT 52.280 1224.920 2172.080 1226.320 ;
        RECT 51.880 1215.440 2172.080 1224.920 ;
        RECT 51.880 1214.040 2171.680 1215.440 ;
        RECT 51.880 1165.800 2172.080 1214.040 ;
        RECT 52.280 1164.400 2172.080 1165.800 ;
        RECT 51.880 1148.800 2172.080 1164.400 ;
        RECT 51.880 1147.400 2171.680 1148.800 ;
        RECT 51.880 1105.280 2172.080 1147.400 ;
        RECT 52.280 1103.880 2172.080 1105.280 ;
        RECT 51.880 1081.480 2172.080 1103.880 ;
        RECT 51.880 1080.080 2171.680 1081.480 ;
        RECT 51.880 1044.760 2172.080 1080.080 ;
        RECT 52.280 1043.360 2172.080 1044.760 ;
        RECT 51.880 1014.840 2172.080 1043.360 ;
        RECT 51.880 1013.440 2171.680 1014.840 ;
        RECT 51.880 984.240 2172.080 1013.440 ;
        RECT 52.280 982.840 2172.080 984.240 ;
        RECT 51.880 947.520 2172.080 982.840 ;
        RECT 51.880 946.120 2171.680 947.520 ;
        RECT 51.880 923.720 2172.080 946.120 ;
        RECT 52.280 922.320 2172.080 923.720 ;
        RECT 51.880 880.880 2172.080 922.320 ;
        RECT 51.880 879.480 2171.680 880.880 ;
        RECT 51.880 863.200 2172.080 879.480 ;
        RECT 52.280 861.800 2172.080 863.200 ;
        RECT 51.880 814.240 2172.080 861.800 ;
        RECT 51.880 812.840 2171.680 814.240 ;
        RECT 51.880 802.000 2172.080 812.840 ;
        RECT 52.280 800.600 2172.080 802.000 ;
        RECT 51.880 746.920 2172.080 800.600 ;
        RECT 51.880 745.520 2171.680 746.920 ;
        RECT 51.880 741.480 2172.080 745.520 ;
        RECT 52.280 740.080 2172.080 741.480 ;
        RECT 51.880 680.960 2172.080 740.080 ;
        RECT 52.280 680.280 2172.080 680.960 ;
        RECT 52.280 679.560 2171.680 680.280 ;
        RECT 51.880 678.880 2171.680 679.560 ;
        RECT 51.880 620.440 2172.080 678.880 ;
        RECT 52.280 619.040 2172.080 620.440 ;
        RECT 51.880 613.640 2172.080 619.040 ;
        RECT 51.880 612.240 2171.680 613.640 ;
        RECT 51.880 559.920 2172.080 612.240 ;
        RECT 52.280 558.520 2172.080 559.920 ;
        RECT 51.880 546.320 2172.080 558.520 ;
        RECT 51.880 544.920 2171.680 546.320 ;
        RECT 51.880 499.400 2172.080 544.920 ;
        RECT 52.280 498.000 2172.080 499.400 ;
        RECT 51.880 479.680 2172.080 498.000 ;
        RECT 51.880 478.280 2171.680 479.680 ;
        RECT 51.880 438.200 2172.080 478.280 ;
        RECT 52.280 436.800 2172.080 438.200 ;
        RECT 51.880 412.360 2172.080 436.800 ;
        RECT 51.880 410.960 2171.680 412.360 ;
        RECT 51.880 377.680 2172.080 410.960 ;
        RECT 52.280 376.280 2172.080 377.680 ;
        RECT 51.880 345.720 2172.080 376.280 ;
        RECT 51.880 344.320 2171.680 345.720 ;
        RECT 51.880 317.160 2172.080 344.320 ;
        RECT 52.280 315.760 2172.080 317.160 ;
        RECT 51.880 279.080 2172.080 315.760 ;
        RECT 51.880 277.680 2171.680 279.080 ;
        RECT 51.880 256.640 2172.080 277.680 ;
        RECT 52.280 255.240 2172.080 256.640 ;
        RECT 51.880 211.760 2172.080 255.240 ;
        RECT 51.880 210.360 2171.680 211.760 ;
        RECT 51.880 196.120 2172.080 210.360 ;
        RECT 52.280 194.720 2172.080 196.120 ;
        RECT 51.880 145.120 2172.080 194.720 ;
        RECT 51.880 143.720 2171.680 145.120 ;
        RECT 51.880 135.600 2172.080 143.720 ;
        RECT 52.280 134.200 2172.080 135.600 ;
        RECT 51.880 78.480 2172.080 134.200 ;
        RECT 51.880 77.080 2171.680 78.480 ;
        RECT 51.880 75.080 2172.080 77.080 ;
        RECT 52.280 73.680 2172.080 75.080 ;
        RECT 51.880 61.295 2172.080 73.680 ;
      LAYER met4 ;
        RECT 0.000 0.000 2223.700 2027.600 ;
      LAYER met5 ;
        RECT 0.000 70.850 2223.700 2027.600 ;
  END
END fpga_top
END LIBRARY

