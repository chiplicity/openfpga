* NGSPICE file created from sb_2__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt sb_2__2_ SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_left_grid_pin_42_
+ bottom_left_grid_pin_43_ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_
+ bottom_left_grid_pin_47_ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ left_top_grid_pin_1_ prog_clk VPWR VGND
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_15.mux_l2_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_48_ bottom_left_grid_pin_46_
+ mux_bottom_track_3.mux_l1_in_0_/S mux_bottom_track_3.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_062_ _062_/HI _062_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_17.mux_l1_in_0_ chanx_left_in[9] bottom_left_grid_pin_45_ mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_29.mux_l2_in_0_ _067_/HI mux_bottom_track_29.mux_l1_in_0_/X mux_bottom_track_29.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_5 chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _111_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_3.mux_l1_in_0_ bottom_left_grid_pin_44_ bottom_left_grid_pin_42_
+ mux_bottom_track_3.mux_l1_in_0_/S mux_bottom_track_3.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_061_ _061_/HI _061_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l2_in_0_/X _088_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X _077_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_35.mux_l1_in_0_/S mux_left_track_35.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_6 chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X _080_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_3.mux_l2_in_1_/S
+ mux_bottom_track_3.mux_l3_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_29.mux_l1_in_0_ chanx_left_in[15] bottom_left_grid_pin_43_ mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ mux_left_track_7.mux_l3_in_0_/S mux_left_track_7.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_060_ _060_/HI _060_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_7.mux_l2_in_1_ _055_/HI left_bottom_grid_pin_40_ mux_left_track_7.mux_l2_in_1_/S
+ mux_left_track_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_112_ _112_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_33.mux_l2_in_0_/S mux_left_track_35.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_3.mux_l1_in_0_/S
+ mux_bottom_track_3.mux_l2_in_1_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_15.mux_l2_in_0_ _040_/HI mux_left_track_15.mux_l1_in_0_/X mux_left_track_15.mux_l2_in_0_/S
+ mux_left_track_15.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_1_/S mux_left_track_7.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_111_ _111_/A chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_8 chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_7.mux_l1_in_1_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_7.mux_l1_in_0_/S
+ mux_left_track_7.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_1.mux_l3_in_0_/S
+ mux_bottom_track_3.mux_l1_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_15.mux_l1_in_0_ left_bottom_grid_pin_36_ chany_bottom_in[6] mux_left_track_15.mux_l1_in_0_/S
+ mux_left_track_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_27.mux_l2_in_0_ _046_/HI mux_left_track_27.mux_l1_in_0_/X mux_left_track_27.mux_l2_in_0_/S
+ mux_left_track_27.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_110_ _110_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_9 chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_7.mux_l1_in_0_ left_bottom_grid_pin_34_ chany_bottom_in[2] mux_left_track_7.mux_l1_in_0_/S
+ mux_left_track_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_11.mux_l2_in_0_/X
+ _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_21.mux_l1_in_0_/S mux_left_track_21.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_7.mux_l3_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_27.mux_l1_in_0_ left_bottom_grid_pin_34_ chany_bottom_in[12] mux_left_track_27.mux_l1_in_0_/S
+ mux_left_track_27.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_39.mux_l2_in_0_ _053_/HI mux_left_track_39.mux_l1_in_0_/X ccff_tail
+ mux_left_track_39.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_13.mux_l2_in_0_ _059_/HI mux_bottom_track_13.mux_l1_in_0_/X mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_13.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_19.mux_l2_in_0_/S mux_left_track_21.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X
+ _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_099_ _099_/A chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_27.mux_l1_in_0_/S mux_left_track_27.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_39.mux_l1_in_0_ left_bottom_grid_pin_40_ chany_bottom_in[18] mux_left_track_39.mux_l1_in_0_/S
+ mux_left_track_39.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_13.mux_l1_in_0_ chanx_left_in[7] bottom_left_grid_pin_43_ mux_bottom_track_13.mux_l1_in_0_/S
+ mux_bottom_track_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_0_/S mux_bottom_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_098_ _098_/A chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_25.mux_l2_in_0_/S mux_left_track_27.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.mux_l2_in_0_ _036_/HI mux_bottom_track_9.mux_l1_in_0_/X mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l1_in_1_ _065_/HI chanx_left_in[13] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X _090_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X _082_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_097_ chanx_left_in[16] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l2_in_0_/X _085_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l1_in_0_ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_
+ mux_bottom_track_25.mux_l1_in_0_/S mux_bottom_track_25.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l1_in_0_ chanx_left_in[5] bottom_right_grid_pin_1_ mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l2_in_0_/X _108_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_1.mux_l1_in_1_/S mux_left_track_1.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.mux_l2_in_1_ _048_/HI left_bottom_grid_pin_40_ mux_left_track_3.mux_l2_in_0_/S
+ mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_096_ chanx_left_in[17] chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_7.mux_l2_in_1_/S mux_left_track_7.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_079_ _079_/A chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_0_ _038_/HI mux_left_track_11.mux_l1_in_0_/X mux_left_track_11.mux_l2_in_0_/S
+ mux_left_track_11.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_13.mux_l1_in_0_/S mux_left_track_13.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_29.mux_l2_in_0_/S mux_left_track_1.mux_l1_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.mux_l1_in_1_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_095_ chanx_left_in[18] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_7.mux_l1_in_0_/S mux_left_track_7.mux_l2_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_078_ _078_/A chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_11.mux_l1_in_0_ left_bottom_grid_pin_34_ chany_bottom_in[4] mux_left_track_11.mux_l1_in_0_/S
+ mux_left_track_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_11.mux_l2_in_0_/S mux_left_track_13.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_23.mux_l2_in_0_ _044_/HI mux_left_track_23.mux_l1_in_0_/X mux_left_track_23.mux_l2_in_0_/S
+ mux_left_track_23.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_0_ left_bottom_grid_pin_34_ chany_bottom_in[0] mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_19.mux_l1_in_0_/S mux_left_track_19.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_094_ chanx_left_in[19] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_5.mux_l3_in_0_/S mux_left_track_7.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_17.mux_l2_in_0_/S mux_left_track_19.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_23.mux_l1_in_0_ left_bottom_grid_pin_40_ chany_bottom_in[10] mux_left_track_23.mux_l1_in_0_/S
+ mux_left_track_23.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_093_ chanx_left_in[0] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_35.mux_l2_in_0_ _051_/HI mux_left_track_35.mux_l1_in_0_/X mux_left_track_35.mux_l2_in_0_/S
+ mux_left_track_35.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_076_ _076_/A chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X
+ _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_31.mux_l1_in_0_/S mux_left_track_31.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ _059_/HI _059_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X
+ _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_5.mux_l2_in_1_ _069_/HI mux_bottom_track_5.mux_l1_in_2_/X mux_bottom_track_5.mux_l2_in_1_/S
+ mux_bottom_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_092_ _092_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_5.mux_l1_in_2_ chanx_left_in[3] bottom_left_grid_pin_49_ mux_bottom_track_5.mux_l1_in_1_/S
+ mux_bottom_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_075_ _075_/A chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_29.mux_l2_in_0_/S mux_left_track_31.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_35.mux_l1_in_0_ left_bottom_grid_pin_38_ chany_bottom_in[16] mux_left_track_35.mux_l1_in_0_/S
+ mux_left_track_35.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_058_ _058_/HI _058_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_19.mux_l2_in_0_ _062_/HI mux_bottom_track_19.mux_l1_in_0_/X mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_21.mux_l2_in_0_ _063_/HI mux_bottom_track_21.mux_l1_in_0_/X mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_37.mux_l1_in_0_/S mux_left_track_37.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X _092_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_5.mux_l2_in_1_/S
+ mux_bottom_track_5.mux_l3_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_091_ _091_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_074_ _074_/A chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_5.mux_l1_in_1_/S mux_bottom_track_5.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_057_ _057_/HI _057_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_25.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_109_ _109_/A chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_35.mux_l2_in_0_/S mux_left_track_37.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l2_in_0_/X _087_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_19.mux_l1_in_0_ chanx_left_in[10] bottom_left_grid_pin_46_ mux_bottom_track_19.mux_l1_in_0_/S
+ mux_bottom_track_19.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_21.mux_l1_in_0_ chanx_left_in[11] bottom_left_grid_pin_47_ mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_5.mux_l1_in_1_/S
+ mux_bottom_track_5.mux_l2_in_1_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_090_ _090_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _110_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_43_ bottom_right_grid_pin_1_
+ mux_bottom_track_5.mux_l1_in_1_/S mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_073_ _073_/A chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_056_ _056_/HI _056_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_108_ _108_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X _076_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_3.mux_l3_in_0_/S
+ mux_bottom_track_5.mux_l1_in_1_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_27.sky130_fd_sc_hd__buf_4_0_ mux_left_track_27.mux_l2_in_0_/X _079_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_072_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_10 chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_107_ _107_/A chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_13.mux_l1_in_0_/S
+ mux_bottom_track_13.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_23.mux_l1_in_0_/S mux_left_track_23.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_071_ _071_/HI SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l2_in_0_ _041_/HI mux_left_track_17.mux_l1_in_0_/X mux_left_track_17.mux_l2_in_0_/S
+ mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_11 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_106_ _106_/A chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l1_in_1_ _056_/HI left_bottom_grid_pin_41_ mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_13.mux_l1_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_070_ _070_/HI SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_21.mux_l2_in_0_/S mux_left_track_23.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_12 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_19.mux_l1_in_0_/S
+ mux_bottom_track_19.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_29.mux_l1_in_0_/S mux_left_track_29.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_105_ _105_/A chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.mux_l1_in_0_ left_bottom_grid_pin_37_ chany_bottom_in[7] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_29.mux_l2_in_0_ _047_/HI mux_left_track_29.mux_l1_in_0_/X mux_left_track_29.mux_l2_in_0_/S
+ mux_left_track_29.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_31.mux_l2_in_0_ _049_/HI mux_left_track_31.mux_l1_in_0_/X mux_left_track_31.mux_l2_in_0_/S
+ mux_left_track_31.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[3] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X
+ _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_13 chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l1_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_27.mux_l2_in_0_/S mux_left_track_29.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l2_in_1_ _057_/HI mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_1_/S
+ mux_bottom_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_104_ _104_/A chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l1_in_2_ chanx_left_in[1] bottom_left_grid_pin_49_ mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_29.mux_l1_in_0_ left_bottom_grid_pin_35_ chany_bottom_in[13] mux_left_track_29.mux_l1_in_0_/S
+ mux_left_track_29.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_31.mux_l1_in_0_ left_bottom_grid_pin_36_ chany_bottom_in[14] mux_left_track_31.mux_l1_in_0_/S
+ mux_left_track_31.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_15.mux_l2_in_0_ _060_/HI mux_bottom_track_15.mux_l1_in_0_/X mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_14 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_29.mux_l2_in_0_/X
+ _098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_103_ _103_/A chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_1.mux_l1_in_1_/S mux_bottom_track_1.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_3.mux_l1_in_1_/S mux_left_track_3.mux_l2_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_15.mux_l1_in_0_ chanx_left_in[8] bottom_left_grid_pin_44_ mux_bottom_track_15.mux_l1_in_0_/S
+ mux_bottom_track_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_27.mux_l2_in_0_ _066_/HI mux_bottom_track_27.mux_l1_in_0_/X mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _112_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_102_ _102_/A chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_43_ bottom_right_grid_pin_1_
+ mux_bottom_track_1.mux_l1_in_1_/S mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_15.mux_l1_in_0_/S mux_left_track_15.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_1.mux_l3_in_0_/S mux_left_track_3.mux_l1_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X _089_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_101_ _101_/A chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X _081_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_27.mux_l1_in_0_ chanx_left_in[14] bottom_left_grid_pin_42_ mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X _084_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_13.mux_l2_in_0_/S mux_left_track_15.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_1_ _054_/HI mux_left_track_5.mux_l1_in_2_/X mux_left_track_5.mux_l2_in_1_/S
+ mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_7.mux_l3_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ _100_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_41_ left_bottom_grid_pin_39_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_13.mux_l2_in_0_ _039_/HI mux_left_track_13.mux_l1_in_0_/X mux_left_track_13.mux_l2_in_0_/S
+ mux_left_track_13.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X _073_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l1_in_1_ left_bottom_grid_pin_37_ left_bottom_grid_pin_35_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_1.mux_l2_in_1_/S
+ mux_bottom_track_1.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_13.mux_l1_in_0_ left_bottom_grid_pin_35_ chany_bottom_in[5] mux_left_track_13.mux_l1_in_0_/S
+ mux_left_track_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[1] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_25.mux_l1_in_1_ _045_/HI left_bottom_grid_pin_41_ mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_089_ _089_/A chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_31.mux_l2_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l2_in_1_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_39.mux_l1_in_0_/S ccff_tail
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_7.mux_l2_in_0_/S
+ mux_bottom_track_7.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[11] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_088_ _088_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_37.mux_l2_in_0_ _052_/HI mux_left_track_37.mux_l1_in_0_/X mux_left_track_37.mux_l2_in_0_/S
+ mux_left_track_37.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_11.mux_l2_in_0_ _058_/HI mux_bottom_track_11.mux_l1_in_0_/X mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l2_in_0_/X
+ _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_bottom_track_1.mux_l1_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_37.mux_l2_in_0_/S mux_left_track_39.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X
+ _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_7.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_7.mux_l1_in_1_/S
+ mux_bottom_track_7.mux_l2_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_7.mux_l2_in_1_ _035_/HI chanx_left_in[4] mux_bottom_track_7.mux_l2_in_0_/S
+ mux_bottom_track_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_087_ _087_/A chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_37.mux_l1_in_0_ left_bottom_grid_pin_39_ chany_bottom_in[17] mux_left_track_37.mux_l1_in_0_/S
+ mux_left_track_37.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_11.mux_l1_in_0_ chanx_left_in[6] bottom_left_grid_pin_42_ mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_23.mux_l2_in_0_ _064_/HI mux_bottom_track_23.mux_l1_in_0_/X mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_5.mux_l3_in_0_/S
+ mux_bottom_track_7.mux_l1_in_1_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_0_/S mux_bottom_track_7.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_086_ _086_/A chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X _091_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_069_ _069_/HI _069_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_7.mux_l1_in_1_ bottom_left_grid_pin_48_ bottom_left_grid_pin_46_
+ mux_bottom_track_7.mux_l1_in_1_/S mux_bottom_track_7.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l2_in_0_/X _086_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_6_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_23.mux_l1_in_0_ chanx_left_in[12] bottom_left_grid_pin_48_ mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_15.mux_l1_in_0_/S
+ mux_bottom_track_15.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_085_ _085_/A chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X _109_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_068_ _068_/HI _068_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_7.mux_l1_in_0_ bottom_left_grid_pin_44_ bottom_left_grid_pin_42_
+ mux_bottom_track_7.mux_l1_in_1_/S mux_bottom_track_7.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_1.mux_l2_in_1_ _037_/HI mux_left_track_1.mux_l1_in_2_/X mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_2_ left_bottom_grid_pin_41_ left_bottom_grid_pin_39_ mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l1_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X _075_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_084_ _084_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_23.mux_l2_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X _078_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_067_ _067_/HI _067_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_0 SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_1_ left_bottom_grid_pin_37_ left_bottom_grid_pin_35_ mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_083_ _083_/A chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_6_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_066_ _066_/HI _066_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_19.mux_l2_in_0_ _042_/HI mux_left_track_19.mux_l1_in_0_/X mux_left_track_19.mux_l2_in_0_/S
+ mux_left_track_19.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_21.mux_l2_in_0_ _043_/HI mux_left_track_21.mux_l1_in_0_/X mux_left_track_21.mux_l2_in_0_/S
+ mux_left_track_21.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 bottom_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[19] mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_082_ _082_/A chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_3_5_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ _065_/HI _065_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_11.mux_l1_in_0_/S mux_left_track_11.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_19.mux_l1_in_0_ left_bottom_grid_pin_38_ chany_bottom_in[8] mux_left_track_19.mux_l1_in_0_/S
+ mux_left_track_19.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_21.mux_l1_in_0_ left_bottom_grid_pin_39_ chany_bottom_in[9] mux_left_track_21.mux_l1_in_0_/S
+ mux_left_track_21.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l2_in_0_ _050_/HI mux_left_track_33.mux_l1_in_0_/X mux_left_track_33.mux_l2_in_0_/S
+ mux_left_track_33.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X
+ _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_081_ _081_/A chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_5.mux_l1_in_0_/S mux_left_track_5.mux_l2_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X
+ _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_064_ _064_/HI _064_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_9.mux_l2_in_0_/S mux_left_track_11.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l2_in_1_ _068_/HI chanx_left_in[2] mux_bottom_track_3.mux_l2_in_1_/S
+ mux_bottom_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ _080_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_3.mux_l3_in_0_/S mux_left_track_5.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l1_in_0_ left_bottom_grid_pin_37_ chany_bottom_in[15] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_063_ _063_/HI _063_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_0_ _061_/HI mux_bottom_track_17.mux_l1_in_0_/X mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_4 chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_1_/S mux_bottom_track_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

