* NGSPICE file created from cbx_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt cbx_1__0_ bottom_grid_pin_0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ prog_clk top_grid_pin_16_ top_grid_pin_17_ top_grid_pin_18_ top_grid_pin_19_ top_grid_pin_20_
+ top_grid_pin_21_ top_grid_pin_22_ top_grid_pin_23_ top_grid_pin_24_ top_grid_pin_25_
+ top_grid_pin_26_ top_grid_pin_27_ top_grid_pin_28_ top_grid_pin_29_ top_grid_pin_30_
+ top_grid_pin_31_ vpwr vgnd
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__D mux_bottom_ipin_15.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_1__S mux_top_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_26_30 vgnd vpwr scs8hd_fill_1
XFILLER_9_159 vgnd vpwr scs8hd_fill_1
XFILLER_13_155 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_12.mux_l2_in_3_ _25_/HI chanx_right_in[16] mux_bottom_ipin_12.mux_l2_in_2_/S
+ mux_bottom_ipin_12.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_280 vgnd vpwr scs8hd_decap_12
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_bottom_ipin_7.mux_l2_in_3_/S
+ mux_bottom_ipin_7.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_169 vgnd vpwr scs8hd_fill_1
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XFILLER_12_65 vgnd vpwr scs8hd_fill_1
XFILLER_18_203 vpwr vgnd scs8hd_fill_2
XFILLER_33_206 vgnd vpwr scs8hd_fill_1
XFILLER_18_269 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
X_66_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_17_291 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S mux_bottom_ipin_4.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__D mux_bottom_ipin_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_86 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_15.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_15.mux_l3_in_0_/S mux_bottom_ipin_15.mux_l4_in_0_/S
+ mem_bottom_ipin_15.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_88 vgnd vpwr scs8hd_decap_12
XFILLER_9_11 vpwr vgnd scs8hd_fill_2
X_49_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_20_231 vpwr vgnd scs8hd_fill_2
XFILLER_20_297 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_12.mux_l4_in_0_ mux_bottom_ipin_12.mux_l3_in_1_/X mux_bottom_ipin_12.mux_l3_in_0_/X
+ mux_bottom_ipin_12.mux_l4_in_0_/S mux_bottom_ipin_12.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_2.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_2.mux_l1_in_0_/X
+ mux_bottom_ipin_2.mux_l2_in_0_/S mux_bottom_ipin_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_97 vpwr vgnd scs8hd_fill_2
XFILLER_11_231 vgnd vpwr scs8hd_decap_12
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XFILLER_22_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S mux_bottom_ipin_13.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S mux_bottom_ipin_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_10.scs8hd_buf_4_0_ mux_bottom_ipin_10.mux_l4_in_0_/X top_grid_pin_26_
+ vgnd vpwr scs8hd_buf_1
XFILLER_29_96 vgnd vpwr scs8hd_decap_3
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_293 vgnd vpwr scs8hd_decap_6
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_12.mux_l3_in_1_ mux_bottom_ipin_12.mux_l2_in_3_/X mux_bottom_ipin_12.mux_l2_in_2_/X
+ mux_bottom_ipin_12.mux_l3_in_1_/S mux_bottom_ipin_12.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S mux_bottom_ipin_9.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_15_87 vpwr vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_31_123 vgnd vpwr scs8hd_fill_1
XFILLER_31_101 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1 mux_bottom_ipin_15.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_101 vgnd vpwr scs8hd_decap_4
XFILLER_22_145 vgnd vpwr scs8hd_decap_4
XFILLER_22_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0 _31_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S mux_bottom_ipin_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__D mux_bottom_ipin_2.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_ipin_12.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[12] mux_bottom_ipin_12.mux_l2_in_2_/S
+ mux_bottom_ipin_12.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0 mux_bottom_ipin_6.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_7.mux_l1_in_0_/X
+ mux_bottom_ipin_7.mux_l2_in_3_/S mux_bottom_ipin_7.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_204 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S mux_bottom_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_292 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XFILLER_18_237 vpwr vgnd scs8hd_fill_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
X_65_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_32_273 vpwr vgnd scs8hd_fill_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_5.mux_l3_in_1_/S mux_bottom_ipin_5.mux_l4_in_0_/S
+ mem_bottom_ipin_5.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S mux_bottom_ipin_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S mux_bottom_ipin_1.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_65 vpwr vgnd scs8hd_fill_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_15.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_15.mux_l2_in_3_/S mux_bottom_ipin_15.mux_l3_in_0_/S
+ mem_bottom_ipin_15.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_23 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.scs8hd_buf_4_0_ mux_bottom_ipin_7.mux_l4_in_0_/X top_grid_pin_23_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_48_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S mux_bottom_ipin_7.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l3_in_0__A0 mux_top_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_210 vpwr vgnd scs8hd_fill_2
XFILLER_20_265 vgnd vpwr scs8hd_decap_3
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XFILLER_11_210 vpwr vgnd scs8hd_fill_2
XFILLER_11_243 vgnd vpwr scs8hd_fill_1
XFILLER_7_269 vgnd vpwr scs8hd_decap_6
XFILLER_15_7 vgnd vpwr scs8hd_decap_4
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0 mux_bottom_ipin_10.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_75 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__D mux_bottom_ipin_3.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_19_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_14.scs8hd_buf_4_0__A mux_bottom_ipin_14.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_12.mux_l3_in_0_ mux_bottom_ipin_12.mux_l2_in_1_/X mux_bottom_ipin_12.mux_l2_in_0_/X
+ mux_bottom_ipin_12.mux_l3_in_1_/S mux_bottom_ipin_12.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_2.mux_l1_in_0_/S
+ mux_bottom_ipin_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_165 vpwr vgnd scs8hd_fill_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_31_65 vgnd vpwr scs8hd_decap_12
XFILLER_31_21 vpwr vgnd scs8hd_fill_2
XFILLER_31_87 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_3
XFILLER_16_176 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vpwr vgnd scs8hd_fill_2
XFILLER_22_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_26_65 vgnd vpwr scs8hd_decap_4
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1 mux_bottom_ipin_6.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_12.mux_l2_in_1_ chanx_left_in[12] mux_bottom_ipin_12.mux_l1_in_2_/X
+ mux_bottom_ipin_12.mux_l2_in_2_/S mux_bottom_ipin_12.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_290 vpwr vgnd scs8hd_fill_2
XFILLER_8_172 vgnd vpwr scs8hd_decap_12
XFILLER_12_190 vgnd vpwr scs8hd_fill_1
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A1 mux_top_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_271 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
X_64_ chanx_left_in[9] chanx_right_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_32_285 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S mux_bottom_ipin_15.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_5.mux_l2_in_3_/S mux_bottom_ipin_5.mux_l3_in_1_/S
+ mem_bottom_ipin_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_296 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_12.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_bottom_ipin_12.mux_l1_in_2_/S
+ mux_bottom_ipin_12.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_22 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__D mux_bottom_ipin_5.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_15.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_15.mux_l1_in_0_/S mux_bottom_ipin_15.mux_l2_in_3_/S
+ mem_bottom_ipin_15.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_ipin_7.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_7.mux_l1_in_0_/S
+ mux_bottom_ipin_7.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_14_285 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.scs8hd_buf_4_0__A mux_bottom_ipin_6.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
X_47_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_0.mux_l3_in_0__A1 mux_top_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_244 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S mux_bottom_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S mux_bottom_ipin_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1 mux_bottom_ipin_10.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_54 vgnd vpwr scs8hd_decap_4
XFILLER_34_166 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0 mux_bottom_ipin_1.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_177 vgnd vpwr scs8hd_decap_4
XFILLER_25_100 vgnd vpwr scs8hd_decap_3
XFILLER_31_77 vgnd vpwr scs8hd_decap_6
XFILLER_31_55 vpwr vgnd scs8hd_fill_2
XFILLER_0_298 vgnd vpwr scs8hd_fill_1
XFILLER_31_169 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vgnd vpwr scs8hd_decap_3
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S mux_bottom_ipin_13.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S mux_bottom_ipin_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_44 vpwr vgnd scs8hd_fill_2
XFILLER_26_88 vpwr vgnd scs8hd_fill_2
XFILLER_13_147 vgnd vpwr scs8hd_decap_8
XFILLER_13_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_12.mux_l2_in_0_ mux_bottom_ipin_12.mux_l1_in_1_/X mux_bottom_ipin_12.mux_l1_in_0_/X
+ mux_bottom_ipin_12.mux_l2_in_2_/S mux_bottom_ipin_12.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__D mux_bottom_ipin_7.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_261 vgnd vpwr scs8hd_decap_12
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.scs8hd_buf_4_0_ mux_bottom_ipin_2.mux_l4_in_0_/X top_grid_pin_18_
+ vgnd vpwr scs8hd_buf_1
XFILLER_5_7 vgnd vpwr scs8hd_decap_12
XFILLER_12_24 vgnd vpwr scs8hd_decap_4
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_24_209 vgnd vpwr scs8hd_decap_3
X_63_ chanx_left_in[10] chanx_right_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_297 vpwr vgnd scs8hd_fill_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_5.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_5.mux_l1_in_0_/S mux_bottom_ipin_5.mux_l2_in_3_/S
+ mem_bottom_ipin_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S mux_bottom_ipin_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S mux_bottom_ipin_12.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_275 vgnd vpwr scs8hd_fill_1
XFILLER_23_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S mux_bottom_ipin_4.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_12.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_12.mux_l1_in_2_/S
+ mux_bottom_ipin_12.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_15.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_14.mux_l4_in_0_/S mux_bottom_ipin_15.mux_l1_in_0_/S
+ mem_bottom_ipin_15.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_47 vgnd vpwr scs8hd_decap_4
XFILLER_14_297 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
X_46_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_20_289 vgnd vpwr scs8hd_decap_8
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_3
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_18_78 vgnd vpwr scs8hd_decap_4
XFILLER_18_89 vgnd vpwr scs8hd_decap_3
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XFILLER_11_267 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1 mux_bottom_ipin_1.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
X_29_ _29_/HI _29_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S mux_bottom_ipin_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_33 vpwr vgnd scs8hd_fill_2
XFILLER_29_11 vpwr vgnd scs8hd_fill_2
XFILLER_20_46 vgnd vpwr scs8hd_decap_3
XFILLER_20_57 vgnd vpwr scs8hd_decap_4
XFILLER_28_131 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_10.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_10.mux_l3_in_1_/S mux_bottom_ipin_10.mux_l4_in_0_/S
+ mem_bottom_ipin_10.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__D mux_bottom_ipin_10.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0 mux_bottom_ipin_8.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__D mux_bottom_ipin_8.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_8
XFILLER_34_123 vpwr vgnd scs8hd_fill_2
XFILLER_19_142 vgnd vpwr scs8hd_decap_4
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S mux_bottom_ipin_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1 mux_bottom_ipin_1.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_13 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_112 vgnd vpwr scs8hd_decap_4
XFILLER_16_189 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0 mux_bottom_ipin_8.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_23 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_8_196 vpwr vgnd scs8hd_fill_2
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XFILLER_35_273 vgnd vpwr scs8hd_decap_6
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_36 vgnd vpwr scs8hd_decap_3
XFILLER_12_58 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_207 vgnd vpwr scs8hd_decap_4
XFILLER_26_251 vgnd vpwr scs8hd_decap_4
XFILLER_26_240 vpwr vgnd scs8hd_fill_2
X_62_ chanx_left_in[11] chanx_right_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_17_262 vpwr vgnd scs8hd_fill_2
XFILLER_32_265 vgnd vpwr scs8hd_decap_8
XFILLER_17_295 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_5.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_4.mux_l4_in_0_/S mux_bottom_ipin_5.mux_l1_in_0_/S
+ mem_bottom_ipin_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0 mux_bottom_ipin_12.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_12.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_12.mux_l1_in_2_/S
+ mux_bottom_ipin_12.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_35 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
XFILLER_14_243 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__D mux_bottom_ipin_11.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__D mux_bottom_ipin_9.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
X_45_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_9_291 vpwr vgnd scs8hd_fill_2
XFILLER_18_46 vgnd vpwr scs8hd_fill_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S mux_bottom_ipin_11.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_279 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0 mux_bottom_ipin_12.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_0.mux_l3_in_0_/S mux_bottom_ipin_0.mux_l4_in_0_/S
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
X_28_ _28_/HI _28_/LO vgnd vpwr scs8hd_conb_1
Xmem_bottom_ipin_10.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_10.mux_l2_in_3_/S mux_bottom_ipin_10.mux_l3_in_1_/S
+ mem_bottom_ipin_10.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_89 vgnd vpwr scs8hd_decap_4
XFILLER_28_154 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1 mux_bottom_ipin_8.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_19_132 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.scs8hd_buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X bottom_grid_pin_0_ vgnd
+ vpwr scs8hd_buf_1
Xmux_bottom_ipin_3.mux_l2_in_3_ _30_/HI chanx_right_in[15] mux_bottom_ipin_3.mux_l2_in_2_/S
+ mux_bottom_ipin_3.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1 mux_bottom_ipin_14.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S mux_bottom_ipin_10.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_127 vpwr vgnd scs8hd_fill_2
XFILLER_22_149 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0 mux_bottom_ipin_5.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1 mux_bottom_ipin_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__D mux_bottom_ipin_12.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_193 vpwr vgnd scs8hd_fill_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_26_285 vgnd vpwr scs8hd_decap_12
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S mux_bottom_ipin_1.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_61_ chanx_left_in[12] chanx_right_out[12] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_3.mux_l4_in_0_ mux_bottom_ipin_3.mux_l3_in_1_/X mux_bottom_ipin_3.mux_l3_in_0_/X
+ mux_bottom_ipin_3.mux_l4_in_0_/S mux_bottom_ipin_3.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S mux_bottom_ipin_15.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1 mux_bottom_ipin_12.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_288 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l4_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_23_69 vpwr vgnd scs8hd_fill_2
XFILLER_14_255 vgnd vpwr scs8hd_decap_8
X_44_ chanx_right_in[9] chanx_left_out[9] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0 mux_bottom_ipin_3.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_8.mux_l2_in_3_ _18_/HI chanx_right_in[18] mux_bottom_ipin_8.mux_l2_in_3_/S
+ mux_bottom_ipin_8.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_36 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S mux_bottom_ipin_10.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l3_in_1_ mux_bottom_ipin_3.mux_l2_in_3_/X mux_bottom_ipin_3.mux_l2_in_2_/X
+ mux_bottom_ipin_3.mux_l3_in_1_/S mux_bottom_ipin_3.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S mux_bottom_ipin_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1 mux_bottom_ipin_12.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XFILLER_10_280 vgnd vpwr scs8hd_decap_12
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_0.mux_l2_in_1_/S mux_bottom_ipin_0.mux_l3_in_0_/S
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
X_27_ _27_/HI _27_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S mux_bottom_ipin_14.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_10.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_10.mux_l1_in_0_/S mux_bottom_ipin_10.mux_l2_in_3_/S
+ mem_bottom_ipin_10.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__34__A chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.scs8hd_buf_4_0__A mux_bottom_ipin_1.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0 mux_bottom_ipin_3.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_10_70 vpwr vgnd scs8hd_fill_2
XFILLER_10_81 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__D mux_bottom_ipin_14.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_169 vpwr vgnd scs8hd_fill_2
XFILLER_25_136 vgnd vpwr scs8hd_decap_4
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_26 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_bottom_ipin_3.mux_l2_in_2_/S
+ mux_bottom_ipin_3.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_8.mux_l4_in_0_ mux_bottom_ipin_8.mux_l3_in_1_/X mux_bottom_ipin_8.mux_l3_in_0_/X
+ mux_bottom_ipin_8.mux_l4_in_0_/S mux_bottom_ipin_8.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_12
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1 mux_bottom_ipin_5.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S mux_bottom_ipin_5.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_294 vgnd vpwr scs8hd_decap_4
XFILLER_29_250 vpwr vgnd scs8hd_fill_2
XFILLER_8_154 vgnd vpwr scs8hd_fill_1
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XFILLER_32_90 vpwr vgnd scs8hd_fill_2
XFILLER_27_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D mux_bottom_ipin_0.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_242 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S mux_bottom_ipin_9.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_8.mux_l3_in_1_ mux_bottom_ipin_8.mux_l2_in_3_/X mux_bottom_ipin_8.mux_l2_in_2_/X
+ mux_bottom_ipin_8.mux_l3_in_1_/S mux_bottom_ipin_8.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_297 vpwr vgnd scs8hd_fill_2
XANTENNA__42__A chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_1__D mux_top_ipin_0.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
X_60_ chanx_left_in[13] chanx_right_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_32_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_278 vgnd vpwr scs8hd_fill_1
XFILLER_23_245 vgnd vpwr scs8hd_decap_4
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA__37__A chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_14_267 vgnd vpwr scs8hd_decap_6
X_43_ chanx_right_in[10] chanx_left_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_215 vgnd vpwr scs8hd_decap_3
XFILLER_20_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1 mux_bottom_ipin_3.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_8.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_bottom_ipin_8.mux_l2_in_3_/S
+ mux_bottom_ipin_8.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S mux_bottom_ipin_8.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.mux_l3_in_0_ mux_bottom_ipin_3.mux_l2_in_1_/X mux_bottom_ipin_3.mux_l2_in_0_/X
+ mux_bottom_ipin_3.mux_l3_in_1_/S mux_bottom_ipin_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_ipin_8.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_8.mux_l3_in_1_/S mux_bottom_ipin_8.mux_l4_in_0_/S
+ mem_bottom_ipin_8.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_296 vgnd vpwr scs8hd_decap_3
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
XFILLER_10_292 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_0.mux_l1_in_2_/S mux_bottom_ipin_0.mux_l2_in_1_/S
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
X_26_ _26_/HI _26_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_58 vgnd vpwr scs8hd_fill_1
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XFILLER_28_123 vpwr vgnd scs8hd_fill_2
XFILLER_28_112 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_10.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_9.mux_l4_in_0_/S mux_bottom_ipin_10.mux_l1_in_0_/S
+ mem_bottom_ipin_10.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0 _27_/HI vgnd vpwr scs8hd_diode_2
XFILLER_6_29 vpwr vgnd scs8hd_fill_2
XANTENNA__50__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1 mux_bottom_ipin_3.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0 mux_bottom_ipin_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__D mux_bottom_ipin_2.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_3.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_bottom_ipin_3.mux_l2_in_2_/S
+ mux_bottom_ipin_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_137 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_159 vpwr vgnd scs8hd_fill_2
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__45__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_107 vgnd vpwr scs8hd_fill_1
XFILLER_26_26 vpwr vgnd scs8hd_fill_2
XFILLER_26_15 vpwr vgnd scs8hd_fill_2
XFILLER_29_273 vgnd vpwr scs8hd_decap_3
XFILLER_16_70 vpwr vgnd scs8hd_fill_2
XFILLER_35_298 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_28 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_8.mux_l3_in_0_ mux_bottom_ipin_8.mux_l2_in_1_/X mux_bottom_ipin_8.mux_l2_in_0_/X
+ mux_bottom_ipin_8.mux_l3_in_1_/S mux_bottom_ipin_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S mux_bottom_ipin_12.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_287 vpwr vgnd scs8hd_fill_2
XFILLER_23_202 vpwr vgnd scs8hd_fill_2
XFILLER_31_290 vpwr vgnd scs8hd_fill_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_13.mux_l2_in_3_ _26_/HI chanx_right_in[17] mux_bottom_ipin_13.mux_l2_in_2_/S
+ mux_bottom_ipin_13.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__53__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_224 vgnd vpwr scs8hd_decap_12
XFILLER_13_82 vpwr vgnd scs8hd_fill_2
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
X_42_ chanx_right_in[11] chanx_left_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_227 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_8.mux_l2_in_1_ chanx_left_in[12] mux_bottom_ipin_8.mux_l1_in_2_/X
+ mux_bottom_ipin_8.mux_l2_in_3_/S mux_bottom_ipin_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_283 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__D mux_bottom_ipin_3.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_8.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_8.mux_l2_in_3_/S mux_bottom_ipin_8.mux_l3_in_1_/S
+ mem_bottom_ipin_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_227 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_11.scs8hd_buf_4_0_ mux_bottom_ipin_11.mux_l4_in_0_/X top_grid_pin_27_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S mux_bottom_ipin_11.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__48__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_bottom_ipin_0.mux_l1_in_2_/S
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
X_25_ _25_/HI _25_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.scs8hd_buf_4_0__A mux_bottom_ipin_9.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S mux_bottom_ipin_7.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_37 vpwr vgnd scs8hd_fill_2
XFILLER_28_179 vgnd vpwr scs8hd_decap_6
XFILLER_28_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1 mux_bottom_ipin_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_19_102 vgnd vpwr scs8hd_decap_3
XFILLER_34_127 vgnd vpwr scs8hd_decap_12
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_146 vgnd vpwr scs8hd_fill_1
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_8.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_bottom_ipin_8.mux_l1_in_0_/S
+ mux_bottom_ipin_8.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_3.mux_l1_in_0_/X
+ mux_bottom_ipin_3.mux_l2_in_2_/S mux_bottom_ipin_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_13.mux_l4_in_0_ mux_bottom_ipin_13.mux_l3_in_1_/X mux_bottom_ipin_13.mux_l3_in_0_/X
+ mux_bottom_ipin_13.mux_l4_in_0_/S mux_bottom_ipin_13.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0 _32_/HI vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S mux_bottom_ipin_10.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_119 vgnd vpwr scs8hd_decap_3
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_182 vpwr vgnd scs8hd_fill_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__61__A chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0 mux_bottom_ipin_7.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XFILLER_30_130 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vgnd vpwr scs8hd_decap_4
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S mux_bottom_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_163 vgnd vpwr scs8hd_decap_3
XANTENNA__56__A chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_4
XFILLER_32_70 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_13.mux_l3_in_1_ mux_bottom_ipin_13.mux_l2_in_3_/X mux_bottom_ipin_13.mux_l2_in_2_/X
+ mux_bottom_ipin_13.mux_l3_in_1_/S mux_bottom_ipin_13.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XFILLER_12_18 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__D mux_bottom_ipin_4.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S mux_bottom_ipin_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_8.scs8hd_buf_4_0_ mux_bottom_ipin_8.mux_l4_in_0_/X top_grid_pin_24_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_3
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S mux_bottom_ipin_5.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_13.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[13] mux_bottom_ipin_13.mux_l2_in_2_/S
+ mux_bottom_ipin_13.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_19 vpwr vgnd scs8hd_fill_2
XFILLER_14_236 vpwr vgnd scs8hd_fill_2
XFILLER_14_247 vpwr vgnd scs8hd_fill_2
X_41_ chanx_right_in[12] chanx_left_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_9_295 vgnd vpwr scs8hd_decap_4
XFILLER_13_291 vpwr vgnd scs8hd_fill_2
XFILLER_20_206 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_8.mux_l2_in_0_ mux_bottom_ipin_8.mux_l1_in_1_/X mux_bottom_ipin_8.mux_l1_in_0_/X
+ mux_bottom_ipin_8.mux_l2_in_3_/S mux_bottom_ipin_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_8.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_8.mux_l1_in_0_/S mux_bottom_ipin_8.mux_l2_in_3_/S
+ mem_bottom_ipin_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0 mux_bottom_ipin_11.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__64__A chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_6_276 vgnd vpwr scs8hd_decap_12
XFILLER_10_272 vgnd vpwr scs8hd_decap_3
X_24_ _24_/HI _24_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S mux_bottom_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S mux_bottom_ipin_4.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XANTENNA__59__A chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_8.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_8.mux_l1_in_0_/S
+ mux_bottom_ipin_8.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_139 vgnd vpwr scs8hd_decap_12
XFILLER_34_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_19_158 vpwr vgnd scs8hd_fill_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_194 vpwr vgnd scs8hd_fill_2
XFILLER_33_172 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__D mux_bottom_ipin_6.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1 mux_bottom_ipin_7.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_13.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_13.mux_l3_in_1_/S mux_bottom_ipin_13.mux_l4_in_0_/S
+ mem_bottom_ipin_13.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_21_83 vgnd vpwr scs8hd_decap_3
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_161 vpwr vgnd scs8hd_fill_2
XFILLER_30_186 vpwr vgnd scs8hd_fill_2
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_26_39 vgnd vpwr scs8hd_decap_3
XFILLER_21_142 vpwr vgnd scs8hd_fill_2
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_231 vpwr vgnd scs8hd_fill_2
XANTENNA__72__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_83 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_82 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_13.mux_l3_in_0_ mux_bottom_ipin_13.mux_l2_in_1_/X mux_bottom_ipin_13.mux_l2_in_0_/X
+ mux_bottom_ipin_13.mux_l3_in_1_/S mux_bottom_ipin_13.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_168 vpwr vgnd scs8hd_fill_2
XFILLER_12_186 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_3.mux_l1_in_0_/S
+ mux_bottom_ipin_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_267 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_1__S mux_top_ipin_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA__67__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_17_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vpwr vgnd scs8hd_fill_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_215 vpwr vgnd scs8hd_fill_2
XFILLER_23_18 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_13.mux_l2_in_1_ chanx_left_in[13] mux_bottom_ipin_13.mux_l1_in_2_/X
+ mux_bottom_ipin_13.mux_l2_in_2_/S mux_bottom_ipin_13.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_62 vgnd vpwr scs8hd_fill_1
X_40_ chanx_right_in[13] chanx_left_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1 mux_bottom_ipin_11.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__D mux_bottom_ipin_8.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_8.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_7.mux_l4_in_0_/S mux_bottom_ipin_8.mux_l1_in_0_/S
+ mem_bottom_ipin_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0 _21_/HI vgnd vpwr scs8hd_diode_2
XFILLER_10_240 vgnd vpwr scs8hd_decap_12
XFILLER_6_288 vgnd vpwr scs8hd_decap_8
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
X_23_ _23_/HI _23_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0 mux_bottom_ipin_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_13.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_bottom_ipin_13.mux_l1_in_2_/S
+ mux_bottom_ipin_13.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_269 vgnd vpwr scs8hd_decap_12
XFILLER_10_41 vgnd vpwr scs8hd_decap_12
XFILLER_10_74 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_8.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_8.mux_l1_in_0_/S
+ mux_bottom_ipin_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_170 vpwr vgnd scs8hd_fill_2
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_18_170 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_3.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_3.mux_l3_in_1_/S mux_bottom_ipin_3.mux_l4_in_0_/S
+ mem_bottom_ipin_3.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S mux_bottom_ipin_13.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S mux_bottom_ipin_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_173 vpwr vgnd scs8hd_fill_2
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_13.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_13.mux_l2_in_2_/S mux_bottom_ipin_13.mux_l3_in_1_/S
+ mem_bottom_ipin_13.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_151 vgnd vpwr scs8hd_decap_4
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.scs8hd_buf_4_0_ mux_bottom_ipin_3.mux_l4_in_0_/X top_grid_pin_19_
+ vgnd vpwr scs8hd_buf_1
XFILLER_29_298 vgnd vpwr scs8hd_fill_1
XFILLER_29_243 vgnd vpwr scs8hd_fill_1
XFILLER_29_210 vgnd vpwr scs8hd_decap_4
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_40 vpwr vgnd scs8hd_fill_2
XFILLER_8_158 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__D mux_bottom_ipin_11.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_257 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S mux_bottom_ipin_12.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S mux_bottom_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_32_205 vgnd vpwr scs8hd_decap_8
XFILLER_17_224 vpwr vgnd scs8hd_fill_2
XFILLER_17_279 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.scs8hd_buf_4_0__A mux_bottom_ipin_12.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_23_249 vgnd vpwr scs8hd_fill_1
XFILLER_23_238 vpwr vgnd scs8hd_fill_2
XFILLER_31_282 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S mux_bottom_ipin_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_13.mux_l2_in_0_ mux_bottom_ipin_13.mux_l1_in_1_/X mux_bottom_ipin_13.mux_l1_in_0_/X
+ mux_bottom_ipin_13.mux_l2_in_2_/S mux_bottom_ipin_13.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_22_271 vpwr vgnd scs8hd_fill_2
XFILLER_13_271 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0 mux_bottom_ipin_9.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S mux_bottom_ipin_1.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XFILLER_10_252 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_1_11 vgnd vpwr scs8hd_decap_12
X_22_ _22_/HI _22_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1 mux_bottom_ipin_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_127 vpwr vgnd scs8hd_fill_2
XFILLER_28_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S mux_bottom_ipin_7.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_13.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_13.mux_l1_in_2_/S
+ mux_bottom_ipin_13.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S mux_bottom_ipin_15.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_10_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_3
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
XFILLER_33_152 vgnd vpwr scs8hd_decap_12
XFILLER_18_193 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_3.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_3.mux_l2_in_2_/S mux_bottom_ipin_3.mux_l3_in_1_/S
+ mem_bottom_ipin_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0 mux_bottom_ipin_9.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__D mux_bottom_ipin_12.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_16_108 vpwr vgnd scs8hd_fill_2
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_13.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_13.mux_l1_in_2_/S mux_bottom_ipin_13.mux_l2_in_2_/S
+ mem_bottom_ipin_13.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S mux_bottom_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S mux_bottom_ipin_0.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.scs8hd_buf_4_0__A mux_bottom_ipin_4.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_166 vgnd vpwr scs8hd_fill_1
XFILLER_30_144 vgnd vpwr scs8hd_decap_6
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_26_19 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S mux_bottom_ipin_6.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0 mux_bottom_ipin_13.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_247 vpwr vgnd scs8hd_fill_2
XFILLER_26_236 vpwr vgnd scs8hd_fill_2
XFILLER_34_291 vgnd vpwr scs8hd_decap_8
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XFILLER_25_291 vpwr vgnd scs8hd_fill_2
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_31_294 vgnd vpwr scs8hd_decap_4
XFILLER_14_206 vpwr vgnd scs8hd_fill_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0 mux_bottom_ipin_13.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
XFILLER_13_283 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__D mux_bottom_ipin_13.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1 mux_bottom_ipin_9.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_41 vgnd vpwr scs8hd_decap_3
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.scs8hd_buf_4_0__A mux_top_ipin_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_220 vpwr vgnd scs8hd_fill_2
XFILLER_10_264 vgnd vpwr scs8hd_decap_8
XFILLER_1_23 vgnd vpwr scs8hd_decap_12
X_21_ _21_/HI _21_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_ipin_13.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_13.mux_l1_in_2_/S
+ mux_bottom_ipin_13.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1 mux_bottom_ipin_15.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_74 vpwr vgnd scs8hd_fill_2
XFILLER_33_164 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_3.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_3.mux_l1_in_0_/S mux_bottom_ipin_3.mux_l2_in_2_/S
+ mem_bottom_ipin_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1 mux_bottom_ipin_9.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S mux_bottom_ipin_14.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_13.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_12.mux_l4_in_0_/S mux_bottom_ipin_13.mux_l1_in_2_/S
+ mem_bottom_ipin_13.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_134 vgnd vpwr scs8hd_decap_8
XFILLER_7_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_101 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_29_278 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_41 vgnd vpwr scs8hd_fill_1
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1 mux_bottom_ipin_13.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_3_ _31_/HI chanx_right_in[14] mux_bottom_ipin_4.mux_l2_in_2_/S
+ mux_bottom_ipin_4.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S mux_bottom_ipin_13.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__D mux_bottom_ipin_15.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_2__S mux_top_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_27_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0__A0 mux_top_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_74 vpwr vgnd scs8hd_fill_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0 mux_bottom_ipin_4.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_240 vpwr vgnd scs8hd_fill_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1 mux_bottom_ipin_13.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_211 vgnd vpwr scs8hd_decap_12
XFILLER_13_295 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S mux_bottom_ipin_4.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S mux_bottom_ipin_12.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_75 vpwr vgnd scs8hd_fill_2
XFILLER_10_210 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__D mux_bottom_ipin_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_298 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0 mux_bottom_ipin_4.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l4_in_0_ mux_bottom_ipin_4.mux_l3_in_1_/X mux_bottom_ipin_4.mux_l3_in_0_/X
+ mux_bottom_ipin_4.mux_l4_in_0_/S mux_bottom_ipin_4.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_35 vgnd vpwr scs8hd_decap_12
X_20_ _20_/HI _20_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_22 vpwr vgnd scs8hd_fill_2
XFILLER_10_66 vpwr vgnd scs8hd_fill_2
XFILLER_19_42 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_9.mux_l2_in_3_ _19_/HI chanx_right_in[19] mux_bottom_ipin_9.mux_l2_in_0_/S
+ mux_bottom_ipin_9.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
XFILLER_33_198 vpwr vgnd scs8hd_fill_2
XFILLER_33_176 vgnd vpwr scs8hd_fill_1
XFILLER_33_132 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_3.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_2.mux_l4_in_0_/S mux_bottom_ipin_3.mux_l1_in_0_/S
+ mem_bottom_ipin_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1 mux_bottom_ipin_6.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S mux_bottom_ipin_13.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_4.mux_l3_in_1_ mux_bottom_ipin_4.mux_l2_in_3_/X mux_bottom_ipin_4.mux_l2_in_2_/X
+ mux_bottom_ipin_4.mux_l3_in_1_/S mux_bottom_ipin_4.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S mux_bottom_ipin_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S mux_bottom_ipin_11.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_23 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S mux_bottom_ipin_9.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_146 vpwr vgnd scs8hd_fill_2
XFILLER_21_168 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_87 vpwr vgnd scs8hd_fill_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XFILLER_20_190 vgnd vpwr scs8hd_decap_4
XFILLER_35_249 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_bottom_ipin_4.mux_l2_in_2_/S
+ mux_bottom_ipin_4.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_205 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_9.mux_l4_in_0_ mux_bottom_ipin_9.mux_l3_in_1_/X mux_bottom_ipin_9.mux_l3_in_0_/X
+ mux_bottom_ipin_9.mux_l4_in_0_/S mux_bottom_ipin_9.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S mux_bottom_ipin_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0__A1 mux_top_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__D mux_bottom_ipin_3.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_23_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1 mux_bottom_ipin_4.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S mux_bottom_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_285 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1 mux_bottom_ipin_10.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_223 vgnd vpwr scs8hd_decap_12
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XFILLER_13_241 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_9.mux_l3_in_1_ mux_bottom_ipin_9.mux_l2_in_3_/X mux_bottom_ipin_9.mux_l2_in_2_/X
+ mux_bottom_ipin_9.mux_l3_in_1_/S mux_bottom_ipin_9.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0 _28_/HI vgnd vpwr scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0 mux_bottom_ipin_1.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1 mux_bottom_ipin_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_47 vgnd vpwr scs8hd_decap_12
XFILLER_10_78 vgnd vpwr scs8hd_fill_1
XFILLER_10_89 vgnd vpwr scs8hd_decap_3
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vpwr vgnd scs8hd_fill_2
XFILLER_27_174 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_9.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_bottom_ipin_9.mux_l2_in_0_/S
+ mux_bottom_ipin_9.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_144 vgnd vpwr scs8hd_fill_1
XFILLER_24_177 vgnd vpwr scs8hd_decap_3
XFILLER_24_111 vgnd vpwr scs8hd_fill_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_4.mux_l3_in_0_ mux_bottom_ipin_4.mux_l2_in_1_/X mux_bottom_ipin_4.mux_l2_in_0_/X
+ mux_bottom_ipin_4.mux_l3_in_1_/S mux_bottom_ipin_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_11 vpwr vgnd scs8hd_fill_2
XFILLER_30_103 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__D mux_bottom_ipin_4.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_35 vgnd vpwr scs8hd_decap_12
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_214 vgnd vpwr scs8hd_fill_1
XFILLER_16_11 vgnd vpwr scs8hd_fill_1
XFILLER_16_44 vgnd vpwr scs8hd_decap_3
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_32_54 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vpwr vgnd scs8hd_fill_2
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S mux_bottom_ipin_10.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_bottom_ipin_4.mux_l1_in_2_/X
+ mux_bottom_ipin_4.mux_l2_in_2_/S mux_bottom_ipin_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_291 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_17_228 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_231 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_261 vpwr vgnd scs8hd_fill_2
XFILLER_31_286 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_12.scs8hd_buf_4_0_ mux_bottom_ipin_12.mux_l4_in_0_/X top_grid_pin_28_
+ vgnd vpwr scs8hd_buf_1
XFILLER_13_45 vpwr vgnd scs8hd_fill_2
XFILLER_22_297 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_4.mux_l1_in_1_/S
+ mux_bottom_ipin_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_235 vgnd vpwr scs8hd_decap_8
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_9_279 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_9.mux_l3_in_0_ mux_bottom_ipin_9.mux_l2_in_1_/X mux_bottom_ipin_9.mux_l2_in_0_/X
+ mux_bottom_ipin_9.mux_l3_in_1_/S mux_bottom_ipin_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_ipin_0.mux_l3_in_0__S mux_top_ipin_0.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1 mux_bottom_ipin_1.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__D mux_bottom_ipin_5.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0 _33_/HI vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_14.mux_l2_in_3_ _27_/HI chanx_right_in[18] mux_bottom_ipin_14.mux_l2_in_0_/S
+ mux_bottom_ipin_14.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S mux_bottom_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0 mux_bottom_ipin_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_9.mux_l2_in_1_ chanx_left_in[13] mux_bottom_ipin_9.mux_l1_in_2_/X
+ mux_bottom_ipin_9.mux_l2_in_0_/S mux_bottom_ipin_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_296 vgnd vpwr scs8hd_decap_3
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_142 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S mux_bottom_ipin_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_112 vgnd vpwr scs8hd_decap_4
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XFILLER_7_47 vgnd vpwr scs8hd_decap_12
XFILLER_21_159 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_6.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_6.mux_l3_in_1_/S mux_bottom_ipin_6.mux_l4_in_0_/S
+ mem_bottom_ipin_6.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_9.mux_l1_in_2_ chanx_right_in[9] chanx_left_in[9] mux_bottom_ipin_9.mux_l1_in_2_/S
+ mux_bottom_ipin_9.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_159 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A0 _20_/HI vgnd vpwr scs8hd_diode_2
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_9.scs8hd_buf_4_0_ mux_bottom_ipin_9.mux_l4_in_0_/X top_grid_pin_25_
+ vgnd vpwr scs8hd_buf_1
Xmux_bottom_ipin_14.mux_l4_in_0_ mux_bottom_ipin_14.mux_l3_in_1_/X mux_bottom_ipin_14.mux_l3_in_0_/X
+ mux_bottom_ipin_14.mux_l4_in_0_/S mux_bottom_ipin_14.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_4.mux_l2_in_0_ mux_bottom_ipin_4.mux_l1_in_1_/X mux_bottom_ipin_4.mux_l1_in_0_/X
+ mux_bottom_ipin_4.mux_l2_in_2_/S mux_bottom_ipin_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S mux_bottom_ipin_13.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S mux_bottom_ipin_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_66 vpwr vgnd scs8hd_fill_2
XFILLER_25_251 vpwr vgnd scs8hd_fill_2
XFILLER_25_295 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__D mux_bottom_ipin_7.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0 _23_/HI vgnd vpwr scs8hd_diode_2
XFILLER_31_243 vgnd vpwr scs8hd_fill_1
XFILLER_31_298 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S mux_bottom_ipin_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0 mux_bottom_ipin_12.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_210 vpwr vgnd scs8hd_fill_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_13_221 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_14.mux_l3_in_1_ mux_bottom_ipin_14.mux_l2_in_3_/X mux_bottom_ipin_14.mux_l2_in_2_/X
+ mux_bottom_ipin_14.mux_l3_in_0_/S mux_bottom_ipin_14.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_4.mux_l1_in_1_/S
+ mux_bottom_ipin_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_269 vgnd vpwr scs8hd_decap_4
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1 mux_bottom_ipin_8.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.scs8hd_buf_4_0__A mux_bottom_ipin_15.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_280 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S mux_bottom_ipin_4.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_283 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S mux_bottom_ipin_8.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_14.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_bottom_ipin_14.mux_l2_in_0_/S
+ mux_bottom_ipin_14.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_143 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vgnd vpwr scs8hd_decap_4
XFILLER_19_34 vpwr vgnd scs8hd_fill_2
XFILLER_19_78 vgnd vpwr scs8hd_decap_3
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1 mux_bottom_ipin_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_9.mux_l2_in_0_ mux_bottom_ipin_9.mux_l1_in_1_/X mux_bottom_ipin_9.mux_l1_in_0_/X
+ mux_bottom_ipin_9.mux_l2_in_0_/S mux_bottom_ipin_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vgnd vpwr scs8hd_decap_3
XFILLER_24_135 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_35 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_21_79 vpwr vgnd scs8hd_fill_2
XFILLER_15_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__D mux_bottom_ipin_10.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__D mux_bottom_ipin_9.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_190 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S mux_bottom_ipin_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S mux_bottom_ipin_7.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_6.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_6.mux_l2_in_3_/S mux_bottom_ipin_6.mux_l3_in_1_/S
+ mem_bottom_ipin_6.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_32_23 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_9.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_9.mux_l1_in_2_/S
+ mux_bottom_ipin_9.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1 mux_bottom_ipin_12.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_28_271 vgnd vpwr scs8hd_fill_1
XFILLER_28_260 vpwr vgnd scs8hd_fill_2
XFILLER_11_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.scs8hd_buf_4_0__A mux_bottom_ipin_7.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_25_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_241 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_16_285 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1 mux_bottom_ipin_12.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_14 vpwr vgnd scs8hd_fill_2
XFILLER_22_244 vpwr vgnd scs8hd_fill_2
XFILLER_8_7 vpwr vgnd scs8hd_fill_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_14.mux_l3_in_0_ mux_bottom_ipin_14.mux_l2_in_1_/X mux_bottom_ipin_14.mux_l2_in_0_/X
+ mux_bottom_ipin_14.mux_l3_in_0_/S mux_bottom_ipin_14.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0 _22_/HI vgnd vpwr scs8hd_diode_2
XFILLER_13_255 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_4.mux_l1_in_1_/S
+ mux_bottom_ipin_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0 mux_bottom_ipin_3.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_292 vgnd vpwr scs8hd_decap_6
XFILLER_24_79 vpwr vgnd scs8hd_fill_2
XFILLER_24_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__D mux_bottom_ipin_12.mux_l1_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_295 vgnd vpwr scs8hd_decap_4
XFILLER_10_26 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_14.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_bottom_ipin_14.mux_l2_in_0_/S
+ mux_bottom_ipin_14.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_276 vgnd vpwr scs8hd_decap_12
XFILLER_18_122 vpwr vgnd scs8hd_fill_2
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_166 vpwr vgnd scs8hd_fill_2
XFILLER_18_199 vpwr vgnd scs8hd_fill_2
XFILLER_24_114 vpwr vgnd scs8hd_fill_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
X_59_ chanx_left_in[14] chanx_right_out[14] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_4.scs8hd_buf_4_0_ mux_bottom_ipin_4.mux_l4_in_0_/X top_grid_pin_20_
+ vgnd vpwr scs8hd_buf_1
XFILLER_24_147 vgnd vpwr scs8hd_decap_6
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_29_239 vgnd vpwr scs8hd_decap_4
XFILLER_29_217 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_6.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_6.mux_l1_in_0_/S mux_bottom_ipin_6.mux_l2_in_3_/S
+ mem_bottom_ipin_6.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_16_36 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_9.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_9.mux_l1_in_2_/S
+ mux_bottom_ipin_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_194 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S mux_bottom_ipin_10.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S mux_bottom_ipin_6.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_264 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__D mux_bottom_ipin_13.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_253 vpwr vgnd scs8hd_fill_2
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XFILLER_16_297 vpwr vgnd scs8hd_fill_2
XFILLER_22_267 vpwr vgnd scs8hd_fill_2
XFILLER_22_289 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_11.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_11.mux_l3_in_0_/S mux_bottom_ipin_11.mux_l4_in_0_/S
+ mem_bottom_ipin_11.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S mux_bottom_ipin_1.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_4
XFILLER_13_267 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1 mux_bottom_ipin_3.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S mux_bottom_ipin_15.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_69 vgnd vpwr scs8hd_decap_4
XFILLER_10_215 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S mux_bottom_ipin_5.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_14.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_14.mux_l1_in_0_/X
+ mux_bottom_ipin_14.mux_l2_in_0_/S mux_bottom_ipin_14.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA__40__A chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_2_288 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S mux_bottom_ipin_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_101 vpwr vgnd scs8hd_fill_2
XFILLER_18_134 vpwr vgnd scs8hd_fill_2
XFILLER_33_148 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_58_ chanx_left_in[15] chanx_right_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_21_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S mux_bottom_ipin_4.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_107 vgnd vpwr scs8hd_decap_4
XANTENNA__35__A chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_30_9 vgnd vpwr scs8hd_decap_3
XFILLER_11_92 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__D mux_bottom_ipin_14.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vgnd vpwr scs8hd_decap_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0 mux_bottom_ipin_14.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_5.mux_l4_in_0_/S mux_bottom_ipin_6.mux_l1_in_0_/S
+ mem_bottom_ipin_6.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XFILLER_32_58 vgnd vpwr scs8hd_decap_12
XFILLER_28_251 vgnd vpwr scs8hd_decap_3
XFILLER_11_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_295 vgnd vpwr scs8hd_decap_4
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S mux_bottom_ipin_5.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S mux_bottom_ipin_3.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0 mux_bottom_ipin_14.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_90 vpwr vgnd scs8hd_fill_2
XFILLER_31_257 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D mux_bottom_ipin_0.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S mux_bottom_ipin_9.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_1.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_1.mux_l3_in_0_/S mux_bottom_ipin_1.mux_l4_in_0_/S
+ mem_bottom_ipin_1.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_bottom_ipin_11.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_11.mux_l2_in_3_/S mux_bottom_ipin_11.mux_l3_in_0_/S
+ mem_bottom_ipin_11.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__43__A chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_2__D mux_top_ipin_0.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_279 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__38__A chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_10.scs8hd_buf_4_0__A mux_bottom_ipin_10.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_3_ _21_/HI chanx_right_in[16] mux_bottom_ipin_0.mux_l2_in_1_/S
+ mux_bottom_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
X_57_ chanx_left_in[16] chanx_right_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_32_171 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_127 vgnd vpwr scs8hd_decap_12
XFILLER_23_171 vpwr vgnd scs8hd_fill_2
XANTENNA__51__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_14.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_14.mux_l1_in_0_/S
+ mux_bottom_ipin_14.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1 mux_bottom_ipin_14.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__D mux_bottom_ipin_2.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_37 vgnd vpwr scs8hd_decap_4
XFILLER_32_15 vgnd vpwr scs8hd_decap_8
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_130 vgnd vpwr scs8hd_decap_4
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_20_163 vpwr vgnd scs8hd_fill_2
XFILLER_28_285 vpwr vgnd scs8hd_fill_2
XFILLER_28_274 vgnd vpwr scs8hd_fill_1
XANTENNA__46__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_22_70 vgnd vpwr scs8hd_decap_3
XFILLER_19_263 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0 mux_bottom_ipin_5.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_26 vpwr vgnd scs8hd_fill_2
XFILLER_25_233 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l4_in_0_ mux_bottom_ipin_0.mux_l3_in_1_/X mux_bottom_ipin_0.mux_l3_in_0_/X
+ mux_bottom_ipin_0.mux_l4_in_0_/S mux_bottom_ipin_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_17_92 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1 mux_bottom_ipin_14.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_1.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_1.mux_l2_in_0_/S mux_bottom_ipin_1.mux_l3_in_0_/S
+ mem_bottom_ipin_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_207 vpwr vgnd scs8hd_fill_2
XFILLER_13_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S mux_bottom_ipin_12.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_11.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_11.mux_l1_in_0_/S mux_bottom_ipin_11.mux_l2_in_3_/S
+ mem_bottom_ipin_11.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0 mux_bottom_ipin_5.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S mux_bottom_ipin_2.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_291 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.scs8hd_buf_4_0__A mux_bottom_ipin_2.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_280 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l2_in_3_ _32_/HI chanx_right_in[15] mux_bottom_ipin_5.mux_l2_in_3_/S
+ mux_bottom_ipin_5.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_206 vpwr vgnd scs8hd_fill_2
XFILLER_10_228 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l3_in_1_ mux_bottom_ipin_0.mux_l2_in_3_/X mux_bottom_ipin_0.mux_l2_in_2_/X
+ mux_bottom_ipin_0.mux_l3_in_0_/S mux_bottom_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_7 vpwr vgnd scs8hd_fill_2
XANTENNA__54__A chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_6
X_73_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1 mux_bottom_ipin_7.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__D mux_bottom_ipin_4.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_147 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S mux_bottom_ipin_11.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__49__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S mux_bottom_ipin_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_106 vgnd vpwr scs8hd_decap_6
XFILLER_26_180 vgnd vpwr scs8hd_decap_4
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_bottom_ipin_0.mux_l2_in_1_/S
+ mux_bottom_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
X_56_ chanx_left_in[17] chanx_right_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_32_150 vgnd vpwr scs8hd_fill_1
XFILLER_24_139 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S mux_bottom_ipin_15.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_21_39 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_5.mux_l4_in_0_ mux_bottom_ipin_5.mux_l3_in_1_/X mux_bottom_ipin_5.mux_l3_in_0_/X
+ mux_bottom_ipin_5.mux_l4_in_0_/S mux_bottom_ipin_5.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_139 vgnd vpwr scs8hd_decap_12
XFILLER_7_19 vpwr vgnd scs8hd_fill_2
XFILLER_11_50 vpwr vgnd scs8hd_fill_2
XFILLER_14_194 vgnd vpwr scs8hd_fill_1
X_39_ chanx_right_in[14] chanx_left_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_186 vpwr vgnd scs8hd_fill_2
XFILLER_28_297 vpwr vgnd scs8hd_fill_2
XFILLER_7_157 vgnd vpwr scs8hd_decap_12
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XANTENNA__62__A chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S mux_bottom_ipin_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1 mux_bottom_ipin_5.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_5.mux_l3_in_1_ mux_bottom_ipin_5.mux_l2_in_3_/X mux_bottom_ipin_5.mux_l2_in_2_/X
+ mux_bottom_ipin_5.mux_l3_in_1_/S mux_bottom_ipin_5.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_25_245 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S mux_bottom_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S mux_bottom_ipin_14.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_9.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_9.mux_l3_in_1_/S mux_bottom_ipin_9.mux_l4_in_0_/S
+ mem_bottom_ipin_9.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__57__A chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1 mux_bottom_ipin_11.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_267 vgnd vpwr scs8hd_decap_6
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_33_81 vgnd vpwr scs8hd_decap_6
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_1.mux_l1_in_1_/S mux_bottom_ipin_1.mux_l2_in_0_/S
+ mem_bottom_ipin_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__D mux_bottom_ipin_5.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_11.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_10.mux_l4_in_0_/S mux_bottom_ipin_11.mux_l1_in_0_/S
+ mem_bottom_ipin_11.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S mux_bottom_ipin_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1 mux_bottom_ipin_5.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_bottom_ipin_5.mux_l2_in_3_/S
+ mux_bottom_ipin_5.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l3_in_0_ mux_bottom_ipin_0.mux_l2_in_1_/X mux_bottom_ipin_0.mux_l2_in_0_/X
+ mux_bottom_ipin_0.mux_l3_in_0_/S mux_bottom_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S mux_bottom_ipin_5.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_83 vpwr vgnd scs8hd_fill_2
XANTENNA__70__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_fill_1
XFILLER_30_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
X_72_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_60 vgnd vpwr scs8hd_fill_1
XANTENNA__65__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_126 vgnd vpwr scs8hd_decap_8
XFILLER_18_148 vgnd vpwr scs8hd_fill_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_107 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_bottom_ipin_0.mux_l1_in_2_/X
+ mux_bottom_ipin_0.mux_l2_in_1_/S mux_bottom_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
X_55_ chanx_left_in[18] chanx_right_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_32_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0 mux_bottom_ipin_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_3
X_38_ chanx_right_in[15] chanx_left_out[15] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__D mux_bottom_ipin_6.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_28_210 vpwr vgnd scs8hd_fill_2
XFILLER_7_169 vgnd vpwr scs8hd_decap_12
XFILLER_7_147 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XFILLER_34_279 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0 mux_bottom_ipin_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l3_in_0_ mux_bottom_ipin_5.mux_l2_in_1_/X mux_bottom_ipin_5.mux_l2_in_0_/X
+ mux_bottom_ipin_5.mux_l3_in_1_/S mux_bottom_ipin_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_13.scs8hd_buf_4_0_ mux_bottom_ipin_13.mux_l4_in_0_/X top_grid_pin_29_
+ vgnd vpwr scs8hd_buf_1
XFILLER_25_268 vpwr vgnd scs8hd_fill_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_9.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_9.mux_l2_in_0_/S mux_bottom_ipin_9.mux_l3_in_1_/S
+ mem_bottom_ipin_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XFILLER_16_235 vgnd vpwr scs8hd_decap_6
XFILLER_16_257 vpwr vgnd scs8hd_fill_2
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__73__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_1.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_0.mux_l4_in_0_/S mux_bottom_ipin_1.mux_l1_in_1_/S
+ mem_bottom_ipin_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_271 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_10.mux_l2_in_3_ _23_/HI chanx_right_in[14] mux_bottom_ipin_10.mux_l2_in_3_/S
+ mux_bottom_ipin_10.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S mux_bottom_ipin_13.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1 mux_bottom_ipin_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_2__S mux_top_ipin_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_21_260 vpwr vgnd scs8hd_fill_2
XANTENNA__68__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l2_in_1_ chanx_left_in[9] mux_bottom_ipin_5.mux_l1_in_2_/X
+ mux_bottom_ipin_5.mux_l2_in_3_/S mux_bottom_ipin_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_260 vgnd vpwr scs8hd_decap_3
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_31 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0 _17_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0 mux_bottom_ipin_9.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
X_71_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_29 vgnd vpwr scs8hd_decap_3
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__D mux_bottom_ipin_8.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_5.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_bottom_ipin_5.mux_l1_in_0_/S
+ mux_bottom_ipin_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S mux_bottom_ipin_12.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_138 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_10.mux_l4_in_0_ mux_bottom_ipin_10.mux_l3_in_1_/X mux_bottom_ipin_10.mux_l3_in_0_/X
+ mux_bottom_ipin_10.mux_l4_in_0_/S mux_bottom_ipin_10.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_0.mux_l2_in_0_ mux_bottom_ipin_0.mux_l1_in_1_/X mux_bottom_ipin_0.mux_l1_in_0_/X
+ mux_bottom_ipin_0.mux_l2_in_1_/S mux_bottom_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
X_54_ chanx_left_in[19] chanx_right_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_32_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1 mux_bottom_ipin_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_108 vpwr vgnd scs8hd_fill_2
XFILLER_23_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
X_37_ chanx_right_in[16] chanx_left_out[16] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_15.mux_l2_in_3_ _28_/HI chanx_right_in[19] mux_bottom_ipin_15.mux_l2_in_3_/S
+ mux_bottom_ipin_15.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_20_111 vpwr vgnd scs8hd_fill_2
XFILLER_20_122 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S mux_bottom_ipin_11.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_155 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_10.mux_l3_in_1_ mux_bottom_ipin_10.mux_l2_in_3_/X mux_bottom_ipin_10.mux_l2_in_2_/X
+ mux_bottom_ipin_10.mux_l3_in_1_/S mux_bottom_ipin_10.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_40 vgnd vpwr scs8hd_decap_4
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0 _24_/HI vgnd vpwr scs8hd_diode_2
XFILLER_19_255 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1 mux_bottom_ipin_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0 mux_bottom_ipin_13.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_203 vpwr vgnd scs8hd_fill_2
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_9.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_9.mux_l1_in_2_/S mux_bottom_ipin_9.mux_l2_in_0_/S
+ mem_bottom_ipin_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_40 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_94 vgnd vpwr scs8hd_decap_12
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1 mux_bottom_ipin_9.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__D mux_bottom_ipin_11.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_10.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_bottom_ipin_10.mux_l2_in_3_/S
+ mux_bottom_ipin_10.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S mux_bottom_ipin_12.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_217 vpwr vgnd scs8hd_fill_2
XFILLER_21_250 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S mux_bottom_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S mux_bottom_ipin_10.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_61 vpwr vgnd scs8hd_fill_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_15.mux_l4_in_0_ mux_bottom_ipin_15.mux_l3_in_1_/X mux_bottom_ipin_15.mux_l3_in_0_/X
+ mux_bottom_ipin_15.mux_l4_in_0_/S mux_bottom_ipin_15.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l2_in_0_ mux_bottom_ipin_5.mux_l1_in_1_/X mux_bottom_ipin_5.mux_l1_in_0_/X
+ mux_bottom_ipin_5.mux_l2_in_3_/S mux_bottom_ipin_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_298 vgnd vpwr scs8hd_fill_1
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S mux_bottom_ipin_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1 mux_bottom_ipin_9.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_41 vpwr vgnd scs8hd_fill_2
XFILLER_5_279 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_14.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_14.mux_l3_in_0_/S mux_bottom_ipin_14.mux_l4_in_0_/S
+ mem_bottom_ipin_14.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
X_70_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_15.mux_l3_in_1_ mux_bottom_ipin_15.mux_l2_in_3_/X mux_bottom_ipin_15.mux_l2_in_2_/X
+ mux_bottom_ipin_15.mux_l3_in_0_/S mux_bottom_ipin_15.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_5.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_5.mux_l1_in_0_/S
+ mux_bottom_ipin_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_150 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XFILLER_25_62 vgnd vpwr scs8hd_decap_4
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S mux_bottom_ipin_1.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_53_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_142 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S mux_bottom_ipin_7.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1 mux_bottom_ipin_13.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_20 vpwr vgnd scs8hd_fill_2
XFILLER_11_42 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
XFILLER_14_164 vpwr vgnd scs8hd_fill_2
XFILLER_14_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
X_36_ chanx_right_in[17] chanx_left_out[17] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_15.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_bottom_ipin_15.mux_l2_in_3_/S
+ mux_bottom_ipin_15.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__D mux_bottom_ipin_13.mux_l1_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_190 vpwr vgnd scs8hd_fill_2
XFILLER_20_145 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_28_289 vgnd vpwr scs8hd_decap_8
XFILLER_28_267 vgnd vpwr scs8hd_decap_4
XFILLER_28_256 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_10.mux_l3_in_0_ mux_bottom_ipin_10.mux_l2_in_1_/X mux_bottom_ipin_10.mux_l2_in_0_/X
+ mux_bottom_ipin_10.mux_l3_in_1_/S mux_bottom_ipin_10.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_19_212 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_fill_1
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_65 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
X_19_ _19_/HI _19_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1 mux_bottom_ipin_13.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_237 vpwr vgnd scs8hd_fill_2
XFILLER_25_215 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_9.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_8.mux_l4_in_0_/S mux_bottom_ipin_9.mux_l1_in_2_/S
+ mem_bottom_ipin_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0 _29_/HI vgnd vpwr scs8hd_diode_2
XFILLER_24_270 vpwr vgnd scs8hd_fill_2
XFILLER_17_30 vpwr vgnd scs8hd_fill_2
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_292 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0 mux_bottom_ipin_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_10.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_bottom_ipin_10.mux_l2_in_3_/S
+ mux_bottom_ipin_10.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_229 vgnd vpwr scs8hd_decap_12
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XFILLER_21_295 vgnd vpwr scs8hd_decap_4
XFILLER_28_84 vgnd vpwr scs8hd_decap_6
XFILLER_28_73 vpwr vgnd scs8hd_fill_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_8_200 vpwr vgnd scs8hd_fill_2
XFILLER_5_55 vgnd vpwr scs8hd_decap_6
XFILLER_12_284 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_4.mux_l3_in_1_/S mux_bottom_ipin_4.mux_l4_in_0_/S
+ mem_bottom_ipin_4.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_6
XFILLER_14_64 vpwr vgnd scs8hd_fill_2
XFILLER_14_75 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_14.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_14.mux_l2_in_0_/S mux_bottom_ipin_14.mux_l3_in_0_/S
+ mem_bottom_ipin_14.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_ipin_5.scs8hd_buf_4_0_ mux_bottom_ipin_5.mux_l4_in_0_/X top_grid_pin_21_
+ vgnd vpwr scs8hd_buf_1
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_15.mux_l3_in_0_ mux_bottom_ipin_15.mux_l2_in_1_/X mux_bottom_ipin_15.mux_l2_in_0_/X
+ mux_bottom_ipin_15.mux_l3_in_0_/S mux_bottom_ipin_15.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__D mux_bottom_ipin_14.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l2_in_0__S mux_top_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_5.mux_l1_in_0_/S
+ mux_bottom_ipin_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XFILLER_25_52 vpwr vgnd scs8hd_fill_2
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
X_52_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_1_283 vgnd vpwr scs8hd_decap_12
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XFILLER_23_198 vpwr vgnd scs8hd_fill_2
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XFILLER_11_54 vgnd vpwr scs8hd_decap_4
XFILLER_14_154 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_13.scs8hd_buf_4_0__A mux_bottom_ipin_13.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
X_35_ chanx_right_in[18] chanx_left_out[18] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_15.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_bottom_ipin_15.mux_l2_in_3_/S
+ mux_bottom_ipin_15.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1 mux_bottom_ipin_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_224 vpwr vgnd scs8hd_fill_2
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__D mux_bottom_ipin_0.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_97 vpwr vgnd scs8hd_fill_2
XFILLER_19_235 vpwr vgnd scs8hd_fill_2
XFILLER_19_268 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XFILLER_8_11 vpwr vgnd scs8hd_fill_2
XFILLER_8_77 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_18_ _18_/HI _18_/LO vgnd vpwr scs8hd_conb_1
XFILLER_33_282 vgnd vpwr scs8hd_decap_12
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_219 vgnd vpwr scs8hd_decap_12
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_12_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_30_285 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1 mux_bottom_ipin_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_219 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_10.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_10.mux_l1_in_0_/X
+ mux_bottom_ipin_10.mux_l2_in_3_/S mux_bottom_ipin_10.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__D mux_bottom_ipin_15.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S mux_bottom_ipin_13.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__S mux_top_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_41 vgnd vpwr scs8hd_fill_1
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XFILLER_8_212 vpwr vgnd scs8hd_fill_2
XFILLER_12_296 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S mux_bottom_ipin_9.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_4.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_4.mux_l2_in_2_/S mux_bottom_ipin_4.mux_l3_in_1_/S
+ mem_bottom_ipin_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_30_86 vgnd vpwr scs8hd_decap_4
XFILLER_30_75 vgnd vpwr scs8hd_decap_4
XFILLER_30_64 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_14.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_14.mux_l1_in_0_/S mux_bottom_ipin_14.mux_l2_in_0_/S
+ mem_bottom_ipin_14.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.scs8hd_buf_4_0__A mux_bottom_ipin_5.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S mux_bottom_ipin_12.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S mux_bottom_ipin_4.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_163 vpwr vgnd scs8hd_fill_2
XFILLER_25_20 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__D mux_bottom_ipin_1.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
X_51_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_1_295 vgnd vpwr scs8hd_decap_4
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_188 vpwr vgnd scs8hd_fill_2
XFILLER_32_166 vgnd vpwr scs8hd_decap_3
XFILLER_17_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0 mux_bottom_ipin_15.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S mux_bottom_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_15.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_15.mux_l1_in_0_/X
+ mux_bottom_ipin_15.mux_l2_in_3_/S mux_bottom_ipin_15.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
X_34_ chanx_right_in[19] chanx_left_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_20_158 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S mux_bottom_ipin_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_147 vgnd vpwr scs8hd_decap_8
XFILLER_11_158 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0 mux_bottom_ipin_15.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_27_291 vpwr vgnd scs8hd_fill_2
XFILLER_8_56 vgnd vpwr scs8hd_fill_1
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
X_17_ _17_/HI _17_/LO vgnd vpwr scs8hd_conb_1
XFILLER_33_294 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S mux_bottom_ipin_7.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XFILLER_16_228 vgnd vpwr scs8hd_decap_4
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_30_297 vpwr vgnd scs8hd_fill_2
XFILLER_15_272 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_0.mux_l2_in_3_ _20_/HI chanx_right_in[16] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_264 vpwr vgnd scs8hd_fill_2
XFILLER_28_20 vgnd vpwr scs8hd_decap_4
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.scs8hd_buf_4_0_ mux_bottom_ipin_0.mux_l4_in_0_/X top_grid_pin_16_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__D mux_bottom_ipin_3.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0 mux_bottom_ipin_8.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S mux_bottom_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_4.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_4.mux_l1_in_1_/S mux_bottom_ipin_4.mux_l2_in_2_/S
+ mem_bottom_ipin_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_290 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S mux_bottom_ipin_6.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_4
XFILLER_29_161 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_14.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_13.mux_l4_in_0_/S mux_bottom_ipin_14.mux_l1_in_0_/S
+ mem_bottom_ipin_14.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_ipin_10.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_10.mux_l1_in_0_/S
+ mux_bottom_ipin_10.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_197 vgnd vpwr scs8hd_decap_8
XFILLER_26_186 vpwr vgnd scs8hd_fill_2
XFILLER_26_131 vgnd vpwr scs8hd_decap_4
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_43 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ ccff_tail mux_top_ipin_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_50_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1 mux_bottom_ipin_15.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_101 vpwr vgnd scs8hd_fill_2
XFILLER_14_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0 mux_bottom_ipin_6.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
X_33_ _33_/HI _33_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_126 vpwr vgnd scs8hd_fill_2
XFILLER_11_104 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_0_/S mux_top_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_22 vgnd vpwr scs8hd_decap_4
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0 mux_bottom_ipin_12.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1 mux_bottom_ipin_15.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__D mux_bottom_ipin_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.mux_l2_in_3_ _22_/HI chanx_right_in[17] mux_bottom_ipin_1.mux_l2_in_0_/S
+ mux_bottom_ipin_1.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XFILLER_25_229 vpwr vgnd scs8hd_fill_2
XFILLER_25_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_88 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_65 vpwr vgnd scs8hd_fill_2
XFILLER_33_21 vgnd vpwr scs8hd_decap_12
XFILLER_33_10 vgnd vpwr scs8hd_decap_4
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0 mux_bottom_ipin_6.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_15.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_15.mux_l1_in_0_/S
+ mux_bottom_ipin_15.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_15_284 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_ipin_0.mux_l3_in_1__A0 mux_top_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_287 vpwr vgnd scs8hd_fill_2
XFILLER_28_65 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_12_210 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1 mux_bottom_ipin_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_4.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_3.mux_l4_in_0_/S mux_bottom_ipin_4.mux_l1_in_1_/S
+ mem_bottom_ipin_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_ipin_1.mux_l4_in_0_ mux_bottom_ipin_1.mux_l3_in_1_/X mux_bottom_ipin_1.mux_l3_in_0_/X
+ mux_bottom_ipin_1.mux_l4_in_0_/S mux_bottom_ipin_1.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0 mux_bottom_ipin_10.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_173 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l4_in_0__A0 mux_top_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l3_in_1__S mux_top_ipin_0.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S mux_bottom_ipin_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_25_66 vgnd vpwr scs8hd_fill_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_6.mux_l2_in_3_ _33_/HI chanx_right_in[18] mux_bottom_ipin_6.mux_l2_in_3_/S
+ mux_bottom_ipin_6.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__D mux_bottom_ipin_6.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l3_in_1_ mux_bottom_ipin_1.mux_l2_in_3_/X mux_bottom_ipin_1.mux_l2_in_2_/X
+ mux_bottom_ipin_1.mux_l3_in_0_/S mux_bottom_ipin_1.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0 mux_bottom_ipin_10.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_24 vgnd vpwr scs8hd_decap_3
XFILLER_14_168 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S mux_bottom_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1 mux_bottom_ipin_6.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
X_32_ _32_/HI _32_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_194 vpwr vgnd scs8hd_fill_2
XFILLER_13_190 vpwr vgnd scs8hd_fill_2
XFILLER_20_149 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_0_/S mux_top_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S mux_bottom_ipin_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_116 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S mux_bottom_ipin_4.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1 mux_bottom_ipin_12.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_36 vgnd vpwr scs8hd_decap_12
XFILLER_10_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_bottom_ipin_1.mux_l2_in_0_/S
+ mux_bottom_ipin_1.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_219 vgnd vpwr scs8hd_fill_1
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_6.mux_l4_in_0_ mux_bottom_ipin_6.mux_l3_in_1_/X mux_bottom_ipin_6.mux_l3_in_0_/X
+ mux_bottom_ipin_6.mux_l4_in_0_/S mux_bottom_ipin_6.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1 mux_bottom_ipin_6.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_230 vgnd vpwr scs8hd_decap_8
XFILLER_17_34 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_33 vgnd vpwr scs8hd_decap_3
XFILLER_24_285 vpwr vgnd scs8hd_fill_2
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_30_255 vgnd vpwr scs8hd_fill_1
XFILLER_30_211 vgnd vpwr scs8hd_decap_3
XFILLER_15_230 vpwr vgnd scs8hd_fill_2
XFILLER_15_296 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_ipin_0.mux_l3_in_1__A1 mux_top_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S mux_bottom_ipin_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__D mux_bottom_ipin_9.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__D mux_bottom_ipin_7.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l3_in_1_ mux_bottom_ipin_6.mux_l2_in_3_/X mux_bottom_ipin_6.mux_l2_in_2_/X
+ mux_bottom_ipin_6.mux_l3_in_1_/S mux_bottom_ipin_6.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S mux_bottom_ipin_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_23 vgnd vpwr scs8hd_fill_1
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1 mux_bottom_ipin_10.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_0.mux_l1_in_0_/S
+ mux_top_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_ipin_0.mux_l4_in_0__A1 mux_top_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0 mux_bottom_ipin_1.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XFILLER_26_144 vgnd vpwr scs8hd_decap_6
XFILLER_26_111 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_56 vgnd vpwr scs8hd_decap_4
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S mux_bottom_ipin_4.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S mux_bottom_ipin_2.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_bottom_ipin_6.mux_l2_in_3_/S
+ mux_bottom_ipin_6.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_155 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l3_in_0_ mux_bottom_ipin_1.mux_l2_in_1_/X mux_bottom_ipin_1.mux_l2_in_0_/X
+ mux_bottom_ipin_1.mux_l3_in_0_/S mux_bottom_ipin_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1 mux_bottom_ipin_10.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S mux_bottom_ipin_8.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_11_58 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A mux_bottom_ipin_0.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_191 vpwr vgnd scs8hd_fill_2
X_31_ _31_/HI _31_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0 mux_bottom_ipin_1.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_14.scs8hd_buf_4_0_ mux_bottom_ipin_14.mux_l4_in_0_/X top_grid_pin_30_
+ vgnd vpwr scs8hd_buf_1
XFILLER_28_228 vgnd vpwr scs8hd_decap_4
XFILLER_28_206 vpwr vgnd scs8hd_fill_2
XFILLER_22_46 vgnd vpwr scs8hd_fill_1
XFILLER_19_239 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__D mux_bottom_ipin_10.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_59 vgnd vpwr scs8hd_decap_4
XFILLER_8_48 vgnd vpwr scs8hd_decap_8
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.mux_l2_in_1_ chanx_left_in[11] mux_bottom_ipin_1.mux_l1_in_2_/X
+ mux_bottom_ipin_1.mux_l2_in_0_/S mux_bottom_ipin_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__D mux_bottom_ipin_9.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_261 vpwr vgnd scs8hd_fill_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1 mux_bottom_ipin_3.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_253 vpwr vgnd scs8hd_fill_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_24_297 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_30_289 vgnd vpwr scs8hd_decap_8
XFILLER_30_267 vpwr vgnd scs8hd_fill_2
XFILLER_15_264 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0 _18_/HI vgnd vpwr scs8hd_diode_2
XFILLER_21_245 vgnd vpwr scs8hd_decap_3
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_1.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_bottom_ipin_1.mux_l1_in_1_/S
+ mux_bottom_ipin_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_12_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l3_in_0_ mux_bottom_ipin_6.mux_l2_in_1_/X mux_bottom_ipin_6.mux_l2_in_0_/X
+ mux_bottom_ipin_6.mux_l3_in_1_/S mux_bottom_ipin_6.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_58 vgnd vpwr scs8hd_decap_4
XFILLER_30_79 vgnd vpwr scs8hd_fill_1
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_29_197 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_0.mux_l1_in_0_/S
+ mux_top_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_296 vgnd vpwr scs8hd_decap_3
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_11.mux_l2_in_3_ _24_/HI chanx_right_in[15] mux_bottom_ipin_11.mux_l2_in_3_/S
+ mux_bottom_ipin_11.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1 mux_bottom_ipin_1.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_167 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_7.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_7.mux_l3_in_0_/S mux_bottom_ipin_7.mux_l4_in_0_/S
+ mem_bottom_ipin_7.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_57 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_6.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_bottom_ipin_6.mux_l2_in_3_/S
+ mux_bottom_ipin_6.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__D mux_bottom_ipin_12.mux_l2_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_31_192 vpwr vgnd scs8hd_fill_2
XFILLER_23_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S mux_bottom_ipin_1.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0 _25_/HI vgnd vpwr scs8hd_diode_2
X_30_ _30_/HI _30_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1 mux_bottom_ipin_1.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0 mux_bottom_ipin_14.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S mux_bottom_ipin_15.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_36 vpwr vgnd scs8hd_fill_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_207 vgnd vpwr scs8hd_decap_3
XFILLER_27_295 vgnd vpwr scs8hd_decap_4
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_11.mux_l4_in_0_ mux_bottom_ipin_11.mux_l3_in_1_/X mux_bottom_ipin_11.mux_l3_in_0_/X
+ mux_bottom_ipin_11.mux_l4_in_0_/S mux_bottom_ipin_11.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_162 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_1.mux_l2_in_0_ mux_bottom_ipin_1.mux_l1_in_1_/X mux_bottom_ipin_1.mux_l1_in_0_/X
+ mux_bottom_ipin_1.mux_l2_in_0_/S mux_bottom_ipin_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_254 vpwr vgnd scs8hd_fill_2
XFILLER_33_210 vpwr vgnd scs8hd_fill_2
XFILLER_33_298 vgnd vpwr scs8hd_fill_1
XFILLER_33_265 vpwr vgnd scs8hd_fill_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S mux_bottom_ipin_10.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S mux_bottom_ipin_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_235 vgnd vpwr scs8hd_decap_12
XFILLER_30_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_24_3 vgnd vpwr scs8hd_fill_1
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_21_213 vpwr vgnd scs8hd_fill_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_11.mux_l3_in_1_ mux_bottom_ipin_11.mux_l2_in_3_/X mux_bottom_ipin_11.mux_l2_in_2_/X
+ mux_bottom_ipin_11.mux_l3_in_0_/S mux_bottom_ipin_11.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S mux_bottom_ipin_14.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_1.mux_l1_in_1_/S
+ mux_bottom_ipin_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_12_224 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__D mux_bottom_ipin_14.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_58 vgnd vpwr scs8hd_decap_4
XFILLER_30_36 vgnd vpwr scs8hd_fill_1
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_0.mux_l1_in_0_/S
+ mux_top_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_11.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_bottom_ipin_11.mux_l2_in_3_/S
+ mux_bottom_ipin_11.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S mux_bottom_ipin_15.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S mux_bottom_ipin_13.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_135 vgnd vpwr scs8hd_fill_1
XFILLER_26_102 vgnd vpwr scs8hd_decap_3
XFILLER_25_69 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S mux_bottom_ipin_5.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_36 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_7.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_7.mux_l2_in_3_/S mux_bottom_ipin_7.mux_l3_in_0_/S
+ mem_bottom_ipin_7.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_6.mux_l1_in_0_/X
+ mux_bottom_ipin_6.mux_l2_in_3_/S mux_bottom_ipin_6.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D mux_bottom_ipin_0.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_8.scs8hd_buf_4_0__A mux_bottom_ipin_8.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_160 vgnd vpwr scs8hd_decap_6
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XFILLER_11_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XANTENNA__41__A chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_0__D mux_bottom_ipin_15.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_171 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S mux_bottom_ipin_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1 mux_bottom_ipin_14.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S mux_bottom_ipin_4.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0 _30_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__36__A chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_12_81 vgnd vpwr scs8hd_decap_8
XFILLER_18_230 vgnd vpwr scs8hd_decap_4
XFILLER_18_241 vgnd vpwr scs8hd_fill_1
XFILLER_18_274 vgnd vpwr scs8hd_fill_1
XFILLER_18_285 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0 mux_bottom_ipin_5.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_69 vgnd vpwr scs8hd_decap_12
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_266 vpwr vgnd scs8hd_fill_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_30_203 vpwr vgnd scs8hd_fill_2
XFILLER_15_222 vpwr vgnd scs8hd_fill_2
XFILLER_30_247 vgnd vpwr scs8hd_decap_8
XFILLER_15_288 vpwr vgnd scs8hd_fill_2
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_203 vpwr vgnd scs8hd_fill_2
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_36 vgnd vpwr scs8hd_decap_3
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_11.mux_l3_in_0_ mux_bottom_ipin_11.mux_l2_in_1_/X mux_bottom_ipin_11.mux_l2_in_0_/X
+ mux_bottom_ipin_11.mux_l3_in_0_/S mux_bottom_ipin_11.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_28_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_1.mux_l1_in_1_/S
+ mux_bottom_ipin_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_236 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_291 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.scs8hd_buf_4_0_ mux_bottom_ipin_6.mux_l4_in_0_/X top_grid_pin_22_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__D mux_bottom_ipin_1.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_30_26 vgnd vpwr scs8hd_decap_3
XFILLER_30_15 vpwr vgnd scs8hd_fill_2
XANTENNA__44__A chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_3__D mux_top_ipin_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_276 vgnd vpwr scs8hd_decap_12
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_11.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_bottom_ipin_11.mux_l2_in_3_/S
+ mux_bottom_ipin_11.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_59 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_7.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_7.mux_l1_in_0_/S mux_bottom_ipin_7.mux_l2_in_3_/S
+ mem_bottom_ipin_7.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_25_48 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__39__A chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_279 vpwr vgnd scs8hd_fill_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_147 vgnd vpwr scs8hd_decap_6
XFILLER_31_91 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1 mux_bottom_ipin_5.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S mux_bottom_ipin_12.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_183 vpwr vgnd scs8hd_fill_2
XFILLER_13_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_6.mux_l1_in_0_/S
+ mux_bottom_ipin_6.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_27_264 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_12.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_12.mux_l3_in_1_/S mux_bottom_ipin_12.mux_l4_in_0_/S
+ mem_bottom_ipin_12.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__52__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XFILLER_18_220 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1 mux_bottom_ipin_5.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_278 vpwr vgnd scs8hd_fill_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_6
XFILLER_18_297 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__D mux_bottom_ipin_2.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_289 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S mux_bottom_ipin_11.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__47__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_15_234 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_3
XFILLER_0_85 vgnd vpwr scs8hd_decap_8
XFILLER_9_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_28_26 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_19 vgnd vpwr scs8hd_decap_12
XFILLER_12_248 vgnd vpwr scs8hd_decap_12
XFILLER_20_270 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S mux_bottom_ipin_10.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA__60__A chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_4_288 vgnd vpwr scs8hd_decap_8
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_11.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_11.mux_l1_in_0_/X
+ mux_bottom_ipin_11.mux_l2_in_3_/S mux_bottom_ipin_11.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_ipin_7.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_6.mux_l4_in_0_/S mux_bottom_ipin_7.mux_l1_in_0_/S
+ mem_bottom_ipin_7.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_1_269 vgnd vpwr scs8hd_decap_6
XFILLER_32_107 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_0.scs8hd_dfxbp_1_3_ prog_clk mux_top_ipin_0.mux_l3_in_0_/S ccff_tail
+ mem_top_ipin_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__55__A chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_17_159 vpwr vgnd scs8hd_fill_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_0_280 vgnd vpwr scs8hd_decap_12
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_3
XFILLER_31_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__D mux_bottom_ipin_4.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0 mux_bottom_ipin_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_22_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S mux_bottom_ipin_11.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S mux_bottom_ipin_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_100 vgnd vpwr scs8hd_decap_12
XFILLER_13_162 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_4
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_2.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_2.mux_l3_in_0_/S mux_bottom_ipin_2.mux_l4_in_0_/S
+ mem_bottom_ipin_2.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S mux_bottom_ipin_15.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_ipin_12.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_12.mux_l2_in_2_/S mux_bottom_ipin_12.mux_l3_in_1_/S
+ mem_bottom_ipin_12.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_19 vpwr vgnd scs8hd_fill_2
XFILLER_10_154 vgnd vpwr scs8hd_decap_8
XFILLER_10_165 vpwr vgnd scs8hd_fill_2
XFILLER_33_202 vgnd vpwr scs8hd_decap_4
XFILLER_18_265 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_38 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.scs8hd_buf_4_0_ mux_bottom_ipin_1.mux_l4_in_0_/X top_grid_pin_17_
+ vgnd vpwr scs8hd_buf_1
XANTENNA__63__A chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S mux_bottom_ipin_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_268 vgnd vpwr scs8hd_decap_4
XFILLER_23_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0 mux_bottom_ipin_9.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_62 vgnd vpwr scs8hd_fill_1
XFILLER_28_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S mux_bottom_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__58__A chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_18_82 vgnd vpwr scs8hd_fill_1
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XFILLER_11_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_11.scs8hd_buf_4_0__A mux_bottom_ipin_11.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_275 vgnd vpwr scs8hd_fill_1
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__D mux_bottom_ipin_6.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1 mux_bottom_ipin_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_61 vgnd vpwr scs8hd_fill_1
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_26_138 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_9_7 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.scs8hd_dfxbp_1_2_ prog_clk mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l3_in_0_/S
+ mem_top_ipin_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__71__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0 mux_bottom_ipin_7.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_292 vgnd vpwr scs8hd_decap_6
XFILLER_16_193 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S mux_bottom_ipin_9.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1 mux_bottom_ipin_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__S mux_top_ipin_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_22_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0 mux_bottom_ipin_13.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__66__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_11.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_11.mux_l1_in_0_/S
+ mux_bottom_ipin_11.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_71 vpwr vgnd scs8hd_fill_2
XFILLER_9_112 vgnd vpwr scs8hd_decap_8
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_2.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_2.mux_l2_in_0_/S mux_bottom_ipin_2.mux_l3_in_0_/S
+ mem_bottom_ipin_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0 mux_bottom_ipin_7.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_200 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_12.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_12.mux_l1_in_2_/S mux_bottom_ipin_12.mux_l2_in_2_/S
+ mem_bottom_ipin_12.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_62 vgnd vpwr scs8hd_fill_1
XFILLER_33_214 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_3.scs8hd_buf_4_0__A mux_bottom_ipin_3.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_18_211 vgnd vpwr scs8hd_fill_1
XFILLER_33_269 vgnd vpwr scs8hd_decap_6
XFILLER_33_258 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_17 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_69_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__D mux_bottom_ipin_7.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1 mux_bottom_ipin_9.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0 mux_bottom_ipin_11.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_261 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l2_in_3_ _29_/HI chanx_right_in[14] mux_bottom_ipin_2.mux_l2_in_0_/S
+ mux_bottom_ipin_2.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_61 vpwr vgnd scs8hd_fill_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XFILLER_11_283 vpwr vgnd scs8hd_fill_2
XFILLER_7_298 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_29_136 vgnd vpwr scs8hd_decap_4
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S mux_bottom_ipin_13.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XANTENNA__69__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_29_93 vgnd vpwr scs8hd_fill_1
XFILLER_29_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0 mux_bottom_ipin_11.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_17_106 vpwr vgnd scs8hd_fill_2
XFILLER_25_161 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.scs8hd_dfxbp_1_1_ prog_clk mux_top_ipin_0.mux_l1_in_0_/S mux_top_ipin_0.mux_l2_in_2_/S
+ mem_top_ipin_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_83 vgnd vpwr scs8hd_fill_1
XFILLER_15_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1 mux_bottom_ipin_7.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_109 vgnd vpwr scs8hd_decap_3
XFILLER_16_172 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l4_in_0_ mux_bottom_ipin_2.mux_l3_in_1_/X mux_bottom_ipin_2.mux_l3_in_0_/X
+ mux_bottom_ipin_2.mux_l4_in_0_/S mux_bottom_ipin_2.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__D mux_bottom_ipin_10.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__D mux_bottom_ipin_8.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S mux_bottom_ipin_12.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1 mux_bottom_ipin_13.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_2.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_2.mux_l1_in_0_/S mux_bottom_ipin_2.mux_l2_in_0_/S
+ mem_bottom_ipin_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S mux_bottom_ipin_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1 mux_bottom_ipin_7.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_3_ _17_/HI chanx_right_in[19] mux_bottom_ipin_7.mux_l2_in_3_/S
+ mux_bottom_ipin_7.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0 mux_bottom_ipin_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_12.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_11.mux_l4_in_0_/S mux_bottom_ipin_12.mux_l1_in_2_/S
+ mem_bottom_ipin_12.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_189 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_33_226 vgnd vpwr scs8hd_decap_12
XFILLER_18_234 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l3_in_1_ mux_bottom_ipin_2.mux_l2_in_3_/X mux_bottom_ipin_2.mux_l2_in_2_/X
+ mux_bottom_ipin_2.mux_l3_in_0_/S mux_bottom_ipin_2.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
X_68_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_24_226 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S mux_bottom_ipin_11.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_30_207 vpwr vgnd scs8hd_fill_2
XFILLER_23_292 vpwr vgnd scs8hd_fill_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
XFILLER_21_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S mux_bottom_ipin_7.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1 mux_bottom_ipin_11.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_40 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_2.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_bottom_ipin_2.mux_l2_in_0_/S
+ mux_bottom_ipin_2.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_295 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_7.mux_l4_in_0_ mux_bottom_ipin_7.mux_l3_in_1_/X mux_bottom_ipin_7.mux_l3_in_0_/X
+ mux_bottom_ipin_7.mux_l4_in_0_/S mux_bottom_ipin_7.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_19 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0 mux_bottom_ipin_2.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__D mux_bottom_ipin_11.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S mux_bottom_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_41 vgnd vpwr scs8hd_decap_3
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_29_50 vpwr vgnd scs8hd_fill_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1 mux_bottom_ipin_11.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_151 vpwr vgnd scs8hd_fill_2
XFILLER_26_107 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_34_195 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S mux_bottom_ipin_6.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_118 vgnd vpwr scs8hd_decap_4
XFILLER_25_173 vpwr vgnd scs8hd_fill_2
XFILLER_15_30 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_15.mux_l4_in_0_/S mux_top_ipin_0.mux_l1_in_0_/S
+ mem_top_ipin_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_51 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l3_in_1_ mux_bottom_ipin_7.mux_l2_in_3_/X mux_bottom_ipin_7.mux_l2_in_2_/X
+ mux_bottom_ipin_7.mux_l3_in_0_/S mux_bottom_ipin_7.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0 mux_bottom_ipin_2.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_143 vgnd vpwr scs8hd_decap_6
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_15.scs8hd_buf_4_0_ mux_bottom_ipin_15.mux_l4_in_0_/X top_grid_pin_31_
+ vgnd vpwr scs8hd_buf_1
XFILLER_22_187 vpwr vgnd scs8hd_fill_2
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_2.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_ipin_1.mux_l4_in_0_/S mux_bottom_ipin_2.mux_l1_in_0_/S
+ mem_bottom_ipin_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S mux_bottom_ipin_7.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1 mux_bottom_ipin_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_bottom_ipin_7.mux_l2_in_3_/S
+ mux_bottom_ipin_7.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_268 vpwr vgnd scs8hd_fill_2
XFILLER_27_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S mux_bottom_ipin_5.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XFILLER_12_75 vgnd vpwr scs8hd_decap_4
XFILLER_33_238 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_2.mux_l3_in_0_ mux_bottom_ipin_2.mux_l2_in_1_/X mux_bottom_ipin_2.mux_l2_in_0_/X
+ mux_bottom_ipin_2.mux_l3_in_0_/S mux_bottom_ipin_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0 _19_/HI vgnd vpwr scs8hd_diode_2
XFILLER_24_205 vpwr vgnd scs8hd_fill_2
X_67_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_24_249 vpwr vgnd scs8hd_fill_2
XFILLER_24_238 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__D mux_bottom_ipin_13.mux_l2_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_23_271 vgnd vpwr scs8hd_decap_4
XFILLER_9_76 vgnd vpwr scs8hd_decap_12
XFILLER_9_43 vpwr vgnd scs8hd_fill_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_20_285 vpwr vgnd scs8hd_fill_2
XFILLER_18_74 vpwr vgnd scs8hd_fill_2
XFILLER_18_85 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_bottom_ipin_2.mux_l2_in_0_/S
+ mux_bottom_ipin_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_40 vpwr vgnd scs8hd_fill_2
XFILLER_7_278 vgnd vpwr scs8hd_decap_12
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1 mux_bottom_ipin_2.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_20_53 vpwr vgnd scs8hd_fill_2
XFILLER_20_64 vgnd vpwr scs8hd_fill_1
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_11 vgnd vpwr scs8hd_decap_4
XFILLER_3_281 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vgnd vpwr scs8hd_fill_1
XFILLER_34_174 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_7.mux_l3_in_0_ mux_bottom_ipin_7.mux_l2_in_1_/X mux_bottom_ipin_7.mux_l2_in_0_/X
+ mux_bottom_ipin_7.mux_l3_in_0_/S mux_bottom_ipin_7.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XFILLER_31_96 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0 _26_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1 mux_bottom_ipin_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_273 vgnd vpwr scs8hd_decap_6
XFILLER_31_177 vgnd vpwr scs8hd_decap_4
XFILLER_31_166 vgnd vpwr scs8hd_fill_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0 mux_bottom_ipin_15.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
.ends

