VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_bottom
  CLASS BLOCK ;
  FOREIGN grid_io_bottom ;
  ORIGIN 0.000 0.000 ;
  SIZE 144.630 BY 120.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 2.400 99.920 ;
    END
  END ccff_tail
  PIN gfpga_pad_GPIO_A
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END gfpga_pad_GPIO_A
  PIN gfpga_pad_GPIO_IE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END gfpga_pad_GPIO_IE
  PIN gfpga_pad_GPIO_OE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 2.400 ;
    END
  END gfpga_pad_GPIO_OE
  PIN gfpga_pad_GPIO_Y
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 2.400 ;
    END
  END gfpga_pad_GPIO_Y
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END prog_clk
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 117.600 74.890 120.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 117.600 125.030 120.000 ;
    END
  END top_width_0_height_0__pin_1_lower
  PIN top_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 117.600 25.210 120.000 ;
    END
  END top_width_0_height_0__pin_1_upper
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.720 10.640 31.320 109.040 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 54.720 10.640 56.320 109.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 108.885 ;
      LAYER met1 ;
        RECT 5.520 9.900 144.440 109.040 ;
      LAYER met2 ;
        RECT 7.450 117.320 24.650 117.600 ;
        RECT 25.490 117.320 74.330 117.600 ;
        RECT 75.170 117.320 124.470 117.600 ;
        RECT 125.310 117.320 131.260 117.600 ;
        RECT 7.450 2.680 131.260 117.320 ;
        RECT 7.450 2.400 18.210 2.680 ;
        RECT 19.050 2.400 55.470 2.680 ;
        RECT 56.310 2.400 93.190 2.680 ;
        RECT 94.030 2.400 130.450 2.680 ;
      LAYER met3 ;
        RECT 2.400 100.320 131.320 108.965 ;
        RECT 2.800 98.920 131.320 100.320 ;
        RECT 2.400 60.200 131.320 98.920 ;
        RECT 2.800 58.800 131.320 60.200 ;
        RECT 2.400 20.760 131.320 58.800 ;
        RECT 2.800 19.360 131.320 20.760 ;
        RECT 2.400 6.975 131.320 19.360 ;
      LAYER met4 ;
        RECT 79.720 10.640 131.320 109.040 ;
  END
END grid_io_bottom
END LIBRARY

