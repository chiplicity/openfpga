magic
tech sky130A
magscale 1 2
timestamp 1606475469
<< locali >>
rect 14381 11679 14415 11849
rect 15945 11747 15979 11849
rect 12265 10523 12299 10693
rect 2053 7735 2087 7905
rect 8401 7259 8435 7497
<< viali >>
rect 1961 20009 1995 20043
rect 4537 20009 4571 20043
rect 5273 20009 5307 20043
rect 5733 20009 5767 20043
rect 9137 20009 9171 20043
rect 13001 20009 13035 20043
rect 14289 20009 14323 20043
rect 14841 20009 14875 20043
rect 15669 20009 15703 20043
rect 16221 20009 16255 20043
rect 16773 20009 16807 20043
rect 17325 20009 17359 20043
rect 17877 20009 17911 20043
rect 18521 20009 18555 20043
rect 19073 20009 19107 20043
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 3525 19873 3559 19907
rect 4445 19873 4479 19907
rect 5641 19873 5675 19907
rect 9045 19873 9079 19907
rect 10149 19873 10183 19907
rect 11989 19873 12023 19907
rect 12817 19873 12851 19907
rect 13369 19873 13403 19907
rect 13645 19873 13679 19907
rect 14105 19873 14139 19907
rect 14657 19873 14691 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 16589 19873 16623 19907
rect 17141 19873 17175 19907
rect 17693 19873 17727 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 4721 19805 4755 19839
rect 5917 19805 5951 19839
rect 9321 19805 9355 19839
rect 10241 19805 10275 19839
rect 10425 19805 10459 19839
rect 2513 19737 2547 19771
rect 8677 19737 8711 19771
rect 12173 19737 12207 19771
rect 4077 19669 4111 19703
rect 9781 19669 9815 19703
rect 2421 19329 2455 19363
rect 13001 19329 13035 19363
rect 13921 19329 13955 19363
rect 16129 19329 16163 19363
rect 17049 19329 17083 19363
rect 18337 19329 18371 19363
rect 1685 19261 1719 19295
rect 2237 19261 2271 19295
rect 3249 19261 3283 19295
rect 5089 19261 5123 19295
rect 7757 19261 7791 19295
rect 9413 19261 9447 19295
rect 10057 19261 10091 19295
rect 10324 19261 10358 19295
rect 11805 19261 11839 19295
rect 12817 19261 12851 19295
rect 13645 19261 13679 19295
rect 14657 19261 14691 19295
rect 14933 19261 14967 19295
rect 15393 19261 15427 19295
rect 15945 19261 15979 19295
rect 16773 19261 16807 19295
rect 18061 19261 18095 19295
rect 18797 19261 18831 19295
rect 19993 19261 20027 19295
rect 3516 19193 3550 19227
rect 5356 19193 5390 19227
rect 8024 19193 8058 19227
rect 20637 19193 20671 19227
rect 1869 19125 1903 19159
rect 4629 19125 4663 19159
rect 6469 19125 6503 19159
rect 9137 19125 9171 19159
rect 11437 19125 11471 19159
rect 11989 19125 12023 19159
rect 15577 19125 15611 19159
rect 18981 19125 19015 19159
rect 1593 18921 1627 18955
rect 3433 18921 3467 18955
rect 4077 18921 4111 18955
rect 4445 18921 4479 18955
rect 4537 18921 4571 18955
rect 6837 18921 6871 18955
rect 13645 18921 13679 18955
rect 14105 18921 14139 18955
rect 15301 18921 15335 18955
rect 2237 18853 2271 18887
rect 5724 18853 5758 18887
rect 12081 18853 12115 18887
rect 12817 18853 12851 18887
rect 16589 18853 16623 18887
rect 18337 18853 18371 18887
rect 19073 18853 19107 18887
rect 1409 18785 1443 18819
rect 1961 18785 1995 18819
rect 3341 18785 3375 18819
rect 7205 18785 7239 18819
rect 8033 18785 8067 18819
rect 8677 18785 8711 18819
rect 10416 18785 10450 18819
rect 11805 18785 11839 18819
rect 12541 18785 12575 18819
rect 14013 18785 14047 18819
rect 15669 18785 15703 18819
rect 16313 18785 16347 18819
rect 17325 18785 17359 18819
rect 18061 18785 18095 18819
rect 18797 18785 18831 18819
rect 3525 18717 3559 18751
rect 4629 18717 4663 18751
rect 5457 18717 5491 18751
rect 8125 18717 8159 18751
rect 8217 18717 8251 18751
rect 8861 18717 8895 18751
rect 10149 18717 10183 18751
rect 14289 18717 14323 18751
rect 15761 18717 15795 18751
rect 15945 18717 15979 18751
rect 17601 18717 17635 18751
rect 2973 18581 3007 18615
rect 7665 18581 7699 18615
rect 11529 18581 11563 18615
rect 5273 18377 5307 18411
rect 8217 18377 8251 18411
rect 11437 18377 11471 18411
rect 15209 18377 15243 18411
rect 5733 18241 5767 18275
rect 5917 18241 5951 18275
rect 8769 18241 8803 18275
rect 15853 18241 15887 18275
rect 1593 18173 1627 18207
rect 2145 18173 2179 18207
rect 2973 18173 3007 18207
rect 7113 18173 7147 18207
rect 8677 18173 8711 18207
rect 10057 18173 10091 18207
rect 13185 18173 13219 18207
rect 15025 18173 15059 18207
rect 15669 18173 15703 18207
rect 2421 18105 2455 18139
rect 3240 18105 3274 18139
rect 5641 18105 5675 18139
rect 6285 18105 6319 18139
rect 7389 18105 7423 18139
rect 10324 18105 10358 18139
rect 13452 18105 13486 18139
rect 1777 18037 1811 18071
rect 4353 18037 4387 18071
rect 8585 18037 8619 18071
rect 14565 18037 14599 18071
rect 15577 18037 15611 18071
rect 1961 17833 1995 17867
rect 3065 17833 3099 17867
rect 3433 17833 3467 17867
rect 6745 17833 6779 17867
rect 8585 17833 8619 17867
rect 10149 17833 10183 17867
rect 16957 17833 16991 17867
rect 17785 17833 17819 17867
rect 7297 17765 7331 17799
rect 9045 17765 9079 17799
rect 13820 17765 13854 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 2881 17697 2915 17731
rect 5632 17697 5666 17731
rect 7021 17697 7055 17731
rect 8953 17697 8987 17731
rect 10057 17697 10091 17731
rect 15844 17697 15878 17731
rect 18153 17697 18187 17731
rect 5365 17629 5399 17663
rect 9229 17629 9263 17663
rect 10333 17629 10367 17663
rect 13093 17629 13127 17663
rect 13553 17629 13587 17663
rect 15577 17629 15611 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 2513 17493 2547 17527
rect 9689 17493 9723 17527
rect 14933 17493 14967 17527
rect 5641 17289 5675 17323
rect 10977 17289 11011 17323
rect 12449 17289 12483 17323
rect 13461 17289 13495 17323
rect 15393 17289 15427 17323
rect 18061 17289 18095 17323
rect 2237 17153 2271 17187
rect 3065 17153 3099 17187
rect 6101 17153 6135 17187
rect 6193 17153 6227 17187
rect 7389 17153 7423 17187
rect 13001 17153 13035 17187
rect 14105 17153 14139 17187
rect 15945 17153 15979 17187
rect 18613 17153 18647 17187
rect 19073 17153 19107 17187
rect 1501 17085 1535 17119
rect 2053 17085 2087 17119
rect 7656 17085 7690 17119
rect 9597 17085 9631 17119
rect 13829 17085 13863 17119
rect 15761 17085 15795 17119
rect 18521 17085 18555 17119
rect 3332 17017 3366 17051
rect 9864 17017 9898 17051
rect 13921 17017 13955 17051
rect 18429 17017 18463 17051
rect 18889 17017 18923 17051
rect 1685 16949 1719 16983
rect 4445 16949 4479 16983
rect 6009 16949 6043 16983
rect 8769 16949 8803 16983
rect 12817 16949 12851 16983
rect 12909 16949 12943 16983
rect 15853 16949 15887 16983
rect 16957 16949 16991 16983
rect 2881 16745 2915 16779
rect 6377 16745 6411 16779
rect 9781 16745 9815 16779
rect 13829 16745 13863 16779
rect 15945 16745 15979 16779
rect 16313 16745 16347 16779
rect 18337 16745 18371 16779
rect 19993 16745 20027 16779
rect 2329 16677 2363 16711
rect 10784 16677 10818 16711
rect 18858 16677 18892 16711
rect 1501 16609 1535 16643
rect 2063 16609 2097 16643
rect 3249 16609 3283 16643
rect 3341 16609 3375 16643
rect 5264 16609 5298 16643
rect 6653 16609 6687 16643
rect 7380 16609 7414 16643
rect 8953 16609 8987 16643
rect 10517 16609 10551 16643
rect 12173 16609 12207 16643
rect 12440 16609 12474 16643
rect 14197 16609 14231 16643
rect 17224 16609 17258 16643
rect 3525 16541 3559 16575
rect 4997 16541 5031 16575
rect 7113 16541 7147 16575
rect 14289 16541 14323 16575
rect 14381 16541 14415 16575
rect 16405 16541 16439 16575
rect 16589 16541 16623 16575
rect 16957 16541 16991 16575
rect 18613 16541 18647 16575
rect 1685 16473 1719 16507
rect 8769 16473 8803 16507
rect 8493 16405 8527 16439
rect 11897 16405 11931 16439
rect 13553 16405 13587 16439
rect 4261 16201 4295 16235
rect 5273 16201 5307 16235
rect 10241 16201 10275 16235
rect 12449 16201 12483 16235
rect 13921 16201 13955 16235
rect 17417 16201 17451 16235
rect 2053 16065 2087 16099
rect 4721 16065 4755 16099
rect 4813 16065 4847 16099
rect 5825 16065 5859 16099
rect 7941 16065 7975 16099
rect 8125 16065 8159 16099
rect 8861 16065 8895 16099
rect 13001 16065 13035 16099
rect 14381 16065 14415 16099
rect 14565 16065 14599 16099
rect 16037 16065 16071 16099
rect 1869 15997 1903 16031
rect 2605 15997 2639 16031
rect 2872 15997 2906 16031
rect 6469 15997 6503 16031
rect 10517 15997 10551 16031
rect 10784 15997 10818 16031
rect 12909 15997 12943 16031
rect 14289 15997 14323 16031
rect 7849 15929 7883 15963
rect 9128 15929 9162 15963
rect 12817 15929 12851 15963
rect 13461 15929 13495 15963
rect 16304 15929 16338 15963
rect 3985 15861 4019 15895
rect 4629 15861 4663 15895
rect 5641 15861 5675 15895
rect 5733 15861 5767 15895
rect 6285 15861 6319 15895
rect 7481 15861 7515 15895
rect 11897 15861 11931 15895
rect 1593 15657 1627 15691
rect 3157 15657 3191 15691
rect 6377 15657 6411 15691
rect 6837 15657 6871 15691
rect 7297 15657 7331 15691
rect 8953 15657 8987 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 12173 15657 12207 15691
rect 12633 15657 12667 15691
rect 13645 15657 13679 15691
rect 14657 15657 14691 15691
rect 15853 15657 15887 15691
rect 2237 15589 2271 15623
rect 7205 15589 7239 15623
rect 10057 15589 10091 15623
rect 11529 15589 11563 15623
rect 1409 15521 1443 15555
rect 1971 15521 2005 15555
rect 4988 15521 5022 15555
rect 8033 15521 8067 15555
rect 8861 15521 8895 15555
rect 11437 15521 11471 15555
rect 12541 15521 12575 15555
rect 13369 15521 13403 15555
rect 14013 15521 14047 15555
rect 14841 15521 14875 15555
rect 16221 15521 16255 15555
rect 17049 15521 17083 15555
rect 4721 15453 4755 15487
rect 7481 15453 7515 15487
rect 9137 15453 9171 15487
rect 10241 15453 10275 15487
rect 11621 15453 11655 15487
rect 12817 15453 12851 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 16313 15453 16347 15487
rect 16497 15453 16531 15487
rect 8493 15385 8527 15419
rect 16865 15385 16899 15419
rect 6101 15317 6135 15351
rect 11069 15317 11103 15351
rect 13185 15317 13219 15351
rect 5641 15113 5675 15147
rect 9873 15113 9907 15147
rect 13093 15113 13127 15147
rect 15669 15113 15703 15147
rect 17417 15113 17451 15147
rect 2789 14977 2823 15011
rect 6285 14977 6319 15011
rect 6837 14977 6871 15011
rect 8493 14977 8527 15011
rect 11621 14977 11655 15011
rect 13737 14977 13771 15011
rect 16037 14977 16071 15011
rect 1409 14909 1443 14943
rect 1961 14909 1995 14943
rect 3056 14909 3090 14943
rect 6101 14909 6135 14943
rect 7104 14909 7138 14943
rect 8760 14909 8794 14943
rect 11529 14909 11563 14943
rect 14289 14909 14323 14943
rect 14545 14909 14579 14943
rect 18153 14909 18187 14943
rect 2237 14841 2271 14875
rect 6009 14841 6043 14875
rect 11437 14841 11471 14875
rect 16304 14841 16338 14875
rect 18420 14841 18454 14875
rect 1593 14773 1627 14807
rect 4169 14773 4203 14807
rect 8217 14773 8251 14807
rect 11069 14773 11103 14807
rect 13461 14773 13495 14807
rect 13553 14773 13587 14807
rect 19533 14773 19567 14807
rect 1777 14569 1811 14603
rect 4537 14569 4571 14603
rect 7665 14569 7699 14603
rect 14565 14569 14599 14603
rect 15669 14569 15703 14603
rect 17049 14569 17083 14603
rect 2421 14501 2455 14535
rect 4445 14501 4479 14535
rect 10692 14501 10726 14535
rect 17417 14501 17451 14535
rect 18328 14501 18362 14535
rect 1593 14433 1627 14467
rect 2145 14433 2179 14467
rect 6009 14433 6043 14467
rect 6276 14433 6310 14467
rect 7849 14433 7883 14467
rect 10425 14433 10459 14467
rect 13185 14433 13219 14467
rect 13441 14433 13475 14467
rect 15761 14433 15795 14467
rect 18061 14433 18095 14467
rect 3341 14365 3375 14399
rect 4629 14365 4663 14399
rect 5549 14365 5583 14399
rect 15945 14365 15979 14399
rect 16497 14365 16531 14399
rect 17509 14365 17543 14399
rect 17693 14365 17727 14399
rect 15301 14297 15335 14331
rect 4077 14229 4111 14263
rect 7389 14229 7423 14263
rect 11805 14229 11839 14263
rect 19441 14229 19475 14263
rect 2513 14025 2547 14059
rect 5733 14025 5767 14059
rect 9413 14025 9447 14059
rect 9781 14025 9815 14059
rect 12633 14025 12667 14059
rect 17049 14025 17083 14059
rect 18061 14025 18095 14059
rect 4905 13957 4939 13991
rect 1961 13889 1995 13923
rect 2973 13889 3007 13923
rect 3157 13889 3191 13923
rect 6377 13889 6411 13923
rect 7481 13889 7515 13923
rect 10425 13889 10459 13923
rect 11253 13889 11287 13923
rect 11437 13889 11471 13923
rect 13277 13889 13311 13923
rect 14289 13889 14323 13923
rect 15209 13889 15243 13923
rect 15669 13889 15703 13923
rect 18705 13889 18739 13923
rect 1777 13821 1811 13855
rect 2881 13821 2915 13855
rect 3525 13821 3559 13855
rect 3792 13821 3826 13855
rect 6101 13821 6135 13855
rect 7297 13821 7331 13855
rect 8033 13821 8067 13855
rect 14105 13821 14139 13855
rect 15117 13821 15151 13855
rect 15936 13821 15970 13855
rect 18429 13821 18463 13855
rect 18889 13821 18923 13855
rect 8300 13753 8334 13787
rect 10149 13753 10183 13787
rect 11161 13753 11195 13787
rect 13001 13753 13035 13787
rect 15025 13753 15059 13787
rect 19073 13753 19107 13787
rect 6193 13685 6227 13719
rect 6837 13685 6871 13719
rect 7205 13685 7239 13719
rect 10241 13685 10275 13719
rect 10793 13685 10827 13719
rect 13093 13685 13127 13719
rect 13645 13685 13679 13719
rect 14013 13685 14047 13719
rect 14657 13685 14691 13719
rect 18521 13685 18555 13719
rect 1593 13481 1627 13515
rect 6561 13481 6595 13515
rect 7757 13481 7791 13515
rect 14197 13481 14231 13515
rect 14473 13481 14507 13515
rect 15669 13481 15703 13515
rect 16681 13481 16715 13515
rect 17141 13481 17175 13515
rect 10793 13413 10827 13447
rect 12541 13413 12575 13447
rect 17049 13413 17083 13447
rect 1409 13345 1443 13379
rect 1961 13345 1995 13379
rect 5448 13345 5482 13379
rect 7389 13345 7423 13379
rect 7941 13345 7975 13379
rect 8401 13345 8435 13379
rect 9045 13345 9079 13379
rect 13084 13345 13118 13379
rect 14657 13345 14691 13379
rect 16037 13345 16071 13379
rect 2145 13277 2179 13311
rect 5181 13277 5215 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 12817 13277 12851 13311
rect 16129 13277 16163 13311
rect 16313 13277 16347 13311
rect 17233 13277 17267 13311
rect 7205 13141 7239 13175
rect 8033 13141 8067 13175
rect 2513 12937 2547 12971
rect 6101 12937 6135 12971
rect 6837 12937 6871 12971
rect 9321 12937 9355 12971
rect 11437 12937 11471 12971
rect 13093 12937 13127 12971
rect 17233 12937 17267 12971
rect 1961 12869 1995 12903
rect 11529 12869 11563 12903
rect 4721 12801 4755 12835
rect 7389 12801 7423 12835
rect 12081 12801 12115 12835
rect 13645 12801 13679 12835
rect 1777 12733 1811 12767
rect 2329 12733 2363 12767
rect 7941 12733 7975 12767
rect 10057 12733 10091 12767
rect 10324 12733 10358 12767
rect 15853 12733 15887 12767
rect 18061 12733 18095 12767
rect 18328 12733 18362 12767
rect 4988 12665 5022 12699
rect 7205 12665 7239 12699
rect 8208 12665 8242 12699
rect 11897 12665 11931 12699
rect 12449 12665 12483 12699
rect 13461 12665 13495 12699
rect 14105 12665 14139 12699
rect 16120 12665 16154 12699
rect 4261 12597 4295 12631
rect 7297 12597 7331 12631
rect 11989 12597 12023 12631
rect 13553 12597 13587 12631
rect 19441 12597 19475 12631
rect 1593 12393 1627 12427
rect 7573 12393 7607 12427
rect 8585 12393 8619 12427
rect 9045 12393 9079 12427
rect 13001 12393 13035 12427
rect 16773 12393 16807 12427
rect 17049 12393 17083 12427
rect 18153 12393 18187 12427
rect 18705 12393 18739 12427
rect 2237 12325 2271 12359
rect 2973 12325 3007 12359
rect 6000 12325 6034 12359
rect 10762 12325 10796 12359
rect 12541 12325 12575 12359
rect 13369 12325 13403 12359
rect 15649 12325 15683 12359
rect 19073 12325 19107 12359
rect 1409 12257 1443 12291
rect 1961 12257 1995 12291
rect 2697 12257 2731 12291
rect 4333 12257 4367 12291
rect 7941 12257 7975 12291
rect 8033 12257 8067 12291
rect 8953 12257 8987 12291
rect 10517 12257 10551 12291
rect 12265 12257 12299 12291
rect 14473 12257 14507 12291
rect 18061 12257 18095 12291
rect 4077 12189 4111 12223
rect 5733 12189 5767 12223
rect 8217 12189 8251 12223
rect 9137 12189 9171 12223
rect 13461 12189 13495 12223
rect 13645 12189 13679 12223
rect 14565 12189 14599 12223
rect 15393 12189 15427 12223
rect 18337 12189 18371 12223
rect 19165 12189 19199 12223
rect 19257 12189 19291 12223
rect 17693 12121 17727 12155
rect 5457 12053 5491 12087
rect 7113 12053 7147 12087
rect 11897 12053 11931 12087
rect 14289 12053 14323 12087
rect 4353 11849 4387 11883
rect 5641 11849 5675 11883
rect 9321 11849 9355 11883
rect 11161 11849 11195 11883
rect 13461 11849 13495 11883
rect 14381 11849 14415 11883
rect 15853 11849 15887 11883
rect 15945 11849 15979 11883
rect 16129 11849 16163 11883
rect 4077 11781 4111 11815
rect 10149 11781 10183 11815
rect 1869 11713 1903 11747
rect 4905 11713 4939 11747
rect 6193 11713 6227 11747
rect 7389 11713 7423 11747
rect 10701 11713 10735 11747
rect 11713 11713 11747 11747
rect 13001 11713 13035 11747
rect 14105 11713 14139 11747
rect 17141 11781 17175 11815
rect 15945 11713 15979 11747
rect 16681 11713 16715 11747
rect 18061 11713 18095 11747
rect 19717 11713 19751 11747
rect 1685 11645 1719 11679
rect 2697 11645 2731 11679
rect 6101 11645 6135 11679
rect 7941 11645 7975 11679
rect 10609 11645 10643 11679
rect 11529 11645 11563 11679
rect 12817 11645 12851 11679
rect 13829 11645 13863 11679
rect 14381 11645 14415 11679
rect 14473 11645 14507 11679
rect 14729 11645 14763 11679
rect 16589 11645 16623 11679
rect 17325 11645 17359 11679
rect 18328 11645 18362 11679
rect 2964 11577 2998 11611
rect 4813 11577 4847 11611
rect 7297 11577 7331 11611
rect 8208 11577 8242 11611
rect 9689 11577 9723 11611
rect 10517 11577 10551 11611
rect 12909 11577 12943 11611
rect 19984 11577 20018 11611
rect 4721 11509 4755 11543
rect 6009 11509 6043 11543
rect 6837 11509 6871 11543
rect 7205 11509 7239 11543
rect 11621 11509 11655 11543
rect 12449 11509 12483 11543
rect 13921 11509 13955 11543
rect 16497 11509 16531 11543
rect 17509 11509 17543 11543
rect 19441 11509 19475 11543
rect 21097 11509 21131 11543
rect 1593 11305 1627 11339
rect 4077 11305 4111 11339
rect 9045 11305 9079 11339
rect 11897 11305 11931 11339
rect 14933 11305 14967 11339
rect 15301 11305 15335 11339
rect 15761 11305 15795 11339
rect 17785 11305 17819 11339
rect 18153 11305 18187 11339
rect 7021 11237 7055 11271
rect 9689 11237 9723 11271
rect 12357 11237 12391 11271
rect 1409 11169 1443 11203
rect 1961 11169 1995 11203
rect 3249 11169 3283 11203
rect 4445 11169 4479 11203
rect 5089 11169 5123 11203
rect 5733 11169 5767 11203
rect 7932 11169 7966 11203
rect 10508 11169 10542 11203
rect 12265 11169 12299 11203
rect 13093 11169 13127 11203
rect 13820 11169 13854 11203
rect 15669 11169 15703 11203
rect 2145 11101 2179 11135
rect 3341 11101 3375 11135
rect 3525 11101 3559 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 7113 11101 7147 11135
rect 7297 11101 7331 11135
rect 7665 11101 7699 11135
rect 10241 11101 10275 11135
rect 12449 11101 12483 11135
rect 13553 11101 13587 11135
rect 15853 11101 15887 11135
rect 18245 11101 18279 11135
rect 18429 11101 18463 11135
rect 6653 11033 6687 11067
rect 11621 11033 11655 11067
rect 12909 11033 12943 11067
rect 17601 11033 17635 11067
rect 2881 10965 2915 10999
rect 5549 10965 5583 10999
rect 2053 10761 2087 10795
rect 4077 10761 4111 10795
rect 8493 10761 8527 10795
rect 12081 10761 12115 10795
rect 14381 10761 14415 10795
rect 16497 10761 16531 10795
rect 8217 10693 8251 10727
rect 12265 10693 12299 10727
rect 15485 10693 15519 10727
rect 2697 10625 2731 10659
rect 3709 10625 3743 10659
rect 4721 10625 4755 10659
rect 6837 10625 6871 10659
rect 9045 10625 9079 10659
rect 10701 10625 10735 10659
rect 2513 10557 2547 10591
rect 4537 10557 4571 10591
rect 8861 10557 8895 10591
rect 15945 10625 15979 10659
rect 16129 10625 16163 10659
rect 16957 10625 16991 10659
rect 17049 10625 17083 10659
rect 18061 10625 18095 10659
rect 13001 10557 13035 10591
rect 18328 10557 18362 10591
rect 7104 10489 7138 10523
rect 10968 10489 11002 10523
rect 12265 10489 12299 10523
rect 13268 10489 13302 10523
rect 15853 10489 15887 10523
rect 2421 10421 2455 10455
rect 3065 10421 3099 10455
rect 3433 10421 3467 10455
rect 3525 10421 3559 10455
rect 4445 10421 4479 10455
rect 8953 10421 8987 10455
rect 16865 10421 16899 10455
rect 19441 10421 19475 10455
rect 3433 10217 3467 10251
rect 13369 10217 13403 10251
rect 13645 10217 13679 10251
rect 2044 10149 2078 10183
rect 8309 10149 8343 10183
rect 12234 10149 12268 10183
rect 1777 10081 1811 10115
rect 4077 10081 4111 10115
rect 4344 10081 4378 10115
rect 5733 10081 5767 10115
rect 6000 10081 6034 10115
rect 7849 10081 7883 10115
rect 8401 10081 8435 10115
rect 11989 10081 12023 10115
rect 14013 10081 14047 10115
rect 16221 10081 16255 10115
rect 16488 10081 16522 10115
rect 8585 10013 8619 10047
rect 14105 10013 14139 10047
rect 14197 10013 14231 10047
rect 3157 9877 3191 9911
rect 5457 9877 5491 9911
rect 7113 9877 7147 9911
rect 7665 9877 7699 9911
rect 7941 9877 7975 9911
rect 17601 9877 17635 9911
rect 3157 9673 3191 9707
rect 17049 9673 17083 9707
rect 4169 9605 4203 9639
rect 5733 9605 5767 9639
rect 10057 9605 10091 9639
rect 10333 9605 10367 9639
rect 3801 9537 3835 9571
rect 4813 9537 4847 9571
rect 6377 9537 6411 9571
rect 7481 9537 7515 9571
rect 10885 9537 10919 9571
rect 13369 9537 13403 9571
rect 17325 9537 17359 9571
rect 6193 9469 6227 9503
rect 8677 9469 8711 9503
rect 8944 9469 8978 9503
rect 15669 9469 15703 9503
rect 3525 9401 3559 9435
rect 4537 9401 4571 9435
rect 6101 9401 6135 9435
rect 10793 9401 10827 9435
rect 15936 9401 15970 9435
rect 3617 9333 3651 9367
rect 4629 9333 4663 9367
rect 6837 9333 6871 9367
rect 7205 9333 7239 9367
rect 7297 9333 7331 9367
rect 10701 9333 10735 9367
rect 1961 9129 1995 9163
rect 4721 9129 4755 9163
rect 5273 9129 5307 9163
rect 6377 9129 6411 9163
rect 9689 9129 9723 9163
rect 1777 8993 1811 9027
rect 5181 8993 5215 9027
rect 8197 8993 8231 9027
rect 10057 8993 10091 9027
rect 5365 8925 5399 8959
rect 7941 8925 7975 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 9321 8857 9355 8891
rect 4813 8789 4847 8823
rect 8585 8585 8619 8619
rect 1685 8449 1719 8483
rect 4721 8449 4755 8483
rect 5733 8449 5767 8483
rect 7205 8449 7239 8483
rect 9413 8449 9447 8483
rect 1409 8381 1443 8415
rect 2145 8381 2179 8415
rect 2412 8381 2446 8415
rect 4629 8381 4663 8415
rect 9229 8381 9263 8415
rect 9321 8381 9355 8415
rect 4537 8313 4571 8347
rect 5549 8313 5583 8347
rect 5641 8313 5675 8347
rect 7472 8313 7506 8347
rect 3525 8245 3559 8279
rect 4169 8245 4203 8279
rect 5181 8245 5215 8279
rect 8861 8245 8895 8279
rect 1777 8041 1811 8075
rect 4537 8041 4571 8075
rect 8953 8041 8987 8075
rect 18613 8041 18647 8075
rect 1593 7905 1627 7939
rect 2053 7905 2087 7939
rect 2155 7905 2189 7939
rect 4445 7905 4479 7939
rect 5448 7905 5482 7939
rect 7104 7905 7138 7939
rect 8861 7905 8895 7939
rect 18429 7905 18463 7939
rect 2329 7837 2363 7871
rect 4721 7837 4755 7871
rect 5181 7837 5215 7871
rect 6837 7837 6871 7871
rect 9045 7837 9079 7871
rect 6561 7769 6595 7803
rect 2053 7701 2087 7735
rect 4077 7701 4111 7735
rect 8217 7701 8251 7735
rect 8493 7701 8527 7735
rect 6009 7497 6043 7531
rect 8401 7497 8435 7531
rect 19165 7497 19199 7531
rect 8125 7361 8159 7395
rect 2973 7293 3007 7327
rect 4629 7293 4663 7327
rect 9137 7361 9171 7395
rect 8953 7293 8987 7327
rect 18981 7293 19015 7327
rect 3240 7225 3274 7259
rect 4874 7225 4908 7259
rect 7021 7225 7055 7259
rect 7849 7225 7883 7259
rect 8401 7225 8435 7259
rect 8861 7225 8895 7259
rect 4353 7157 4387 7191
rect 7481 7157 7515 7191
rect 7941 7157 7975 7191
rect 8493 7157 8527 7191
rect 7573 6953 7607 6987
rect 8309 6953 8343 6987
rect 4445 6817 4479 6851
rect 5089 6817 5123 6851
rect 7665 6817 7699 6851
rect 8677 6817 8711 6851
rect 19441 6817 19475 6851
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 7757 6749 7791 6783
rect 8769 6749 8803 6783
rect 8953 6749 8987 6783
rect 4077 6681 4111 6715
rect 19625 6681 19659 6715
rect 7205 6613 7239 6647
rect 20085 6409 20119 6443
rect 19901 6205 19935 6239
rect 20453 5865 20487 5899
rect 20269 5729 20303 5763
rect 20729 5321 20763 5355
rect 20545 5117 20579 5151
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2866 20040 2872 20052
rect 1995 20012 2872 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 5261 20043 5319 20049
rect 5261 20040 5273 20043
rect 4571 20012 5273 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 5261 20009 5273 20012
rect 5307 20009 5319 20043
rect 5261 20003 5319 20009
rect 5626 20000 5632 20052
rect 5684 20040 5690 20052
rect 5721 20043 5779 20049
rect 5721 20040 5733 20043
rect 5684 20012 5733 20040
rect 5684 20000 5690 20012
rect 5721 20009 5733 20012
rect 5767 20009 5779 20043
rect 5721 20003 5779 20009
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9306 20040 9312 20052
rect 9171 20012 9312 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9306 20000 9312 20012
rect 9364 20000 9370 20052
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 12989 20043 13047 20049
rect 12989 20040 13001 20043
rect 12952 20012 13001 20040
rect 12952 20000 12958 20012
rect 12989 20009 13001 20012
rect 13035 20009 13047 20043
rect 12989 20003 13047 20009
rect 13354 20000 13360 20052
rect 13412 20040 13418 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 13412 20012 14289 20040
rect 13412 20000 13418 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 14829 20043 14887 20049
rect 14829 20009 14841 20043
rect 14875 20040 14887 20043
rect 15194 20040 15200 20052
rect 14875 20012 15200 20040
rect 14875 20009 14887 20012
rect 14829 20003 14887 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15654 20040 15660 20052
rect 15615 20012 15660 20040
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16209 20043 16267 20049
rect 16209 20040 16221 20043
rect 16172 20012 16221 20040
rect 16172 20000 16178 20012
rect 16209 20009 16221 20012
rect 16255 20009 16267 20043
rect 16209 20003 16267 20009
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16761 20043 16819 20049
rect 16761 20040 16773 20043
rect 16632 20012 16773 20040
rect 16632 20000 16638 20012
rect 16761 20009 16773 20012
rect 16807 20009 16819 20043
rect 16761 20003 16819 20009
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 17313 20043 17371 20049
rect 17313 20040 17325 20043
rect 17092 20012 17325 20040
rect 17092 20000 17098 20012
rect 17313 20009 17325 20012
rect 17359 20009 17371 20043
rect 17313 20003 17371 20009
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 17865 20043 17923 20049
rect 17865 20040 17877 20043
rect 17552 20012 17877 20040
rect 17552 20000 17558 20012
rect 17865 20009 17877 20012
rect 17911 20009 17923 20043
rect 17865 20003 17923 20009
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18472 20012 18521 20040
rect 18472 20000 18478 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18509 20003 18567 20009
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 19061 20043 19119 20049
rect 19061 20040 19073 20043
rect 18932 20012 19073 20040
rect 18932 20000 18938 20012
rect 19061 20009 19073 20012
rect 19107 20009 19119 20043
rect 19061 20003 19119 20009
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 3513 19907 3571 19913
rect 3513 19873 3525 19907
rect 3559 19904 3571 19907
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3559 19876 4445 19904
rect 3559 19873 3571 19876
rect 3513 19867 3571 19873
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19904 5687 19907
rect 5994 19904 6000 19916
rect 5675 19876 6000 19904
rect 5675 19873 5687 19876
rect 5629 19867 5687 19873
rect 5994 19864 6000 19876
rect 6052 19904 6058 19916
rect 9033 19907 9091 19913
rect 9033 19904 9045 19907
rect 6052 19876 9045 19904
rect 6052 19864 6058 19876
rect 9033 19873 9045 19876
rect 9079 19873 9091 19907
rect 9033 19867 9091 19873
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9732 19876 10149 19904
rect 9732 19864 9738 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 11974 19904 11980 19916
rect 11935 19876 11980 19904
rect 10137 19867 10195 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12805 19907 12863 19913
rect 12805 19873 12817 19907
rect 12851 19904 12863 19907
rect 12986 19904 12992 19916
rect 12851 19876 12992 19904
rect 12851 19873 12863 19876
rect 12805 19867 12863 19873
rect 12986 19864 12992 19876
rect 13044 19864 13050 19916
rect 13354 19904 13360 19916
rect 13315 19876 13360 19904
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13679 19876 14105 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 14366 19864 14372 19916
rect 14424 19904 14430 19916
rect 14645 19907 14703 19913
rect 14645 19904 14657 19907
rect 14424 19876 14657 19904
rect 14424 19864 14430 19876
rect 14645 19873 14657 19876
rect 14691 19873 14703 19907
rect 14645 19867 14703 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 15252 19876 15485 19904
rect 15252 19864 15258 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16114 19904 16120 19916
rect 16071 19876 16120 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 16574 19904 16580 19916
rect 16535 19876 16580 19904
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 17126 19904 17132 19916
rect 17087 19876 17132 19904
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19904 17739 19907
rect 17954 19904 17960 19916
rect 17727 19876 17960 19904
rect 17727 19873 17739 19876
rect 17681 19867 17739 19873
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18506 19904 18512 19916
rect 18371 19876 18512 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18506 19864 18512 19876
rect 18564 19864 18570 19916
rect 18874 19904 18880 19916
rect 18835 19876 18880 19904
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4890 19836 4896 19848
rect 4755 19808 4896 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5902 19836 5908 19848
rect 5863 19808 5908 19836
rect 5902 19796 5908 19808
rect 5960 19796 5966 19848
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 9950 19836 9956 19848
rect 9355 19808 9956 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19805 10287 19839
rect 10410 19836 10416 19848
rect 10371 19808 10416 19836
rect 10229 19799 10287 19805
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19768 2559 19771
rect 2774 19768 2780 19780
rect 2547 19740 2780 19768
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 2774 19728 2780 19740
rect 2832 19728 2838 19780
rect 8665 19771 8723 19777
rect 8665 19737 8677 19771
rect 8711 19768 8723 19771
rect 10244 19768 10272 19799
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 8711 19740 10272 19768
rect 12161 19771 12219 19777
rect 8711 19737 8723 19740
rect 8665 19731 8723 19737
rect 12161 19737 12173 19771
rect 12207 19768 12219 19771
rect 14274 19768 14280 19780
rect 12207 19740 14280 19768
rect 12207 19737 12219 19740
rect 12161 19731 12219 19737
rect 14274 19728 14280 19740
rect 14332 19728 14338 19780
rect 2222 19660 2228 19712
rect 2280 19700 2286 19712
rect 4065 19703 4123 19709
rect 4065 19700 4077 19703
rect 2280 19672 4077 19700
rect 2280 19660 2286 19672
rect 4065 19669 4077 19672
rect 4111 19669 4123 19703
rect 9766 19700 9772 19712
rect 9727 19672 9772 19700
rect 4065 19663 4123 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 3476 19468 5028 19496
rect 3476 19456 3482 19468
rect 1762 19320 1768 19372
rect 1820 19360 1826 19372
rect 2409 19363 2467 19369
rect 2409 19360 2421 19363
rect 1820 19332 2421 19360
rect 1820 19320 1826 19332
rect 2409 19329 2421 19332
rect 2455 19329 2467 19363
rect 5000 19360 5028 19468
rect 17862 19388 17868 19440
rect 17920 19428 17926 19440
rect 18046 19428 18052 19440
rect 17920 19400 18052 19428
rect 17920 19388 17926 19400
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 2409 19323 2467 19329
rect 4264 19332 4936 19360
rect 5000 19332 5212 19360
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 3237 19295 3295 19301
rect 3237 19292 3249 19295
rect 2924 19264 3249 19292
rect 2924 19252 2930 19264
rect 3237 19261 3249 19264
rect 3283 19292 3295 19295
rect 4264 19292 4292 19332
rect 3283 19264 4292 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 4338 19252 4344 19304
rect 4396 19292 4402 19304
rect 4798 19292 4804 19304
rect 4396 19264 4804 19292
rect 4396 19252 4402 19264
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 4908 19292 4936 19332
rect 5074 19292 5080 19304
rect 4908 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5184 19292 5212 19332
rect 9950 19320 9956 19372
rect 10008 19360 10014 19372
rect 12986 19360 12992 19372
rect 10008 19332 10180 19360
rect 12947 19332 12992 19360
rect 10008 19320 10014 19332
rect 7374 19292 7380 19304
rect 5184 19264 7380 19292
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7745 19295 7803 19301
rect 7745 19261 7757 19295
rect 7791 19261 7803 19295
rect 7745 19255 7803 19261
rect 9401 19295 9459 19301
rect 9401 19261 9413 19295
rect 9447 19292 9459 19295
rect 9674 19292 9680 19304
rect 9447 19264 9680 19292
rect 9447 19261 9459 19264
rect 9401 19255 9459 19261
rect 198 19184 204 19236
rect 256 19224 262 19236
rect 3142 19224 3148 19236
rect 256 19196 3148 19224
rect 256 19184 262 19196
rect 3142 19184 3148 19196
rect 3200 19184 3206 19236
rect 3504 19227 3562 19233
rect 3504 19193 3516 19227
rect 3550 19224 3562 19227
rect 5344 19227 5402 19233
rect 3550 19196 4936 19224
rect 3550 19193 3562 19196
rect 3504 19187 3562 19193
rect 4908 19168 4936 19196
rect 5344 19193 5356 19227
rect 5390 19224 5402 19227
rect 5902 19224 5908 19236
rect 5390 19196 5908 19224
rect 5390 19193 5402 19196
rect 5344 19187 5402 19193
rect 5902 19184 5908 19196
rect 5960 19224 5966 19236
rect 6822 19224 6828 19236
rect 5960 19196 6828 19224
rect 5960 19184 5966 19196
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 7282 19184 7288 19236
rect 7340 19224 7346 19236
rect 7760 19224 7788 19255
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 10042 19292 10048 19304
rect 10003 19264 10048 19292
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 10152 19292 10180 19332
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 14366 19360 14372 19372
rect 13955 19332 14372 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 16114 19360 16120 19372
rect 16075 19332 16120 19360
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19360 17095 19363
rect 17126 19360 17132 19372
rect 17083 19332 17132 19360
rect 17083 19329 17095 19332
rect 17037 19323 17095 19329
rect 17126 19320 17132 19332
rect 17184 19320 17190 19372
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18506 19360 18512 19372
rect 18371 19332 18512 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 10318 19301 10324 19304
rect 10312 19292 10324 19301
rect 10152 19264 10324 19292
rect 10312 19255 10324 19264
rect 10318 19252 10324 19255
rect 10376 19252 10382 19304
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 12158 19292 12164 19304
rect 11839 19264 12164 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 13170 19292 13176 19304
rect 12851 19264 13176 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 13722 19292 13728 19304
rect 13679 19264 13728 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 14148 19264 14657 19292
rect 14148 19252 14154 19264
rect 14645 19261 14657 19264
rect 14691 19261 14703 19295
rect 14645 19255 14703 19261
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19292 14979 19295
rect 15194 19292 15200 19304
rect 14967 19264 15200 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15378 19292 15384 19304
rect 15339 19264 15384 19292
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15804 19264 15945 19292
rect 15804 19252 15810 19264
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 16758 19292 16764 19304
rect 16719 19264 16764 19292
rect 15933 19255 15991 19261
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18690 19292 18696 19304
rect 18095 19264 18696 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 18690 19252 18696 19264
rect 18748 19252 18754 19304
rect 18785 19295 18843 19301
rect 18785 19261 18797 19295
rect 18831 19292 18843 19295
rect 19058 19292 19064 19304
rect 18831 19264 19064 19292
rect 18831 19261 18843 19264
rect 18785 19255 18843 19261
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 19981 19295 20039 19301
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 22094 19292 22100 19304
rect 20027 19264 22100 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 7340 19196 7788 19224
rect 8012 19227 8070 19233
rect 7340 19184 7346 19196
rect 8012 19193 8024 19227
rect 8058 19224 8070 19227
rect 8754 19224 8760 19236
rect 8058 19196 8760 19224
rect 8058 19193 8070 19196
rect 8012 19187 8070 19193
rect 8754 19184 8760 19196
rect 8812 19184 8818 19236
rect 13906 19224 13912 19236
rect 10336 19196 13912 19224
rect 1857 19159 1915 19165
rect 1857 19125 1869 19159
rect 1903 19156 1915 19159
rect 2958 19156 2964 19168
rect 1903 19128 2964 19156
rect 1903 19125 1915 19128
rect 1857 19119 1915 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 4246 19116 4252 19168
rect 4304 19156 4310 19168
rect 4617 19159 4675 19165
rect 4617 19156 4629 19159
rect 4304 19128 4629 19156
rect 4304 19116 4310 19128
rect 4617 19125 4629 19128
rect 4663 19125 4675 19159
rect 4617 19119 4675 19125
rect 4890 19116 4896 19168
rect 4948 19156 4954 19168
rect 6457 19159 6515 19165
rect 6457 19156 6469 19159
rect 4948 19128 6469 19156
rect 4948 19116 4954 19128
rect 6457 19125 6469 19128
rect 6503 19125 6515 19159
rect 6457 19119 6515 19125
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 9125 19159 9183 19165
rect 9125 19156 9137 19159
rect 8260 19128 9137 19156
rect 8260 19116 8266 19128
rect 9125 19125 9137 19128
rect 9171 19125 9183 19159
rect 9125 19119 9183 19125
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 10336 19156 10364 19196
rect 13906 19184 13912 19196
rect 13964 19184 13970 19236
rect 20622 19224 20628 19236
rect 20583 19196 20628 19224
rect 20622 19184 20628 19196
rect 20680 19184 20686 19236
rect 9272 19128 10364 19156
rect 9272 19116 9278 19128
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 11425 19159 11483 19165
rect 11425 19156 11437 19159
rect 10468 19128 11437 19156
rect 10468 19116 10474 19128
rect 11425 19125 11437 19128
rect 11471 19125 11483 19159
rect 11425 19119 11483 19125
rect 11977 19159 12035 19165
rect 11977 19125 11989 19159
rect 12023 19156 12035 19159
rect 13814 19156 13820 19168
rect 12023 19128 13820 19156
rect 12023 19125 12035 19128
rect 11977 19119 12035 19125
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 15010 19116 15016 19168
rect 15068 19156 15074 19168
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 15068 19128 15577 19156
rect 15068 19116 15074 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 15565 19119 15623 19125
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18104 19128 18981 19156
rect 18104 19116 18110 19128
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 18969 19119 19027 19125
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 3421 18955 3479 18961
rect 1872 18924 3096 18952
rect 1026 18844 1032 18896
rect 1084 18884 1090 18896
rect 1872 18884 1900 18924
rect 1084 18856 1900 18884
rect 2225 18887 2283 18893
rect 1084 18844 1090 18856
rect 2225 18853 2237 18887
rect 2271 18884 2283 18887
rect 2314 18884 2320 18896
rect 2271 18856 2320 18884
rect 2271 18853 2283 18856
rect 2225 18847 2283 18853
rect 2314 18844 2320 18856
rect 2372 18844 2378 18896
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18785 1455 18819
rect 1946 18816 1952 18828
rect 1907 18788 1952 18816
rect 1397 18779 1455 18785
rect 1412 18748 1440 18779
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 2038 18748 2044 18760
rect 1412 18720 2044 18748
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 2961 18615 3019 18621
rect 2961 18612 2973 18615
rect 2188 18584 2973 18612
rect 2188 18572 2194 18584
rect 2961 18581 2973 18584
rect 3007 18581 3019 18615
rect 3068 18612 3096 18924
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 4065 18955 4123 18961
rect 4065 18952 4077 18955
rect 3467 18924 4077 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 4065 18921 4077 18924
rect 4111 18921 4123 18955
rect 4430 18952 4436 18964
rect 4391 18924 4436 18952
rect 4065 18915 4123 18921
rect 4430 18912 4436 18924
rect 4488 18912 4494 18964
rect 4525 18955 4583 18961
rect 4525 18921 4537 18955
rect 4571 18952 4583 18955
rect 5166 18952 5172 18964
rect 4571 18924 5172 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 6822 18952 6828 18964
rect 6783 18924 6828 18952
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 6932 18924 13308 18952
rect 3142 18844 3148 18896
rect 3200 18884 3206 18896
rect 5712 18887 5770 18893
rect 3200 18856 4568 18884
rect 3200 18844 3206 18856
rect 3326 18816 3332 18828
rect 3287 18788 3332 18816
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 4540 18816 4568 18856
rect 5712 18853 5724 18887
rect 5758 18884 5770 18887
rect 5902 18884 5908 18896
rect 5758 18856 5908 18884
rect 5758 18853 5770 18856
rect 5712 18847 5770 18853
rect 5902 18844 5908 18856
rect 5960 18844 5966 18896
rect 6932 18884 6960 18924
rect 6003 18856 6960 18884
rect 6003 18816 6031 18856
rect 7098 18844 7104 18896
rect 7156 18884 7162 18896
rect 7156 18856 11284 18884
rect 7156 18844 7162 18856
rect 4540 18788 6031 18816
rect 7193 18819 7251 18825
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7239 18788 8033 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8665 18819 8723 18825
rect 8665 18785 8677 18819
rect 8711 18816 8723 18819
rect 9766 18816 9772 18828
rect 8711 18788 9772 18816
rect 8711 18785 8723 18788
rect 8665 18779 8723 18785
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 10410 18825 10416 18828
rect 10404 18779 10416 18825
rect 10468 18816 10474 18828
rect 10468 18788 10504 18816
rect 10410 18776 10416 18779
rect 10468 18776 10474 18788
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 10836 18788 11192 18816
rect 10836 18776 10842 18788
rect 3510 18748 3516 18760
rect 3471 18720 3516 18748
rect 3510 18708 3516 18720
rect 3568 18708 3574 18760
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 4304 18720 4629 18748
rect 4304 18708 4310 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 5074 18708 5080 18760
rect 5132 18748 5138 18760
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 5132 18720 5457 18748
rect 5132 18708 5138 18720
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 8110 18748 8116 18760
rect 8071 18720 8116 18748
rect 5445 18711 5503 18717
rect 8110 18708 8116 18720
rect 8168 18708 8174 18760
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8260 18720 8305 18748
rect 8260 18708 8266 18720
rect 8478 18708 8484 18760
rect 8536 18748 8542 18760
rect 8849 18751 8907 18757
rect 8849 18748 8861 18751
rect 8536 18720 8861 18748
rect 8536 18708 8542 18720
rect 8849 18717 8861 18720
rect 8895 18717 8907 18751
rect 8849 18711 8907 18717
rect 10042 18708 10048 18760
rect 10100 18748 10106 18760
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 10100 18720 10149 18748
rect 10100 18708 10106 18720
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 3786 18640 3792 18692
rect 3844 18680 3850 18692
rect 4982 18680 4988 18692
rect 3844 18652 4988 18680
rect 3844 18640 3850 18652
rect 4982 18640 4988 18652
rect 5040 18640 5046 18692
rect 9214 18680 9220 18692
rect 6380 18652 9220 18680
rect 6380 18612 6408 18652
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 11164 18680 11192 18788
rect 11256 18748 11284 18856
rect 11974 18844 11980 18896
rect 12032 18884 12038 18896
rect 12069 18887 12127 18893
rect 12069 18884 12081 18887
rect 12032 18856 12081 18884
rect 12032 18844 12038 18856
rect 12069 18853 12081 18856
rect 12115 18853 12127 18887
rect 12069 18847 12127 18853
rect 12158 18844 12164 18896
rect 12216 18884 12222 18896
rect 12805 18887 12863 18893
rect 12805 18884 12817 18887
rect 12216 18856 12817 18884
rect 12216 18844 12222 18856
rect 12805 18853 12817 18856
rect 12851 18853 12863 18887
rect 13280 18884 13308 18924
rect 13354 18912 13360 18964
rect 13412 18952 13418 18964
rect 13633 18955 13691 18961
rect 13633 18952 13645 18955
rect 13412 18924 13645 18952
rect 13412 18912 13418 18924
rect 13633 18921 13645 18924
rect 13679 18921 13691 18955
rect 13633 18915 13691 18921
rect 14093 18955 14151 18961
rect 14093 18921 14105 18955
rect 14139 18952 14151 18955
rect 15289 18955 15347 18961
rect 15289 18952 15301 18955
rect 14139 18924 15301 18952
rect 14139 18921 14151 18924
rect 14093 18915 14151 18921
rect 15289 18921 15301 18924
rect 15335 18921 15347 18955
rect 15289 18915 15347 18921
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18012 18924 18368 18952
rect 18012 18912 18018 18924
rect 13906 18884 13912 18896
rect 13280 18856 13912 18884
rect 12805 18847 12863 18853
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 16574 18884 16580 18896
rect 16535 18856 16580 18884
rect 16574 18844 16580 18856
rect 16632 18844 16638 18896
rect 17034 18844 17040 18896
rect 17092 18884 17098 18896
rect 18340 18893 18368 18924
rect 18325 18887 18383 18893
rect 17092 18856 18184 18884
rect 17092 18844 17098 18856
rect 11790 18816 11796 18828
rect 11751 18788 11796 18816
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 12526 18816 12532 18828
rect 12487 18788 12532 18816
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 13998 18816 14004 18828
rect 13959 18788 14004 18816
rect 13998 18776 14004 18788
rect 14056 18776 14062 18828
rect 14458 18816 14464 18828
rect 14200 18788 14464 18816
rect 14200 18748 14228 18788
rect 14458 18776 14464 18788
rect 14516 18776 14522 18828
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 16301 18819 16359 18825
rect 16301 18785 16313 18819
rect 16347 18816 16359 18819
rect 16666 18816 16672 18828
rect 16347 18788 16672 18816
rect 16347 18785 16359 18788
rect 16301 18779 16359 18785
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 11256 18720 14228 18748
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14550 18748 14556 18760
rect 14323 18720 14556 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15252 18720 15761 18748
rect 15252 18708 15258 18720
rect 15749 18717 15761 18720
rect 15795 18717 15807 18751
rect 15930 18748 15936 18760
rect 15891 18720 15936 18748
rect 15749 18711 15807 18717
rect 15930 18708 15936 18720
rect 15988 18708 15994 18760
rect 16482 18708 16488 18760
rect 16540 18748 16546 18760
rect 17328 18748 17356 18779
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18049 18819 18107 18825
rect 18049 18816 18061 18819
rect 18012 18788 18061 18816
rect 18012 18776 18018 18788
rect 18049 18785 18061 18788
rect 18095 18785 18107 18819
rect 18156 18816 18184 18856
rect 18325 18853 18337 18887
rect 18371 18853 18383 18887
rect 19058 18884 19064 18896
rect 19019 18856 19064 18884
rect 18325 18847 18383 18853
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 18785 18819 18843 18825
rect 18785 18816 18797 18819
rect 18156 18788 18797 18816
rect 18049 18779 18107 18785
rect 18785 18785 18797 18788
rect 18831 18785 18843 18819
rect 18785 18779 18843 18785
rect 16540 18720 17356 18748
rect 17589 18751 17647 18757
rect 16540 18708 16546 18720
rect 17589 18717 17601 18751
rect 17635 18748 17647 18751
rect 18874 18748 18880 18760
rect 17635 18720 18880 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 20622 18680 20628 18692
rect 11164 18652 20628 18680
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 3068 18584 6408 18612
rect 2961 18575 3019 18581
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7653 18615 7711 18621
rect 7653 18612 7665 18615
rect 7156 18584 7665 18612
rect 7156 18572 7162 18584
rect 7653 18581 7665 18584
rect 7699 18581 7711 18615
rect 7653 18575 7711 18581
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 11517 18615 11575 18621
rect 11517 18612 11529 18615
rect 8812 18584 11529 18612
rect 8812 18572 8818 18584
rect 11517 18581 11529 18584
rect 11563 18581 11575 18615
rect 11517 18575 11575 18581
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 5261 18411 5319 18417
rect 5261 18408 5273 18411
rect 2004 18380 5273 18408
rect 2004 18368 2010 18380
rect 5261 18377 5273 18380
rect 5307 18377 5319 18411
rect 5261 18371 5319 18377
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 8168 18380 8217 18408
rect 8168 18368 8174 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 8205 18371 8263 18377
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 9950 18408 9956 18420
rect 8720 18380 9956 18408
rect 8720 18368 8726 18380
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 11425 18411 11483 18417
rect 11425 18408 11437 18411
rect 10376 18380 11437 18408
rect 10376 18368 10382 18380
rect 11425 18377 11437 18380
rect 11471 18377 11483 18411
rect 15194 18408 15200 18420
rect 15155 18380 15200 18408
rect 11425 18371 11483 18377
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 566 18300 572 18352
rect 624 18340 630 18352
rect 2774 18340 2780 18352
rect 624 18312 2780 18340
rect 624 18300 630 18312
rect 2774 18300 2780 18312
rect 2832 18300 2838 18352
rect 5718 18272 5724 18284
rect 1596 18244 3096 18272
rect 5679 18244 5724 18272
rect 1596 18213 1624 18244
rect 1581 18207 1639 18213
rect 1581 18173 1593 18207
rect 1627 18173 1639 18207
rect 2130 18204 2136 18216
rect 2091 18176 2136 18204
rect 1581 18167 1639 18173
rect 2130 18164 2136 18176
rect 2188 18164 2194 18216
rect 2866 18164 2872 18216
rect 2924 18204 2930 18216
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2924 18176 2973 18204
rect 2924 18164 2930 18176
rect 2961 18173 2973 18176
rect 3007 18173 3019 18207
rect 3068 18204 3096 18244
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 5902 18272 5908 18284
rect 5863 18244 5908 18272
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 8754 18272 8760 18284
rect 8715 18244 8760 18272
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 15838 18272 15844 18284
rect 8996 18244 10180 18272
rect 8996 18232 9002 18244
rect 7098 18204 7104 18216
rect 3068 18176 6408 18204
rect 7059 18176 7104 18204
rect 2961 18167 3019 18173
rect 1670 18096 1676 18148
rect 1728 18136 1734 18148
rect 2409 18139 2467 18145
rect 2409 18136 2421 18139
rect 1728 18108 2421 18136
rect 1728 18096 1734 18108
rect 2409 18105 2421 18108
rect 2455 18105 2467 18139
rect 2409 18099 2467 18105
rect 3228 18139 3286 18145
rect 3228 18105 3240 18139
rect 3274 18136 3286 18139
rect 4246 18136 4252 18148
rect 3274 18108 4252 18136
rect 3274 18105 3286 18108
rect 3228 18099 3286 18105
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 5629 18139 5687 18145
rect 5629 18105 5641 18139
rect 5675 18136 5687 18139
rect 6273 18139 6331 18145
rect 6273 18136 6285 18139
rect 5675 18108 6285 18136
rect 5675 18105 5687 18108
rect 5629 18099 5687 18105
rect 6273 18105 6285 18108
rect 6319 18105 6331 18139
rect 6380 18136 6408 18176
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 8665 18207 8723 18213
rect 8665 18173 8677 18207
rect 8711 18204 8723 18207
rect 8846 18204 8852 18216
rect 8711 18176 8852 18204
rect 8711 18173 8723 18176
rect 8665 18167 8723 18173
rect 8846 18164 8852 18176
rect 8904 18164 8910 18216
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 10042 18204 10048 18216
rect 9732 18176 10048 18204
rect 9732 18164 9738 18176
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10152 18204 10180 18244
rect 13096 18244 13308 18272
rect 15799 18244 15844 18272
rect 13096 18204 13124 18244
rect 10152 18176 13124 18204
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18173 13231 18207
rect 13280 18204 13308 18244
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 14366 18204 14372 18216
rect 13280 18176 14372 18204
rect 13173 18167 13231 18173
rect 7377 18139 7435 18145
rect 7377 18136 7389 18139
rect 6380 18108 7389 18136
rect 6273 18099 6331 18105
rect 7377 18105 7389 18108
rect 7423 18105 7435 18139
rect 9950 18136 9956 18148
rect 7377 18099 7435 18105
rect 7668 18108 9956 18136
rect 1762 18068 1768 18080
rect 1723 18040 1768 18068
rect 1762 18028 1768 18040
rect 1820 18028 1826 18080
rect 3510 18028 3516 18080
rect 3568 18068 3574 18080
rect 4341 18071 4399 18077
rect 4341 18068 4353 18071
rect 3568 18040 4353 18068
rect 3568 18028 3574 18040
rect 4341 18037 4353 18040
rect 4387 18037 4399 18071
rect 4341 18031 4399 18037
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 7668 18068 7696 18108
rect 9950 18096 9956 18108
rect 10008 18096 10014 18148
rect 10318 18145 10324 18148
rect 10312 18136 10324 18145
rect 10279 18108 10324 18136
rect 10312 18099 10324 18108
rect 10318 18096 10324 18099
rect 10376 18096 10382 18148
rect 4488 18040 7696 18068
rect 4488 18028 4494 18040
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 8386 18068 8392 18080
rect 7800 18040 8392 18068
rect 7800 18028 7806 18040
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 8570 18068 8576 18080
rect 8483 18040 8576 18068
rect 8570 18028 8576 18040
rect 8628 18068 8634 18080
rect 8754 18068 8760 18080
rect 8628 18040 8760 18068
rect 8628 18028 8634 18040
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 9030 18028 9036 18080
rect 9088 18068 9094 18080
rect 10594 18068 10600 18080
rect 9088 18040 10600 18068
rect 9088 18028 9094 18040
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 13188 18068 13216 18167
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 15010 18204 15016 18216
rect 14971 18176 15016 18204
rect 15010 18164 15016 18176
rect 15068 18204 15074 18216
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 15068 18176 15669 18204
rect 15068 18164 15074 18176
rect 15657 18173 15669 18176
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 13440 18139 13498 18145
rect 13440 18105 13452 18139
rect 13486 18136 13498 18139
rect 15930 18136 15936 18148
rect 13486 18108 15936 18136
rect 13486 18105 13498 18108
rect 13440 18099 13498 18105
rect 15930 18096 15936 18108
rect 15988 18096 15994 18148
rect 16850 18096 16856 18148
rect 16908 18136 16914 18148
rect 22554 18136 22560 18148
rect 16908 18108 22560 18136
rect 16908 18096 16914 18108
rect 22554 18096 22560 18108
rect 22612 18096 22618 18148
rect 13538 18068 13544 18080
rect 13188 18040 13544 18068
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 14550 18068 14556 18080
rect 14511 18040 14556 18068
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 15565 18071 15623 18077
rect 15565 18068 15577 18071
rect 15528 18040 15577 18068
rect 15528 18028 15534 18040
rect 15565 18037 15577 18040
rect 15611 18037 15623 18071
rect 15565 18031 15623 18037
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 20254 18068 20260 18080
rect 19668 18040 20260 18068
rect 19668 18028 19674 18040
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 3050 17864 3056 17876
rect 3011 17836 3056 17864
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3326 17824 3332 17876
rect 3384 17864 3390 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3384 17836 3433 17864
rect 3384 17824 3390 17836
rect 3421 17833 3433 17836
rect 3467 17833 3479 17867
rect 3421 17827 3479 17833
rect 5902 17824 5908 17876
rect 5960 17864 5966 17876
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 5960 17836 6745 17864
rect 5960 17824 5966 17836
rect 6733 17833 6745 17836
rect 6779 17833 6791 17867
rect 6733 17827 6791 17833
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 8619 17836 10149 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 10137 17833 10149 17836
rect 10183 17833 10195 17867
rect 10137 17827 10195 17833
rect 15930 17824 15936 17876
rect 15988 17864 15994 17876
rect 16945 17867 17003 17873
rect 16945 17864 16957 17867
rect 15988 17836 16957 17864
rect 15988 17824 15994 17836
rect 16945 17833 16957 17836
rect 16991 17833 17003 17867
rect 16945 17827 17003 17833
rect 17773 17867 17831 17873
rect 17773 17833 17785 17867
rect 17819 17864 17831 17867
rect 17954 17864 17960 17876
rect 17819 17836 17960 17864
rect 17819 17833 17831 17836
rect 17773 17827 17831 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 7285 17799 7343 17805
rect 7285 17796 7297 17799
rect 1780 17768 7297 17796
rect 1780 17737 1808 17768
rect 7285 17765 7297 17768
rect 7331 17765 7343 17799
rect 7285 17759 7343 17765
rect 9033 17799 9091 17805
rect 9033 17765 9045 17799
rect 9079 17796 9091 17799
rect 9858 17796 9864 17808
rect 9079 17768 9864 17796
rect 9079 17765 9091 17768
rect 9033 17759 9091 17765
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 13808 17799 13866 17805
rect 13808 17765 13820 17799
rect 13854 17796 13866 17799
rect 14550 17796 14556 17808
rect 13854 17768 14556 17796
rect 13854 17765 13866 17768
rect 13808 17759 13866 17765
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17697 2375 17731
rect 2317 17691 2375 17697
rect 2332 17660 2360 17691
rect 2406 17688 2412 17740
rect 2464 17728 2470 17740
rect 2869 17731 2927 17737
rect 2869 17728 2881 17731
rect 2464 17700 2881 17728
rect 2464 17688 2470 17700
rect 2869 17697 2881 17700
rect 2915 17697 2927 17731
rect 2869 17691 2927 17697
rect 5620 17731 5678 17737
rect 5620 17697 5632 17731
rect 5666 17728 5678 17731
rect 6178 17728 6184 17740
rect 5666 17700 6184 17728
rect 5666 17697 5678 17700
rect 5620 17691 5678 17697
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 7006 17728 7012 17740
rect 6967 17700 7012 17728
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 8941 17731 8999 17737
rect 8941 17697 8953 17731
rect 8987 17697 8999 17731
rect 8941 17691 8999 17697
rect 5258 17660 5264 17672
rect 2332 17632 5264 17660
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 2866 17552 2872 17604
rect 2924 17592 2930 17604
rect 5368 17592 5396 17623
rect 6822 17620 6828 17672
rect 6880 17660 6886 17672
rect 8956 17660 8984 17691
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 15838 17737 15844 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9824 17700 10057 17728
rect 9824 17688 9830 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 15832 17728 15844 17737
rect 15799 17700 15844 17728
rect 10045 17691 10103 17697
rect 15832 17691 15844 17700
rect 15838 17688 15844 17691
rect 15896 17688 15902 17740
rect 18141 17731 18199 17737
rect 18141 17697 18153 17731
rect 18187 17728 18199 17731
rect 19058 17728 19064 17740
rect 18187 17700 19064 17728
rect 18187 17697 18199 17700
rect 18141 17691 18199 17697
rect 19058 17688 19064 17700
rect 19116 17688 19122 17740
rect 6880 17632 8984 17660
rect 9217 17663 9275 17669
rect 6880 17620 6886 17632
rect 9217 17629 9229 17663
rect 9263 17660 9275 17663
rect 9858 17660 9864 17672
rect 9263 17632 9864 17660
rect 9263 17629 9275 17632
rect 9217 17623 9275 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 10318 17660 10324 17672
rect 10279 17632 10324 17660
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13354 17660 13360 17672
rect 13127 17632 13360 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13538 17660 13544 17672
rect 13499 17632 13544 17660
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 15562 17660 15568 17672
rect 15523 17632 15568 17660
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18233 17663 18291 17669
rect 18233 17660 18245 17663
rect 18012 17632 18245 17660
rect 18012 17620 18018 17632
rect 18233 17629 18245 17632
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 18506 17660 18512 17672
rect 18463 17632 18512 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 2924 17564 5396 17592
rect 14476 17564 15608 17592
rect 2924 17552 2930 17564
rect 14476 17536 14504 17564
rect 2498 17524 2504 17536
rect 2459 17496 2504 17524
rect 2498 17484 2504 17496
rect 2556 17484 2562 17536
rect 3786 17484 3792 17536
rect 3844 17524 3850 17536
rect 9677 17527 9735 17533
rect 9677 17524 9689 17527
rect 3844 17496 9689 17524
rect 3844 17484 3850 17496
rect 9677 17493 9689 17496
rect 9723 17493 9735 17527
rect 9677 17487 9735 17493
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 12066 17524 12072 17536
rect 11204 17496 12072 17524
rect 11204 17484 11210 17496
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 14458 17484 14464 17536
rect 14516 17484 14522 17536
rect 14550 17484 14556 17536
rect 14608 17524 14614 17536
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 14608 17496 14933 17524
rect 14608 17484 14614 17496
rect 14921 17493 14933 17496
rect 14967 17493 14979 17527
rect 15580 17524 15608 17564
rect 17862 17524 17868 17536
rect 15580 17496 17868 17524
rect 14921 17487 14979 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 5718 17320 5724 17332
rect 5675 17292 5724 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 8478 17320 8484 17332
rect 5828 17292 8484 17320
rect 5258 17212 5264 17264
rect 5316 17252 5322 17264
rect 5828 17252 5856 17292
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 10318 17280 10324 17332
rect 10376 17320 10382 17332
rect 10965 17323 11023 17329
rect 10965 17320 10977 17323
rect 10376 17292 10977 17320
rect 10376 17280 10382 17292
rect 10965 17289 10977 17292
rect 11011 17289 11023 17323
rect 10965 17283 11023 17289
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 12250 17320 12256 17332
rect 11664 17292 12256 17320
rect 11664 17280 11670 17292
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12526 17320 12532 17332
rect 12483 17292 12532 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 13449 17323 13507 17329
rect 13449 17289 13461 17323
rect 13495 17320 13507 17323
rect 13998 17320 14004 17332
rect 13495 17292 14004 17320
rect 13495 17289 13507 17292
rect 13449 17283 13507 17289
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 15381 17323 15439 17329
rect 15381 17289 15393 17323
rect 15427 17320 15439 17323
rect 15654 17320 15660 17332
rect 15427 17292 15660 17320
rect 15427 17289 15439 17292
rect 15381 17283 15439 17289
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 15930 17280 15936 17332
rect 15988 17280 15994 17332
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 18049 17323 18107 17329
rect 18049 17320 18061 17323
rect 18012 17292 18061 17320
rect 18012 17280 18018 17292
rect 18049 17289 18061 17292
rect 18095 17289 18107 17323
rect 18049 17283 18107 17289
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 19794 17320 19800 17332
rect 19392 17292 19800 17320
rect 19392 17280 19398 17292
rect 19794 17280 19800 17292
rect 19852 17280 19858 17332
rect 15948 17252 15976 17280
rect 5316 17224 5856 17252
rect 14108 17224 15976 17252
rect 5316 17212 5322 17224
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 1504 17156 2237 17184
rect 1504 17125 1532 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 2924 17156 3065 17184
rect 2924 17144 2930 17156
rect 3053 17153 3065 17156
rect 3099 17153 3111 17187
rect 6086 17184 6092 17196
rect 6047 17156 6092 17184
rect 3053 17147 3111 17153
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6178 17144 6184 17196
rect 6236 17184 6242 17196
rect 6236 17156 6281 17184
rect 6236 17144 6242 17156
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7340 17156 7389 17184
rect 7340 17144 7346 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 8444 17156 9720 17184
rect 8444 17144 8450 17156
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 1489 17079 1547 17085
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17116 2099 17119
rect 3786 17116 3792 17128
rect 2087 17088 3792 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 3786 17076 3792 17088
rect 3844 17076 3850 17128
rect 7644 17119 7702 17125
rect 7644 17085 7656 17119
rect 7690 17116 7702 17119
rect 8018 17116 8024 17128
rect 7690 17088 8024 17116
rect 7690 17085 7702 17088
rect 7644 17079 7702 17085
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 9490 17116 9496 17128
rect 8904 17088 9496 17116
rect 8904 17076 8910 17088
rect 9490 17076 9496 17088
rect 9548 17116 9554 17128
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 9548 17088 9597 17116
rect 9548 17076 9554 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9692 17116 9720 17156
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 14108 17193 14136 17224
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 11940 17156 13001 17184
rect 11940 17144 11946 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 15838 17184 15844 17196
rect 15712 17156 15844 17184
rect 15712 17144 15718 17156
rect 15838 17144 15844 17156
rect 15896 17184 15902 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15896 17156 15945 17184
rect 15896 17144 15902 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 18598 17184 18604 17196
rect 18559 17156 18604 17184
rect 15933 17147 15991 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 19058 17184 19064 17196
rect 19019 17156 19064 17184
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 9692 17088 13216 17116
rect 9585 17079 9643 17085
rect 3320 17051 3378 17057
rect 3320 17017 3332 17051
rect 3366 17048 3378 17051
rect 3510 17048 3516 17060
rect 3366 17020 3516 17048
rect 3366 17017 3378 17020
rect 3320 17011 3378 17017
rect 3510 17008 3516 17020
rect 3568 17008 3574 17060
rect 3878 17008 3884 17060
rect 3936 17048 3942 17060
rect 9858 17057 9864 17060
rect 9852 17048 9864 17057
rect 3936 17020 9720 17048
rect 9771 17020 9864 17048
rect 3936 17008 3942 17020
rect 9692 16992 9720 17020
rect 9852 17011 9864 17020
rect 9916 17048 9922 17060
rect 10226 17048 10232 17060
rect 9916 17020 10232 17048
rect 9858 17008 9864 17011
rect 9916 17008 9922 17020
rect 10226 17008 10232 17020
rect 10284 17008 10290 17060
rect 13188 17048 13216 17088
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 13817 17119 13875 17125
rect 13817 17116 13829 17119
rect 13412 17088 13829 17116
rect 13412 17076 13418 17088
rect 13817 17085 13829 17088
rect 13863 17085 13875 17119
rect 13817 17079 13875 17085
rect 15749 17119 15807 17125
rect 15749 17085 15761 17119
rect 15795 17116 15807 17119
rect 16206 17116 16212 17128
rect 15795 17088 16212 17116
rect 15795 17085 15807 17088
rect 15749 17079 15807 17085
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 17920 17088 18521 17116
rect 17920 17076 17926 17088
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 21634 17116 21640 17128
rect 20956 17088 21640 17116
rect 20956 17076 20962 17088
rect 21634 17076 21640 17088
rect 21692 17076 21698 17128
rect 13909 17051 13967 17057
rect 13909 17048 13921 17051
rect 13188 17020 13921 17048
rect 13909 17017 13921 17020
rect 13955 17017 13967 17051
rect 18414 17048 18420 17060
rect 18375 17020 18420 17048
rect 13909 17011 13967 17017
rect 18414 17008 18420 17020
rect 18472 17048 18478 17060
rect 18877 17051 18935 17057
rect 18877 17048 18889 17051
rect 18472 17020 18889 17048
rect 18472 17008 18478 17020
rect 18877 17017 18889 17020
rect 18923 17017 18935 17051
rect 18877 17011 18935 17017
rect 20714 17008 20720 17060
rect 20772 17048 20778 17060
rect 20990 17048 20996 17060
rect 20772 17020 20996 17048
rect 20772 17008 20778 17020
rect 20990 17008 20996 17020
rect 21048 17008 21054 17060
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 4212 16952 4445 16980
rect 4212 16940 4218 16952
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4433 16943 4491 16949
rect 5902 16940 5908 16992
rect 5960 16980 5966 16992
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 5960 16952 6009 16980
rect 5960 16940 5966 16952
rect 5997 16949 6009 16952
rect 6043 16980 6055 16983
rect 6822 16980 6828 16992
rect 6043 16952 6828 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8260 16952 8769 16980
rect 8260 16940 8266 16952
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 8757 16943 8815 16949
rect 9674 16940 9680 16992
rect 9732 16940 9738 16992
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 12952 16952 12997 16980
rect 12952 16940 12958 16952
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 15838 16980 15844 16992
rect 13320 16952 15844 16980
rect 13320 16940 13326 16952
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 16298 16940 16304 16992
rect 16356 16980 16362 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16356 16952 16957 16980
rect 16356 16940 16362 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2056 16748 2881 16776
rect 1486 16640 1492 16652
rect 1447 16612 1492 16640
rect 1486 16600 1492 16612
rect 1544 16600 1550 16652
rect 2056 16649 2084 16748
rect 2869 16745 2881 16748
rect 2915 16745 2927 16779
rect 2869 16739 2927 16745
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 6236 16748 6377 16776
rect 6236 16736 6242 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 9766 16776 9772 16788
rect 9727 16748 9772 16776
rect 6365 16739 6423 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13817 16779 13875 16785
rect 13817 16776 13829 16779
rect 12952 16748 13829 16776
rect 12952 16736 12958 16748
rect 13817 16745 13829 16748
rect 13863 16745 13875 16779
rect 13817 16739 13875 16745
rect 15933 16779 15991 16785
rect 15933 16745 15945 16779
rect 15979 16745 15991 16779
rect 16298 16776 16304 16788
rect 16259 16748 16304 16776
rect 15933 16739 15991 16745
rect 2317 16711 2375 16717
rect 2317 16677 2329 16711
rect 2363 16708 2375 16711
rect 2406 16708 2412 16720
rect 2363 16680 2412 16708
rect 2363 16677 2375 16680
rect 2317 16671 2375 16677
rect 2406 16668 2412 16680
rect 2464 16668 2470 16720
rect 7098 16668 7104 16720
rect 7156 16708 7162 16720
rect 10772 16711 10830 16717
rect 7156 16680 8984 16708
rect 7156 16668 7162 16680
rect 2051 16643 2109 16649
rect 2051 16609 2063 16643
rect 2097 16609 2109 16643
rect 3234 16640 3240 16652
rect 3195 16612 3240 16640
rect 2051 16603 2109 16609
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16640 3387 16643
rect 4246 16640 4252 16652
rect 3375 16612 4252 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 5252 16643 5310 16649
rect 5252 16609 5264 16643
rect 5298 16640 5310 16643
rect 5810 16640 5816 16652
rect 5298 16612 5816 16640
rect 5298 16609 5310 16612
rect 5252 16603 5310 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 7190 16640 7196 16652
rect 6687 16612 7196 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7368 16643 7426 16649
rect 7368 16609 7380 16643
rect 7414 16640 7426 16643
rect 8202 16640 8208 16652
rect 7414 16612 8208 16640
rect 7414 16609 7426 16612
rect 7368 16603 7426 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8956 16649 8984 16680
rect 10772 16677 10784 16711
rect 10818 16708 10830 16711
rect 12986 16708 12992 16720
rect 10818 16680 12992 16708
rect 10818 16677 10830 16680
rect 10772 16671 10830 16677
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 15948 16708 15976 16739
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 18325 16779 18383 16785
rect 18325 16745 18337 16779
rect 18371 16745 18383 16779
rect 18325 16739 18383 16745
rect 16758 16708 16764 16720
rect 15948 16680 16764 16708
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 18340 16708 18368 16739
rect 18506 16736 18512 16788
rect 18564 16776 18570 16788
rect 19981 16779 20039 16785
rect 19981 16776 19993 16779
rect 18564 16748 19993 16776
rect 18564 16736 18570 16748
rect 19981 16745 19993 16748
rect 20027 16745 20039 16779
rect 19981 16739 20039 16745
rect 18598 16708 18604 16720
rect 18340 16680 18604 16708
rect 18598 16668 18604 16680
rect 18656 16708 18662 16720
rect 18846 16711 18904 16717
rect 18846 16708 18858 16711
rect 18656 16680 18858 16708
rect 18656 16668 18662 16680
rect 18846 16677 18858 16680
rect 18892 16677 18904 16711
rect 18846 16671 18904 16677
rect 12434 16649 12440 16652
rect 8941 16643 8999 16649
rect 8941 16609 8953 16643
rect 8987 16609 8999 16643
rect 10505 16643 10563 16649
rect 10505 16640 10517 16643
rect 8941 16603 8999 16609
rect 9048 16612 10517 16640
rect 3513 16575 3571 16581
rect 3513 16541 3525 16575
rect 3559 16572 3571 16575
rect 3970 16572 3976 16584
rect 3559 16544 3976 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 9048 16572 9076 16612
rect 10505 16609 10517 16612
rect 10551 16609 10563 16643
rect 12161 16643 12219 16649
rect 12161 16640 12173 16643
rect 10505 16603 10563 16609
rect 11532 16612 12173 16640
rect 7101 16535 7159 16541
rect 8864 16544 9076 16572
rect 1670 16504 1676 16516
rect 1631 16476 1676 16504
rect 1670 16464 1676 16476
rect 1728 16464 1734 16516
rect 2866 16464 2872 16516
rect 2924 16504 2930 16516
rect 5000 16504 5028 16535
rect 2924 16476 5028 16504
rect 2924 16464 2930 16476
rect 7116 16436 7144 16535
rect 8864 16516 8892 16544
rect 8757 16507 8815 16513
rect 8757 16504 8769 16507
rect 8220 16476 8769 16504
rect 7282 16436 7288 16448
rect 7116 16408 7288 16436
rect 7282 16396 7288 16408
rect 7340 16436 7346 16448
rect 8220 16436 8248 16476
rect 8757 16473 8769 16476
rect 8803 16504 8815 16507
rect 8846 16504 8852 16516
rect 8803 16476 8852 16504
rect 8803 16473 8815 16476
rect 8757 16467 8815 16473
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 7340 16408 8248 16436
rect 7340 16396 7346 16408
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 8481 16439 8539 16445
rect 8481 16436 8493 16439
rect 8352 16408 8493 16436
rect 8352 16396 8358 16408
rect 8481 16405 8493 16408
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 10410 16396 10416 16448
rect 10468 16436 10474 16448
rect 11532 16436 11560 16612
rect 12161 16609 12173 16612
rect 12207 16609 12219 16643
rect 12428 16640 12440 16649
rect 12395 16612 12440 16640
rect 12161 16603 12219 16609
rect 12428 16603 12440 16612
rect 11882 16436 11888 16448
rect 10468 16408 11560 16436
rect 11843 16408 11888 16436
rect 10468 16396 10474 16408
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12176 16436 12204 16603
rect 12434 16600 12440 16603
rect 12492 16600 12498 16652
rect 12894 16600 12900 16652
rect 12952 16640 12958 16652
rect 13538 16640 13544 16652
rect 12952 16612 13544 16640
rect 12952 16600 12958 16612
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 14182 16640 14188 16652
rect 14143 16612 14188 16640
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 17218 16649 17224 16652
rect 17212 16640 17224 16649
rect 16592 16612 17224 16640
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 16390 16572 16396 16584
rect 16351 16544 16396 16572
rect 14369 16535 14427 16541
rect 14384 16504 14412 16535
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 16592 16581 16620 16612
rect 17212 16603 17224 16612
rect 17218 16600 17224 16603
rect 17276 16600 17282 16652
rect 17972 16612 18644 16640
rect 16577 16575 16635 16581
rect 16577 16541 16589 16575
rect 16623 16541 16635 16575
rect 16577 16535 16635 16541
rect 16945 16575 17003 16581
rect 16945 16541 16957 16575
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 13556 16476 14412 16504
rect 12894 16436 12900 16448
rect 12176 16408 12900 16436
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 13556 16445 13584 16476
rect 15562 16464 15568 16516
rect 15620 16504 15626 16516
rect 16960 16504 16988 16535
rect 17972 16504 18000 16612
rect 18616 16581 18644 16612
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 15620 16476 16988 16504
rect 15620 16464 15626 16476
rect 13541 16439 13599 16445
rect 13541 16436 13553 16439
rect 13136 16408 13553 16436
rect 13136 16396 13142 16408
rect 13541 16405 13553 16408
rect 13587 16405 13599 16439
rect 16960 16436 16988 16476
rect 17880 16476 18000 16504
rect 17880 16436 17908 16476
rect 16960 16408 17908 16436
rect 13541 16399 13599 16405
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 4246 16232 4252 16244
rect 1872 16204 3547 16232
rect 4207 16204 4252 16232
rect 1872 16037 1900 16204
rect 3519 16164 3547 16204
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 5261 16235 5319 16241
rect 5261 16232 5273 16235
rect 4347 16204 5273 16232
rect 4347 16164 4375 16204
rect 5261 16201 5273 16204
rect 5307 16201 5319 16235
rect 5261 16195 5319 16201
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 10226 16232 10232 16244
rect 7432 16204 9996 16232
rect 10187 16204 10232 16232
rect 7432 16192 7438 16204
rect 3519 16136 4375 16164
rect 4890 16124 4896 16176
rect 4948 16164 4954 16176
rect 8662 16164 8668 16176
rect 4948 16136 8668 16164
rect 4948 16124 4954 16136
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 4706 16096 4712 16108
rect 4667 16068 4712 16096
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16065 4859 16099
rect 5810 16096 5816 16108
rect 5771 16068 5816 16096
rect 4801 16059 4859 16065
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 15997 1915 16031
rect 1857 15991 1915 15997
rect 2593 16031 2651 16037
rect 2593 15997 2605 16031
rect 2639 16028 2651 16031
rect 2860 16031 2918 16037
rect 2639 16000 2820 16028
rect 2639 15997 2651 16000
rect 2593 15991 2651 15997
rect 2792 15972 2820 16000
rect 2860 15997 2872 16031
rect 2906 16028 2918 16031
rect 4154 16028 4160 16040
rect 2906 16000 4160 16028
rect 2906 15997 2918 16000
rect 2860 15991 2918 15997
rect 4154 15988 4160 16000
rect 4212 16028 4218 16040
rect 4816 16028 4844 16059
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7800 16068 7941 16096
rect 7800 16056 7806 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 8113 16099 8171 16105
rect 8113 16065 8125 16099
rect 8159 16096 8171 16099
rect 8202 16096 8208 16108
rect 8159 16068 8208 16096
rect 8159 16065 8171 16068
rect 8113 16059 8171 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8846 16096 8852 16108
rect 8807 16068 8852 16096
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 4212 16000 4844 16028
rect 6457 16031 6515 16037
rect 4212 15988 4218 16000
rect 6457 15997 6469 16031
rect 6503 16028 6515 16031
rect 7098 16028 7104 16040
rect 6503 16000 7104 16028
rect 6503 15997 6515 16000
rect 6457 15991 6515 15997
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 2774 15920 2780 15972
rect 2832 15920 2838 15972
rect 7837 15963 7895 15969
rect 7837 15960 7849 15963
rect 5184 15932 7849 15960
rect 5184 15904 5212 15932
rect 7837 15929 7849 15932
rect 7883 15929 7895 15963
rect 7837 15923 7895 15929
rect 9116 15963 9174 15969
rect 9116 15929 9128 15963
rect 9162 15960 9174 15963
rect 9858 15960 9864 15972
rect 9162 15932 9864 15960
rect 9162 15929 9174 15932
rect 9116 15923 9174 15929
rect 9858 15920 9864 15932
rect 9916 15920 9922 15972
rect 9968 15960 9996 16204
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12802 16232 12808 16244
rect 12483 16204 12808 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 13909 16235 13967 16241
rect 13909 16201 13921 16235
rect 13955 16232 13967 16235
rect 14182 16232 14188 16244
rect 13955 16204 14188 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 17276 16204 17417 16232
rect 17276 16192 17282 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 15010 16164 15016 16176
rect 12452 16136 15016 16164
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 10505 16031 10563 16037
rect 10505 16028 10517 16031
rect 10468 16000 10517 16028
rect 10468 15988 10474 16000
rect 10505 15997 10517 16000
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 10772 16031 10830 16037
rect 10772 15997 10784 16031
rect 10818 16028 10830 16031
rect 11882 16028 11888 16040
rect 10818 16000 11888 16028
rect 10818 15997 10830 16000
rect 10772 15991 10830 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 12452 16028 12480 16136
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 12986 16096 12992 16108
rect 12947 16068 12992 16096
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 14366 16096 14372 16108
rect 14327 16068 14372 16096
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 15562 16056 15568 16108
rect 15620 16096 15626 16108
rect 16022 16096 16028 16108
rect 15620 16068 16028 16096
rect 15620 16056 15626 16068
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 11992 16000 12480 16028
rect 12544 16000 12909 16028
rect 11992 15960 12020 16000
rect 12544 15960 12572 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 14277 16031 14335 16037
rect 14277 15997 14289 16031
rect 14323 16028 14335 16031
rect 14458 16028 14464 16040
rect 14323 16000 14464 16028
rect 14323 15997 14335 16000
rect 14277 15991 14335 15997
rect 14458 15988 14464 16000
rect 14516 16028 14522 16040
rect 15102 16028 15108 16040
rect 14516 16000 15108 16028
rect 14516 15988 14522 16000
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 9968 15932 12020 15960
rect 12452 15932 12572 15960
rect 12805 15963 12863 15969
rect 3970 15892 3976 15904
rect 3931 15864 3976 15892
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 5166 15892 5172 15904
rect 4663 15864 5172 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 5776 15864 5821 15892
rect 5776 15852 5782 15864
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 6273 15895 6331 15901
rect 6273 15892 6285 15895
rect 6052 15864 6285 15892
rect 6052 15852 6058 15864
rect 6273 15861 6285 15864
rect 6319 15861 6331 15895
rect 6273 15855 6331 15861
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 7469 15895 7527 15901
rect 7469 15892 7481 15895
rect 7340 15864 7481 15892
rect 7340 15852 7346 15864
rect 7469 15861 7481 15864
rect 7515 15861 7527 15895
rect 7469 15855 7527 15861
rect 11606 15852 11612 15904
rect 11664 15892 11670 15904
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11664 15864 11897 15892
rect 11664 15852 11670 15864
rect 11885 15861 11897 15864
rect 11931 15861 11943 15895
rect 11885 15855 11943 15861
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 12452 15892 12480 15932
rect 12805 15929 12817 15963
rect 12851 15960 12863 15963
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 12851 15932 13461 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 13449 15929 13461 15932
rect 13495 15929 13507 15963
rect 16114 15960 16120 15972
rect 13449 15923 13507 15929
rect 13556 15932 16120 15960
rect 12216 15864 12480 15892
rect 12216 15852 12222 15864
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 13556 15892 13584 15932
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 16292 15963 16350 15969
rect 16292 15929 16304 15963
rect 16338 15960 16350 15963
rect 16574 15960 16580 15972
rect 16338 15932 16580 15960
rect 16338 15929 16350 15932
rect 16292 15923 16350 15929
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 12584 15864 13584 15892
rect 12584 15852 12590 15864
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 16850 15892 16856 15904
rect 13688 15864 16856 15892
rect 13688 15852 13694 15864
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 3145 15691 3203 15697
rect 3145 15657 3157 15691
rect 3191 15688 3203 15691
rect 3234 15688 3240 15700
rect 3191 15660 3240 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 6365 15691 6423 15697
rect 6365 15688 6377 15691
rect 5684 15660 6377 15688
rect 5684 15648 5690 15660
rect 6365 15657 6377 15660
rect 6411 15657 6423 15691
rect 6365 15651 6423 15657
rect 6825 15691 6883 15697
rect 6825 15657 6837 15691
rect 6871 15688 6883 15691
rect 7006 15688 7012 15700
rect 6871 15660 7012 15688
rect 6871 15657 6883 15660
rect 6825 15651 6883 15657
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 8941 15691 8999 15697
rect 8941 15657 8953 15691
rect 8987 15688 8999 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 8987 15660 9689 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 10134 15688 10140 15700
rect 10095 15660 10140 15688
rect 9677 15651 9735 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 12158 15688 12164 15700
rect 12119 15660 12164 15688
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 12621 15691 12679 15697
rect 12621 15657 12633 15691
rect 12667 15688 12679 15691
rect 13538 15688 13544 15700
rect 12667 15660 13544 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 14274 15688 14280 15700
rect 13679 15660 14280 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 14645 15691 14703 15697
rect 14645 15657 14657 15691
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 15841 15691 15899 15697
rect 15841 15657 15853 15691
rect 15887 15688 15899 15691
rect 16390 15688 16396 15700
rect 15887 15660 16396 15688
rect 15887 15657 15899 15660
rect 15841 15651 15899 15657
rect 1486 15580 1492 15632
rect 1544 15620 1550 15632
rect 2225 15623 2283 15629
rect 2225 15620 2237 15623
rect 1544 15592 2237 15620
rect 1544 15580 1550 15592
rect 2225 15589 2237 15592
rect 2271 15589 2283 15623
rect 5994 15620 6000 15632
rect 2225 15583 2283 15589
rect 4724 15592 6000 15620
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 1959 15555 2017 15561
rect 1959 15521 1971 15555
rect 2005 15521 2017 15555
rect 1959 15515 2017 15521
rect 1964 15348 1992 15515
rect 3510 15444 3516 15496
rect 3568 15484 3574 15496
rect 4724 15493 4752 15592
rect 5994 15580 6000 15592
rect 6052 15580 6058 15632
rect 7190 15620 7196 15632
rect 7151 15592 7196 15620
rect 7190 15580 7196 15592
rect 7248 15580 7254 15632
rect 10045 15623 10103 15629
rect 10045 15620 10057 15623
rect 7300 15592 10057 15620
rect 4976 15555 5034 15561
rect 4976 15521 4988 15555
rect 5022 15552 5034 15555
rect 6270 15552 6276 15564
rect 5022 15524 6276 15552
rect 5022 15521 5034 15524
rect 4976 15515 5034 15521
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 7300 15552 7328 15592
rect 10045 15589 10057 15592
rect 10091 15589 10103 15623
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 10045 15583 10103 15589
rect 10244 15592 11529 15620
rect 6420 15524 7328 15552
rect 8021 15555 8079 15561
rect 6420 15512 6426 15524
rect 8021 15521 8033 15555
rect 8067 15552 8079 15555
rect 8849 15555 8907 15561
rect 8849 15552 8861 15555
rect 8067 15524 8861 15552
rect 8067 15521 8079 15524
rect 8021 15515 8079 15521
rect 8849 15521 8861 15524
rect 8895 15521 8907 15555
rect 8849 15515 8907 15521
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10244 15552 10272 15592
rect 11517 15589 11529 15592
rect 11563 15620 11575 15623
rect 13262 15620 13268 15632
rect 11563 15592 13268 15620
rect 11563 15589 11575 15592
rect 11517 15583 11575 15589
rect 13262 15580 13268 15592
rect 13320 15580 13326 15632
rect 14660 15620 14688 15651
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 13372 15592 17080 15620
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 10008 15524 10272 15552
rect 10336 15524 11437 15552
rect 10008 15512 10014 15524
rect 4709 15487 4767 15493
rect 4709 15484 4721 15487
rect 3568 15456 4721 15484
rect 3568 15444 3574 15456
rect 4709 15453 4721 15456
rect 4755 15453 4767 15487
rect 4709 15447 4767 15453
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 8294 15484 8300 15496
rect 7515 15456 8300 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9858 15484 9864 15496
rect 9171 15456 9864 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10226 15484 10232 15496
rect 10187 15456 10232 15484
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 8481 15419 8539 15425
rect 8481 15416 8493 15419
rect 5644 15388 8493 15416
rect 5644 15348 5672 15388
rect 8481 15385 8493 15388
rect 8527 15385 8539 15419
rect 8481 15379 8539 15385
rect 1964 15320 5672 15348
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 5868 15320 6101 15348
rect 5868 15308 5874 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 7466 15308 7472 15360
rect 7524 15348 7530 15360
rect 10336 15348 10364 15524
rect 11425 15521 11437 15524
rect 11471 15552 11483 15555
rect 12342 15552 12348 15564
rect 11471 15524 12348 15552
rect 11471 15521 11483 15524
rect 11425 15515 11483 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 12526 15552 12532 15564
rect 12487 15524 12532 15552
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 13372 15561 13400 15592
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14001 15555 14059 15561
rect 14001 15552 14013 15555
rect 13872 15524 14013 15552
rect 13872 15512 13878 15524
rect 14001 15521 14013 15524
rect 14047 15521 14059 15555
rect 14001 15515 14059 15521
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 14516 15524 14841 15552
rect 14516 15512 14522 15524
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 15010 15512 15016 15564
rect 15068 15552 15074 15564
rect 17052 15561 17080 15592
rect 16209 15555 16267 15561
rect 16209 15552 16221 15555
rect 15068 15524 16221 15552
rect 15068 15512 15074 15524
rect 16209 15521 16221 15524
rect 16255 15521 16267 15555
rect 16209 15515 16267 15521
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 11606 15484 11612 15496
rect 11567 15456 11612 15484
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12805 15487 12863 15493
rect 12805 15484 12817 15487
rect 12492 15456 12817 15484
rect 12492 15444 12498 15456
rect 12805 15453 12817 15456
rect 12851 15484 12863 15487
rect 12851 15456 13768 15484
rect 12851 15453 12863 15456
rect 12805 15447 12863 15453
rect 13740 15416 13768 15456
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13964 15456 14105 15484
rect 13964 15444 13970 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 14550 15484 14556 15496
rect 14323 15456 14556 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 14292 15416 14320 15447
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 16301 15487 16359 15493
rect 16301 15484 16313 15487
rect 15896 15456 16313 15484
rect 15896 15444 15902 15456
rect 16301 15453 16313 15456
rect 16347 15453 16359 15487
rect 16301 15447 16359 15453
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15484 16543 15487
rect 16574 15484 16580 15496
rect 16531 15456 16580 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 16574 15444 16580 15456
rect 16632 15484 16638 15496
rect 17402 15484 17408 15496
rect 16632 15456 17408 15484
rect 16632 15444 16638 15456
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 13740 15388 14320 15416
rect 16022 15376 16028 15428
rect 16080 15416 16086 15428
rect 16853 15419 16911 15425
rect 16853 15416 16865 15419
rect 16080 15388 16865 15416
rect 16080 15376 16086 15388
rect 16853 15385 16865 15388
rect 16899 15385 16911 15419
rect 16853 15379 16911 15385
rect 7524 15320 10364 15348
rect 11057 15351 11115 15357
rect 7524 15308 7530 15320
rect 11057 15317 11069 15351
rect 11103 15348 11115 15351
rect 11146 15348 11152 15360
rect 11103 15320 11152 15348
rect 11103 15317 11115 15320
rect 11057 15311 11115 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 13078 15308 13084 15360
rect 13136 15348 13142 15360
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 13136 15320 13185 15348
rect 13136 15308 13142 15320
rect 13173 15317 13185 15320
rect 13219 15317 13231 15351
rect 13173 15311 13231 15317
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 5074 15144 5080 15156
rect 1964 15116 5080 15144
rect 1964 14949 1992 15116
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 5629 15147 5687 15153
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 5718 15144 5724 15156
rect 5675 15116 5724 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 8846 15144 8852 15156
rect 8496 15116 8852 15144
rect 5994 15036 6000 15088
rect 6052 15076 6058 15088
rect 6052 15048 6868 15076
rect 6052 15036 6058 15048
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 6270 15008 6276 15020
rect 2832 14980 2877 15008
rect 6231 14980 6276 15008
rect 2832 14968 2838 14980
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 6840 15017 6868 15048
rect 8496 15017 8524 15116
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9858 15144 9864 15156
rect 9819 15116 9864 15144
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 13081 15147 13139 15153
rect 13081 15113 13093 15147
rect 13127 15144 13139 15147
rect 13170 15144 13176 15156
rect 13127 15116 13176 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 15654 15144 15660 15156
rect 15615 15116 15660 15144
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 17402 15144 17408 15156
rect 17363 15116 17408 15144
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 8481 15011 8539 15017
rect 8481 14977 8493 15011
rect 8527 14977 8539 15011
rect 11606 15008 11612 15020
rect 11567 14980 11612 15008
rect 8481 14971 8539 14977
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 16022 15008 16028 15020
rect 13771 14980 14412 15008
rect 15983 14980 16028 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14909 2007 14943
rect 1949 14903 2007 14909
rect 1412 14872 1440 14903
rect 2225 14875 2283 14881
rect 2225 14872 2237 14875
rect 1412 14844 2237 14872
rect 2225 14841 2237 14844
rect 2271 14841 2283 14875
rect 2792 14872 2820 14968
rect 3044 14943 3102 14949
rect 3044 14909 3056 14943
rect 3090 14940 3102 14943
rect 3970 14940 3976 14952
rect 3090 14912 3976 14940
rect 3090 14909 3102 14912
rect 3044 14903 3102 14909
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6546 14940 6552 14952
rect 6135 14912 6552 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 7092 14943 7150 14949
rect 7092 14909 7104 14943
rect 7138 14940 7150 14943
rect 8294 14940 8300 14952
rect 7138 14912 8300 14940
rect 7138 14909 7150 14912
rect 7092 14903 7150 14909
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 8748 14943 8806 14949
rect 8748 14909 8760 14943
rect 8794 14940 8806 14943
rect 9674 14940 9680 14952
rect 8794 14912 9680 14940
rect 8794 14909 8806 14912
rect 8748 14903 8806 14909
rect 9674 14900 9680 14912
rect 9732 14940 9738 14952
rect 10226 14940 10232 14952
rect 9732 14912 10232 14940
rect 9732 14900 9738 14912
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11112 14912 11529 14940
rect 11112 14900 11118 14912
rect 11517 14909 11529 14912
rect 11563 14940 11575 14943
rect 12342 14940 12348 14952
rect 11563 14912 12348 14940
rect 11563 14909 11575 14912
rect 11517 14903 11575 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14384 14940 14412 14980
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 14550 14949 14556 14952
rect 14533 14943 14556 14949
rect 14533 14940 14545 14943
rect 14384 14912 14545 14940
rect 14277 14903 14335 14909
rect 14533 14909 14545 14912
rect 14608 14940 14614 14952
rect 16040 14940 16068 14968
rect 18046 14940 18052 14952
rect 14608 14912 14681 14940
rect 16040 14912 18052 14940
rect 14533 14903 14556 14909
rect 2792 14844 3096 14872
rect 2225 14835 2283 14841
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 2958 14804 2964 14816
rect 1627 14776 2964 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 2958 14764 2964 14776
rect 3016 14764 3022 14816
rect 3068 14804 3096 14844
rect 5810 14832 5816 14884
rect 5868 14872 5874 14884
rect 5997 14875 6055 14881
rect 5997 14872 6009 14875
rect 5868 14844 6009 14872
rect 5868 14832 5874 14844
rect 5997 14841 6009 14844
rect 6043 14872 6055 14875
rect 6362 14872 6368 14884
rect 6043 14844 6368 14872
rect 6043 14841 6055 14844
rect 5997 14835 6055 14841
rect 6362 14832 6368 14844
rect 6420 14832 6426 14884
rect 11425 14875 11483 14881
rect 11425 14841 11437 14875
rect 11471 14872 11483 14875
rect 14292 14872 14320 14903
rect 14550 14900 14556 14903
rect 14608 14900 14614 14912
rect 16040 14872 16068 14912
rect 18046 14900 18052 14912
rect 18104 14940 18110 14952
rect 18141 14943 18199 14949
rect 18141 14940 18153 14943
rect 18104 14912 18153 14940
rect 18104 14900 18110 14912
rect 18141 14909 18153 14912
rect 18187 14909 18199 14943
rect 18141 14903 18199 14909
rect 11471 14844 14044 14872
rect 14292 14844 16068 14872
rect 16292 14875 16350 14881
rect 11471 14841 11483 14844
rect 11425 14835 11483 14841
rect 3510 14804 3516 14816
rect 3068 14776 3516 14804
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 4154 14804 4160 14816
rect 4115 14776 4160 14804
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 7524 14776 8217 14804
rect 7524 14764 7530 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 11054 14804 11060 14816
rect 11015 14776 11060 14804
rect 8205 14767 8263 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 13446 14804 13452 14816
rect 13407 14776 13452 14804
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 14016 14804 14044 14844
rect 16292 14841 16304 14875
rect 16338 14872 16350 14875
rect 16942 14872 16948 14884
rect 16338 14844 16948 14872
rect 16338 14841 16350 14844
rect 16292 14835 16350 14841
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 18408 14875 18466 14881
rect 18408 14841 18420 14875
rect 18454 14872 18466 14875
rect 18506 14872 18512 14884
rect 18454 14844 18512 14872
rect 18454 14841 18466 14844
rect 18408 14835 18466 14841
rect 18506 14832 18512 14844
rect 18564 14832 18570 14884
rect 15562 14804 15568 14816
rect 13596 14776 13641 14804
rect 14016 14776 15568 14804
rect 13596 14764 13602 14776
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 19518 14804 19524 14816
rect 19479 14776 19524 14804
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1762 14600 1768 14612
rect 1723 14572 1768 14600
rect 1762 14560 1768 14572
rect 1820 14560 1826 14612
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 4798 14600 4804 14612
rect 4571 14572 4804 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7156 14572 7665 14600
rect 7156 14560 7162 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 14550 14600 14556 14612
rect 14511 14572 14556 14600
rect 7653 14563 7711 14569
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 17034 14600 17040 14612
rect 16995 14572 17040 14600
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 1394 14492 1400 14544
rect 1452 14532 1458 14544
rect 2409 14535 2467 14541
rect 2409 14532 2421 14535
rect 1452 14504 2421 14532
rect 1452 14492 1458 14504
rect 2409 14501 2421 14504
rect 2455 14501 2467 14535
rect 2409 14495 2467 14501
rect 4433 14535 4491 14541
rect 4433 14501 4445 14535
rect 4479 14532 4491 14535
rect 7006 14532 7012 14544
rect 4479 14504 7012 14532
rect 4479 14501 4491 14504
rect 4433 14495 4491 14501
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 10680 14535 10738 14541
rect 10680 14501 10692 14535
rect 10726 14532 10738 14535
rect 11606 14532 11612 14544
rect 10726 14504 11612 14532
rect 10726 14501 10738 14504
rect 10680 14495 10738 14501
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 17405 14535 17463 14541
rect 17405 14501 17417 14535
rect 17451 14532 17463 14535
rect 17954 14532 17960 14544
rect 17451 14504 17960 14532
rect 17451 14501 17463 14504
rect 17405 14495 17463 14501
rect 17954 14492 17960 14504
rect 18012 14492 18018 14544
rect 18316 14535 18374 14541
rect 18316 14501 18328 14535
rect 18362 14532 18374 14535
rect 18690 14532 18696 14544
rect 18362 14504 18696 14532
rect 18362 14501 18374 14504
rect 18316 14495 18374 14501
rect 18690 14492 18696 14504
rect 18748 14532 18754 14544
rect 19518 14532 19524 14544
rect 18748 14504 19524 14532
rect 18748 14492 18754 14504
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 1946 14464 1952 14476
rect 1627 14436 1952 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 2498 14464 2504 14476
rect 2179 14436 2504 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 5994 14464 6000 14476
rect 5955 14436 6000 14464
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6264 14467 6322 14473
rect 6264 14433 6276 14467
rect 6310 14464 6322 14467
rect 7466 14464 7472 14476
rect 6310 14436 7472 14464
rect 6310 14433 6322 14436
rect 6264 14427 6322 14433
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 7837 14467 7895 14473
rect 7837 14464 7849 14467
rect 7800 14436 7849 14464
rect 7800 14424 7806 14436
rect 7837 14433 7849 14436
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 10226 14464 10232 14476
rect 8352 14436 10232 14464
rect 8352 14424 8358 14436
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10410 14464 10416 14476
rect 10371 14436 10416 14464
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 13078 14424 13084 14476
rect 13136 14464 13142 14476
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 13136 14436 13185 14464
rect 13136 14424 13142 14436
rect 13173 14433 13185 14436
rect 13219 14433 13231 14467
rect 13173 14427 13231 14433
rect 13262 14424 13268 14476
rect 13320 14464 13326 14476
rect 13429 14467 13487 14473
rect 13429 14464 13441 14467
rect 13320 14436 13441 14464
rect 13320 14424 13326 14436
rect 13429 14433 13441 14436
rect 13475 14433 13487 14467
rect 13429 14427 13487 14433
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 15102 14464 15108 14476
rect 14424 14436 15108 14464
rect 14424 14424 14430 14436
rect 15102 14424 15108 14436
rect 15160 14464 15166 14476
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15160 14436 15761 14464
rect 15160 14424 15166 14436
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 18046 14464 18052 14476
rect 18007 14436 18052 14464
rect 15749 14427 15807 14433
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 3326 14396 3332 14408
rect 3287 14368 3332 14396
rect 3326 14356 3332 14368
rect 3384 14356 3390 14408
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 5534 14396 5540 14408
rect 5495 14368 5540 14396
rect 4617 14359 4675 14365
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 4632 14328 4660 14359
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14396 16543 14399
rect 17034 14396 17040 14408
rect 16531 14368 17040 14396
rect 16531 14365 16543 14368
rect 16485 14359 16543 14365
rect 17034 14356 17040 14368
rect 17092 14356 17098 14408
rect 17494 14396 17500 14408
rect 17455 14368 17500 14396
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14365 17739 14399
rect 17681 14359 17739 14365
rect 4212 14300 4660 14328
rect 15289 14331 15347 14337
rect 4212 14288 4218 14300
rect 15289 14297 15301 14331
rect 15335 14328 15347 14331
rect 17126 14328 17132 14340
rect 15335 14300 17132 14328
rect 15335 14297 15347 14300
rect 15289 14291 15347 14297
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 2958 14220 2964 14272
rect 3016 14260 3022 14272
rect 4065 14263 4123 14269
rect 4065 14260 4077 14263
rect 3016 14232 4077 14260
rect 3016 14220 3022 14232
rect 4065 14229 4077 14232
rect 4111 14229 4123 14263
rect 4065 14223 4123 14229
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 7377 14263 7435 14269
rect 7377 14260 7389 14263
rect 6420 14232 7389 14260
rect 6420 14220 6426 14232
rect 7377 14229 7389 14232
rect 7423 14229 7435 14263
rect 7377 14223 7435 14229
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 11793 14263 11851 14269
rect 11793 14260 11805 14263
rect 11664 14232 11805 14260
rect 11664 14220 11670 14232
rect 11793 14229 11805 14232
rect 11839 14229 11851 14263
rect 17696 14260 17724 14359
rect 18782 14260 18788 14272
rect 17696 14232 18788 14260
rect 11793 14223 11851 14229
rect 18782 14220 18788 14232
rect 18840 14260 18846 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 18840 14232 19441 14260
rect 18840 14220 18846 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2498 14056 2504 14068
rect 2459 14028 2504 14056
rect 2498 14016 2504 14028
rect 2556 14016 2562 14068
rect 3160 14028 4936 14056
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3160 13929 3188 14028
rect 4908 13997 4936 14028
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5132 14028 5733 14056
rect 5132 14016 5138 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 9401 14059 9459 14065
rect 5721 14019 5779 14025
rect 5828 14028 8984 14056
rect 4893 13991 4951 13997
rect 4893 13957 4905 13991
rect 4939 13988 4951 13991
rect 5828 13988 5856 14028
rect 4939 13960 5856 13988
rect 8956 13988 8984 14028
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9674 14056 9680 14068
rect 9447 14028 9680 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 11790 14056 11796 14068
rect 9815 14028 11796 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12621 14059 12679 14065
rect 12621 14025 12633 14059
rect 12667 14056 12679 14059
rect 13538 14056 13544 14068
rect 12667 14028 13544 14056
rect 12667 14025 12679 14028
rect 12621 14019 12679 14025
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 16022 14056 16028 14068
rect 15672 14028 16028 14056
rect 8956 13960 11836 13988
rect 4939 13957 4951 13960
rect 4893 13951 4951 13957
rect 11808 13932 11836 13960
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 6362 13920 6368 13932
rect 6323 13892 6368 13920
rect 3145 13883 3203 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 7466 13920 7472 13932
rect 7427 13892 7472 13920
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 10410 13920 10416 13932
rect 10371 13892 10416 13920
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11241 13923 11299 13929
rect 11241 13920 11253 13923
rect 11112 13892 11253 13920
rect 11112 13880 11118 13892
rect 11241 13889 11253 13892
rect 11287 13889 11299 13923
rect 11241 13883 11299 13889
rect 11425 13923 11483 13929
rect 11425 13889 11437 13923
rect 11471 13920 11483 13923
rect 11606 13920 11612 13932
rect 11471 13892 11612 13920
rect 11471 13889 11483 13892
rect 11425 13883 11483 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11790 13880 11796 13932
rect 11848 13880 11854 13932
rect 13262 13920 13268 13932
rect 13223 13892 13268 13920
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 15672 13929 15700 14028
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 16356 14028 16620 14056
rect 16356 14016 16362 14028
rect 16592 13988 16620 14028
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17037 14059 17095 14065
rect 17037 14056 17049 14059
rect 17000 14028 17049 14056
rect 17000 14016 17006 14028
rect 17037 14025 17049 14028
rect 17083 14025 17095 14059
rect 17037 14019 17095 14025
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 17552 14028 18061 14056
rect 17552 14016 17558 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 16592 13960 17908 13988
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13412 13892 14289 13920
rect 13412 13880 13418 13892
rect 14277 13889 14289 13892
rect 14323 13920 14335 13923
rect 15197 13923 15255 13929
rect 15197 13920 15209 13923
rect 14323 13892 15209 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 15197 13889 15209 13892
rect 15243 13889 15255 13923
rect 15197 13883 15255 13889
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13889 15715 13923
rect 15657 13883 15715 13889
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13852 1823 13855
rect 2869 13855 2927 13861
rect 1811 13824 2820 13852
rect 1811 13821 1823 13824
rect 1765 13815 1823 13821
rect 2792 13784 2820 13824
rect 2869 13821 2881 13855
rect 2915 13852 2927 13855
rect 3326 13852 3332 13864
rect 2915 13824 3332 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 3510 13852 3516 13864
rect 3471 13824 3516 13852
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 3780 13855 3838 13861
rect 3780 13821 3792 13855
rect 3826 13852 3838 13855
rect 4154 13852 4160 13864
rect 3826 13824 4160 13852
rect 3826 13821 3838 13824
rect 3780 13815 3838 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 4264 13824 5488 13852
rect 4264 13784 4292 13824
rect 2792 13756 4292 13784
rect 5460 13784 5488 13824
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5592 13824 6101 13852
rect 5592 13812 5598 13824
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 7006 13852 7012 13864
rect 6089 13815 6147 13821
rect 6196 13824 7012 13852
rect 6196 13784 6224 13824
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 7650 13852 7656 13864
rect 7331 13824 7656 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 8021 13855 8079 13861
rect 8021 13821 8033 13855
rect 8067 13852 8079 13855
rect 8846 13852 8852 13864
rect 8067 13824 8852 13852
rect 8067 13821 8079 13824
rect 8021 13815 8079 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14093 13855 14151 13861
rect 14093 13852 14105 13855
rect 13964 13824 14105 13852
rect 13964 13812 13970 13824
rect 14093 13821 14105 13824
rect 14139 13821 14151 13855
rect 15102 13852 15108 13864
rect 15063 13824 15108 13852
rect 14093 13815 14151 13821
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15930 13861 15936 13864
rect 15924 13852 15936 13861
rect 15843 13824 15936 13852
rect 15924 13815 15936 13824
rect 15988 13852 15994 13864
rect 17218 13852 17224 13864
rect 15988 13824 17224 13852
rect 15930 13812 15936 13815
rect 15988 13812 15994 13824
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 5460 13756 6224 13784
rect 8288 13787 8346 13793
rect 8288 13753 8300 13787
rect 8334 13784 8346 13787
rect 8662 13784 8668 13796
rect 8334 13756 8668 13784
rect 8334 13753 8346 13756
rect 8288 13747 8346 13753
rect 8662 13744 8668 13756
rect 8720 13744 8726 13796
rect 10137 13787 10195 13793
rect 10137 13753 10149 13787
rect 10183 13784 10195 13787
rect 11146 13784 11152 13796
rect 10183 13756 11008 13784
rect 11107 13756 11152 13784
rect 10183 13753 10195 13756
rect 10137 13747 10195 13753
rect 6181 13719 6239 13725
rect 6181 13685 6193 13719
rect 6227 13716 6239 13719
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 6227 13688 6837 13716
rect 6227 13685 6239 13688
rect 6181 13679 6239 13685
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 6825 13679 6883 13685
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 7156 13688 7205 13716
rect 7156 13676 7162 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 10229 13719 10287 13725
rect 10229 13685 10241 13719
rect 10275 13716 10287 13719
rect 10781 13719 10839 13725
rect 10781 13716 10793 13719
rect 10275 13688 10793 13716
rect 10275 13685 10287 13688
rect 10229 13679 10287 13685
rect 10781 13685 10793 13688
rect 10827 13685 10839 13719
rect 10980 13716 11008 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 12526 13784 12532 13796
rect 11296 13756 12532 13784
rect 11296 13744 11302 13756
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 12989 13787 13047 13793
rect 12989 13753 13001 13787
rect 13035 13784 13047 13787
rect 15010 13784 15016 13796
rect 13035 13756 14688 13784
rect 14971 13756 15016 13784
rect 13035 13753 13047 13756
rect 12989 13747 13047 13753
rect 11054 13716 11060 13728
rect 10980 13688 11060 13716
rect 10781 13679 10839 13685
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 13081 13719 13139 13725
rect 13081 13685 13093 13719
rect 13127 13716 13139 13719
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13127 13688 13645 13716
rect 13127 13685 13139 13688
rect 13081 13679 13139 13685
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 13633 13679 13691 13685
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14660 13725 14688 13756
rect 15010 13744 15016 13756
rect 15068 13744 15074 13796
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13872 13688 14013 13716
rect 13872 13676 13878 13688
rect 14001 13685 14013 13688
rect 14047 13685 14059 13719
rect 14001 13679 14059 13685
rect 14645 13719 14703 13725
rect 14645 13685 14657 13719
rect 14691 13685 14703 13719
rect 17880 13716 17908 13960
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 18417 13855 18475 13861
rect 18417 13821 18429 13855
rect 18463 13852 18475 13855
rect 18506 13852 18512 13864
rect 18463 13824 18512 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 18506 13812 18512 13824
rect 18564 13852 18570 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18564 13824 18889 13852
rect 18564 13812 18570 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 19061 13787 19119 13793
rect 19061 13784 19073 13787
rect 18012 13756 19073 13784
rect 18012 13744 18018 13756
rect 19061 13753 19073 13756
rect 19107 13753 19119 13787
rect 19061 13747 19119 13753
rect 18509 13719 18567 13725
rect 18509 13716 18521 13719
rect 17880 13688 18521 13716
rect 14645 13679 14703 13685
rect 18509 13685 18521 13688
rect 18555 13685 18567 13719
rect 18509 13679 18567 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1581 13515 1639 13521
rect 1581 13481 1593 13515
rect 1627 13512 1639 13515
rect 1854 13512 1860 13524
rect 1627 13484 1860 13512
rect 1627 13481 1639 13484
rect 1581 13475 1639 13481
rect 1854 13472 1860 13484
rect 1912 13472 1918 13524
rect 6178 13512 6184 13524
rect 1964 13484 6184 13512
rect 1964 13385 1992 13484
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 6270 13472 6276 13524
rect 6328 13512 6334 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 6328 13484 6561 13512
rect 6328 13472 6334 13484
rect 6549 13481 6561 13484
rect 6595 13481 6607 13515
rect 7742 13512 7748 13524
rect 7703 13484 7748 13512
rect 6549 13475 6607 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 11238 13512 11244 13524
rect 7852 13484 11244 13512
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 7852 13444 7880 13484
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13630 13512 13636 13524
rect 13320 13484 13636 13512
rect 13320 13472 13326 13484
rect 13630 13472 13636 13484
rect 13688 13512 13694 13524
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 13688 13484 14197 13512
rect 13688 13472 13694 13484
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 14458 13512 14464 13524
rect 14419 13484 14464 13512
rect 14185 13475 14243 13481
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 15657 13515 15715 13521
rect 15657 13481 15669 13515
rect 15703 13512 15715 13515
rect 15746 13512 15752 13524
rect 15703 13484 15752 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 16666 13512 16672 13524
rect 16627 13484 16672 13512
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 17126 13512 17132 13524
rect 17087 13484 17132 13512
rect 17126 13472 17132 13484
rect 17184 13472 17190 13524
rect 10778 13444 10784 13456
rect 4120 13416 7880 13444
rect 10739 13416 10784 13444
rect 4120 13404 4126 13416
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13444 12587 13447
rect 17034 13444 17040 13456
rect 12575 13416 14688 13444
rect 16995 13416 17040 13444
rect 12575 13413 12587 13416
rect 12529 13407 12587 13413
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1397 13339 1455 13345
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13345 2007 13379
rect 1949 13339 2007 13345
rect 5436 13379 5494 13385
rect 5436 13345 5448 13379
rect 5482 13376 5494 13379
rect 5994 13376 6000 13388
rect 5482 13348 6000 13376
rect 5482 13345 5494 13348
rect 5436 13339 5494 13345
rect 1412 13308 1440 13339
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13376 7435 13379
rect 7742 13376 7748 13388
rect 7423 13348 7748 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 7929 13379 7987 13385
rect 7929 13345 7941 13379
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 8435 13348 9045 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 9033 13345 9045 13348
rect 9079 13345 9091 13379
rect 9033 13339 9091 13345
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 1412 13280 2145 13308
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 2133 13271 2191 13277
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 4764 13280 5181 13308
rect 4764 13268 4770 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 7944 13240 7972 13339
rect 8478 13308 8484 13320
rect 8439 13280 8484 13308
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 12544 13240 12572 13407
rect 13072 13379 13130 13385
rect 13072 13345 13084 13379
rect 13118 13376 13130 13379
rect 13354 13376 13360 13388
rect 13118 13348 13360 13376
rect 13118 13345 13130 13348
rect 13072 13339 13130 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 14660 13385 14688 13416
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 14645 13379 14703 13385
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 16025 13379 16083 13385
rect 16025 13345 16037 13379
rect 16071 13376 16083 13379
rect 16850 13376 16856 13388
rect 16071 13348 16856 13376
rect 16071 13345 16083 13348
rect 16025 13339 16083 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17000 13348 17264 13376
rect 17000 13336 17006 13348
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 12768 13280 12817 13308
rect 12768 13268 12774 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 15746 13308 15752 13320
rect 13872 13280 15752 13308
rect 13872 13268 13878 13280
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16114 13308 16120 13320
rect 16075 13280 16120 13308
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13308 16359 13311
rect 16758 13308 16764 13320
rect 16347 13280 16764 13308
rect 16347 13277 16359 13280
rect 16301 13271 16359 13277
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 17236 13317 17264 13348
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 7064 13212 7328 13240
rect 7944 13212 12572 13240
rect 7064 13200 7070 13212
rect 7190 13172 7196 13184
rect 7151 13144 7196 13172
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 7300 13172 7328 13212
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 7300 13144 8033 13172
rect 8021 13141 8033 13144
rect 8067 13141 8079 13175
rect 8021 13135 8079 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 2590 12968 2596 12980
rect 2547 12940 2596 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6089 12971 6147 12977
rect 6089 12968 6101 12971
rect 6052 12940 6101 12968
rect 6052 12928 6058 12940
rect 6089 12937 6101 12940
rect 6135 12937 6147 12971
rect 6089 12931 6147 12937
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 2866 12900 2872 12912
rect 1995 12872 2872 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 4706 12832 4712 12844
rect 4667 12804 4712 12832
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 6104 12832 6132 12931
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6236 12940 6837 12968
rect 6236 12928 6242 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 8720 12940 9321 12968
rect 8720 12928 8726 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 11425 12971 11483 12977
rect 11425 12968 11437 12971
rect 10468 12940 11437 12968
rect 10468 12928 10474 12940
rect 11425 12937 11437 12940
rect 11471 12937 11483 12971
rect 11425 12931 11483 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13446 12968 13452 12980
rect 13127 12940 13452 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 17218 12968 17224 12980
rect 17179 12940 17224 12968
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 11517 12903 11575 12909
rect 11517 12900 11529 12903
rect 11112 12872 11529 12900
rect 11112 12860 11118 12872
rect 11517 12869 11529 12872
rect 11563 12869 11575 12903
rect 11517 12863 11575 12869
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6104 12804 7389 12832
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 13630 12832 13636 12844
rect 13591 12804 13636 12832
rect 12069 12795 12127 12801
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2317 12767 2375 12773
rect 2317 12733 2329 12767
rect 2363 12764 2375 12767
rect 2958 12764 2964 12776
rect 2363 12736 2964 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7708 12736 7941 12764
rect 7708 12724 7714 12736
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 10042 12764 10048 12776
rect 10003 12736 10048 12764
rect 7929 12727 7987 12733
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10312 12767 10370 12773
rect 10312 12733 10324 12767
rect 10358 12764 10370 12767
rect 11606 12764 11612 12776
rect 10358 12736 11612 12764
rect 10358 12733 10370 12736
rect 10312 12727 10370 12733
rect 11606 12724 11612 12736
rect 11664 12764 11670 12776
rect 12084 12764 12112 12795
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 11664 12736 12112 12764
rect 11664 12724 11670 12736
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 15378 12764 15384 12776
rect 12584 12736 15384 12764
rect 12584 12724 12590 12736
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 15841 12767 15899 12773
rect 15841 12764 15853 12767
rect 15528 12736 15853 12764
rect 15528 12724 15534 12736
rect 15841 12733 15853 12736
rect 15887 12733 15899 12767
rect 15841 12727 15899 12733
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 18012 12736 18061 12764
rect 18012 12724 18018 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 18316 12767 18374 12773
rect 18316 12733 18328 12767
rect 18362 12764 18374 12767
rect 18782 12764 18788 12776
rect 18362 12736 18788 12764
rect 18362 12733 18374 12736
rect 18316 12727 18374 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 4976 12699 5034 12705
rect 4976 12665 4988 12699
rect 5022 12696 5034 12699
rect 5442 12696 5448 12708
rect 5022 12668 5448 12696
rect 5022 12665 5034 12668
rect 4976 12659 5034 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 5736 12668 7205 12696
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12628 4307 12631
rect 5736 12628 5764 12668
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 8196 12699 8254 12705
rect 8196 12665 8208 12699
rect 8242 12696 8254 12699
rect 9122 12696 9128 12708
rect 8242 12668 9128 12696
rect 8242 12665 8254 12668
rect 8196 12659 8254 12665
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 11885 12699 11943 12705
rect 11885 12665 11897 12699
rect 11931 12696 11943 12699
rect 12437 12699 12495 12705
rect 12437 12696 12449 12699
rect 11931 12668 12449 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 12437 12665 12449 12668
rect 12483 12665 12495 12699
rect 12437 12659 12495 12665
rect 13449 12699 13507 12705
rect 13449 12665 13461 12699
rect 13495 12696 13507 12699
rect 14093 12699 14151 12705
rect 14093 12696 14105 12699
rect 13495 12668 14105 12696
rect 13495 12665 13507 12668
rect 13449 12659 13507 12665
rect 14093 12665 14105 12668
rect 14139 12665 14151 12699
rect 14093 12659 14151 12665
rect 16108 12699 16166 12705
rect 16108 12665 16120 12699
rect 16154 12696 16166 12699
rect 16758 12696 16764 12708
rect 16154 12668 16764 12696
rect 16154 12665 16166 12668
rect 16108 12659 16166 12665
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 4295 12600 5764 12628
rect 4295 12597 4307 12600
rect 4249 12591 4307 12597
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 11974 12628 11980 12640
rect 7340 12600 7385 12628
rect 11935 12600 11980 12628
rect 7340 12588 7346 12600
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 13538 12588 13544 12640
rect 13596 12628 13602 12640
rect 19426 12628 19432 12640
rect 13596 12600 13641 12628
rect 19387 12600 19432 12628
rect 13596 12588 13602 12600
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 3988 12396 7573 12424
rect 1762 12316 1768 12368
rect 1820 12356 1826 12368
rect 2225 12359 2283 12365
rect 2225 12356 2237 12359
rect 1820 12328 2237 12356
rect 1820 12316 1826 12328
rect 2225 12325 2237 12328
rect 2271 12325 2283 12359
rect 2958 12356 2964 12368
rect 2919 12328 2964 12356
rect 2225 12319 2283 12325
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1854 12288 1860 12300
rect 1443 12260 1860 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12257 2007 12291
rect 2682 12288 2688 12300
rect 2643 12260 2688 12288
rect 1949 12251 2007 12257
rect 1964 12220 1992 12251
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 3988 12220 4016 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 7561 12387 7619 12393
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8536 12396 8585 12424
rect 8536 12384 8542 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 8573 12387 8631 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 11974 12424 11980 12436
rect 9140 12396 11980 12424
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 4120 12328 4476 12356
rect 4120 12316 4126 12328
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4321 12291 4379 12297
rect 4321 12288 4333 12291
rect 4212 12260 4333 12288
rect 4212 12248 4218 12260
rect 4321 12257 4333 12260
rect 4367 12257 4379 12291
rect 4448 12288 4476 12328
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 5534 12356 5540 12368
rect 4764 12328 5540 12356
rect 4764 12316 4770 12328
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 5988 12359 6046 12365
rect 5988 12325 6000 12359
rect 6034 12356 6046 12359
rect 6546 12356 6552 12368
rect 6034 12328 6552 12356
rect 6034 12325 6046 12328
rect 5988 12319 6046 12325
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 9140 12356 9168 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13538 12424 13544 12436
rect 13035 12396 13544 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 16758 12424 16764 12436
rect 14056 12396 15976 12424
rect 16719 12396 16764 12424
rect 14056 12384 14062 12396
rect 6656 12328 9168 12356
rect 6656 12288 6684 12328
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 10750 12359 10808 12365
rect 10750 12356 10762 12359
rect 10468 12328 10762 12356
rect 10468 12316 10474 12328
rect 10750 12325 10762 12328
rect 10796 12325 10808 12359
rect 12526 12356 12532 12368
rect 12487 12328 12532 12356
rect 10750 12319 10808 12325
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 15654 12365 15660 12368
rect 13357 12359 13415 12365
rect 13357 12325 13369 12359
rect 13403 12356 13415 12359
rect 15637 12359 15660 12365
rect 13403 12328 13472 12356
rect 13403 12325 13415 12328
rect 13357 12319 13415 12325
rect 4448 12260 6684 12288
rect 4321 12251 4379 12257
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 6880 12260 7941 12288
rect 6880 12248 6886 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12288 8079 12291
rect 8478 12288 8484 12300
rect 8067 12260 8484 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12257 8999 12291
rect 8941 12251 8999 12257
rect 1964 12192 4016 12220
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 2314 12112 2320 12164
rect 2372 12152 2378 12164
rect 4080 12152 4108 12183
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5721 12223 5779 12229
rect 5721 12220 5733 12223
rect 5592 12192 5733 12220
rect 5592 12180 5598 12192
rect 5721 12189 5733 12192
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 8202 12220 8208 12232
rect 7156 12192 7236 12220
rect 8163 12192 8208 12220
rect 7156 12180 7162 12192
rect 2372 12124 4108 12152
rect 2372 12112 2378 12124
rect 4080 12084 4108 12124
rect 5276 12124 5764 12152
rect 4246 12084 4252 12096
rect 4080 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 5276 12084 5304 12124
rect 5442 12084 5448 12096
rect 4764 12056 5304 12084
rect 5403 12056 5448 12084
rect 4764 12044 4770 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5736 12084 5764 12124
rect 7098 12084 7104 12096
rect 5736 12056 7104 12084
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7208 12084 7236 12192
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 7558 12112 7564 12164
rect 7616 12152 7622 12164
rect 8956 12152 8984 12251
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10100 12260 10517 12288
rect 10100 12248 10106 12260
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 10505 12251 10563 12257
rect 11146 12248 11152 12300
rect 11204 12288 11210 12300
rect 12253 12291 12311 12297
rect 12253 12288 12265 12291
rect 11204 12260 12265 12288
rect 11204 12248 11210 12260
rect 12253 12257 12265 12260
rect 12299 12257 12311 12291
rect 13444 12288 13472 12328
rect 15637 12325 15649 12359
rect 15637 12319 15660 12325
rect 15654 12316 15660 12319
rect 15712 12316 15718 12368
rect 15948 12356 15976 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 16908 12396 17049 12424
rect 16908 12384 16914 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 17037 12387 17095 12393
rect 17144 12396 18153 12424
rect 17144 12356 17172 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18141 12387 18199 12393
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 15948 12328 17172 12356
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 19061 12359 19119 12365
rect 19061 12356 19073 12359
rect 17828 12328 19073 12356
rect 17828 12316 17834 12328
rect 19061 12325 19073 12328
rect 19107 12325 19119 12359
rect 19061 12319 19119 12325
rect 13538 12288 13544 12300
rect 13444 12260 13544 12288
rect 12253 12251 12311 12257
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 14458 12288 14464 12300
rect 14419 12260 14464 12288
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 16666 12288 16672 12300
rect 14660 12260 16672 12288
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 10410 12220 10416 12232
rect 9324 12192 10416 12220
rect 7616 12124 8984 12152
rect 7616 12112 7622 12124
rect 9324 12084 9352 12192
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12189 13507 12223
rect 13630 12220 13636 12232
rect 13591 12192 13636 12220
rect 13449 12183 13507 12189
rect 12802 12112 12808 12164
rect 12860 12152 12866 12164
rect 13464 12152 13492 12183
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 13872 12192 14565 12220
rect 13872 12180 13878 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14660 12152 14688 12260
rect 16666 12248 16672 12260
rect 16724 12288 16730 12300
rect 18049 12291 18107 12297
rect 18049 12288 18061 12291
rect 16724 12260 18061 12288
rect 16724 12248 16730 12260
rect 18049 12257 18061 12260
rect 18095 12257 18107 12291
rect 19426 12288 19432 12300
rect 18049 12251 18107 12257
rect 18340 12260 19432 12288
rect 15378 12220 15384 12232
rect 15339 12192 15384 12220
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 18340 12229 18368 12260
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 19153 12223 19211 12229
rect 19153 12189 19165 12223
rect 19199 12189 19211 12223
rect 19153 12183 19211 12189
rect 12860 12124 14688 12152
rect 17681 12155 17739 12161
rect 12860 12112 12866 12124
rect 17681 12121 17693 12155
rect 17727 12152 17739 12155
rect 19168 12152 19196 12183
rect 19242 12180 19248 12232
rect 19300 12220 19306 12232
rect 19300 12192 19345 12220
rect 19300 12180 19306 12192
rect 17727 12124 19196 12152
rect 17727 12121 17739 12124
rect 17681 12115 17739 12121
rect 7208 12056 9352 12084
rect 10502 12044 10508 12096
rect 10560 12084 10566 12096
rect 11882 12084 11888 12096
rect 10560 12056 11888 12084
rect 10560 12044 10566 12056
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 13136 12056 14289 12084
rect 13136 12044 13142 12056
rect 14277 12053 14289 12056
rect 14323 12084 14335 12087
rect 17310 12084 17316 12096
rect 14323 12056 17316 12084
rect 14323 12053 14335 12056
rect 14277 12047 14335 12053
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 2740 11852 4353 11880
rect 2740 11840 2746 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 4341 11843 4399 11849
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 7282 11880 7288 11892
rect 5675 11852 7288 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9309 11883 9367 11889
rect 9309 11880 9321 11883
rect 9180 11852 9321 11880
rect 9180 11840 9186 11852
rect 9309 11849 9321 11852
rect 9355 11849 9367 11883
rect 11146 11880 11152 11892
rect 11107 11852 11152 11880
rect 9309 11843 9367 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 13449 11883 13507 11889
rect 13449 11849 13461 11883
rect 13495 11880 13507 11883
rect 14090 11880 14096 11892
rect 13495 11852 14096 11880
rect 13495 11849 13507 11852
rect 13449 11843 13507 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14369 11883 14427 11889
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 14415 11852 15516 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 15488 11824 15516 11852
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15712 11852 15853 11880
rect 15712 11840 15718 11852
rect 15841 11849 15853 11852
rect 15887 11880 15899 11883
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 15887 11852 15945 11880
rect 15887 11849 15899 11852
rect 15841 11843 15899 11849
rect 15933 11849 15945 11852
rect 15979 11849 15991 11883
rect 16114 11880 16120 11892
rect 16075 11852 16120 11880
rect 15933 11843 15991 11849
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 18064 11852 19748 11880
rect 4065 11815 4123 11821
rect 4065 11781 4077 11815
rect 4111 11812 4123 11815
rect 4154 11812 4160 11824
rect 4111 11784 4160 11812
rect 4111 11781 4123 11784
rect 4065 11775 4123 11781
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 4080 11744 4108 11775
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 10137 11815 10195 11821
rect 4991 11784 7512 11812
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4080 11716 4905 11744
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2685 11679 2743 11685
rect 2685 11676 2697 11679
rect 2372 11648 2697 11676
rect 2372 11636 2378 11648
rect 2685 11645 2697 11648
rect 2731 11645 2743 11679
rect 2685 11639 2743 11645
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 4991 11676 5019 11784
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 6181 11747 6239 11753
rect 6181 11744 6193 11747
rect 5500 11716 6193 11744
rect 5500 11704 5506 11716
rect 6181 11713 6193 11716
rect 6227 11713 6239 11747
rect 6181 11707 6239 11713
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6696 11716 7052 11744
rect 6696 11704 6702 11716
rect 4120 11648 5019 11676
rect 6089 11679 6147 11685
rect 4120 11636 4126 11648
rect 6089 11645 6101 11679
rect 6135 11676 6147 11679
rect 6730 11676 6736 11688
rect 6135 11648 6736 11676
rect 6135 11645 6147 11648
rect 6089 11639 6147 11645
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 7024 11676 7052 11716
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 7156 11716 7389 11744
rect 7156 11704 7162 11716
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 7484 11744 7512 11784
rect 10137 11781 10149 11815
rect 10183 11812 10195 11815
rect 10183 11784 11560 11812
rect 10183 11781 10195 11784
rect 10137 11775 10195 11781
rect 7484 11716 8064 11744
rect 7377 11707 7435 11713
rect 7558 11676 7564 11688
rect 7024 11648 7564 11676
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 7650 11636 7656 11688
rect 7708 11676 7714 11688
rect 7929 11679 7987 11685
rect 7929 11676 7941 11679
rect 7708 11648 7941 11676
rect 7708 11636 7714 11648
rect 7929 11645 7941 11648
rect 7975 11645 7987 11679
rect 8036 11676 8064 11716
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10560 11716 10701 11744
rect 10560 11704 10566 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 11532 11685 11560 11784
rect 15470 11772 15476 11824
rect 15528 11812 15534 11824
rect 16206 11812 16212 11824
rect 15528 11784 16212 11812
rect 15528 11772 15534 11784
rect 16206 11772 16212 11784
rect 16264 11812 16270 11824
rect 17129 11815 17187 11821
rect 17129 11812 17141 11815
rect 16264 11784 17141 11812
rect 16264 11772 16270 11784
rect 17129 11781 17141 11784
rect 17175 11812 17187 11815
rect 17954 11812 17960 11824
rect 17175 11784 17960 11812
rect 17175 11781 17187 11784
rect 17129 11775 17187 11781
rect 17954 11772 17960 11784
rect 18012 11812 18018 11824
rect 18064 11812 18092 11852
rect 18012 11784 18092 11812
rect 18012 11772 18018 11784
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11664 11716 11713 11744
rect 11664 11704 11670 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 11940 11716 13001 11744
rect 11940 11704 11946 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 18064 11753 18092 11784
rect 19720 11753 19748 11852
rect 14093 11747 14151 11753
rect 13688 11716 13952 11744
rect 13688 11704 13694 11716
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 8036 11648 10609 11676
rect 7929 11639 7987 11645
rect 10597 11645 10609 11648
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 11517 11679 11575 11685
rect 11517 11645 11529 11679
rect 11563 11645 11575 11679
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 11517 11639 11575 11645
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 13814 11676 13820 11688
rect 13775 11648 13820 11676
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 13924 11676 13952 11716
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 15933 11747 15991 11753
rect 14139 11716 14596 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14568 11688 14596 11716
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15979 11716 16681 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 14369 11679 14427 11685
rect 13924 11648 14136 11676
rect 2952 11611 3010 11617
rect 2952 11577 2964 11611
rect 2998 11608 3010 11611
rect 4614 11608 4620 11620
rect 2998 11580 4620 11608
rect 2998 11577 3010 11580
rect 2952 11571 3010 11577
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 4801 11611 4859 11617
rect 4801 11577 4813 11611
rect 4847 11608 4859 11611
rect 4847 11580 6868 11608
rect 4847 11577 4859 11580
rect 4801 11571 4859 11577
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5776 11512 6009 11540
rect 5776 11500 5782 11512
rect 5997 11509 6009 11512
rect 6043 11540 6055 11543
rect 6638 11540 6644 11552
rect 6043 11512 6644 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 6840 11549 6868 11580
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 8202 11617 8208 11620
rect 7285 11611 7343 11617
rect 7285 11608 7297 11611
rect 6972 11580 7297 11608
rect 6972 11568 6978 11580
rect 7285 11577 7297 11580
rect 7331 11577 7343 11611
rect 8196 11608 8208 11617
rect 8115 11580 8208 11608
rect 7285 11571 7343 11577
rect 8196 11571 8208 11580
rect 8260 11608 8266 11620
rect 9030 11608 9036 11620
rect 8260 11580 9036 11608
rect 8202 11568 8208 11571
rect 8260 11568 8266 11580
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 9677 11611 9735 11617
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 10505 11611 10563 11617
rect 10505 11608 10517 11611
rect 9723 11580 10517 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 10505 11577 10517 11580
rect 10551 11577 10563 11611
rect 10505 11571 10563 11577
rect 12897 11611 12955 11617
rect 12897 11577 12909 11611
rect 12943 11608 12955 11611
rect 13998 11608 14004 11620
rect 12943 11580 14004 11608
rect 12943 11577 12955 11580
rect 12897 11571 12955 11577
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 14108 11608 14136 11648
rect 14369 11645 14381 11679
rect 14415 11676 14427 11679
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 14415 11648 14473 11676
rect 14415 11645 14427 11648
rect 14369 11639 14427 11645
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 14717 11679 14775 11685
rect 14717 11676 14729 11679
rect 14608 11648 14729 11676
rect 14608 11636 14614 11648
rect 14717 11645 14729 11648
rect 14763 11645 14775 11679
rect 14717 11639 14775 11645
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 16577 11679 16635 11685
rect 16577 11676 16589 11679
rect 15620 11648 16589 11676
rect 15620 11636 15626 11648
rect 16577 11645 16589 11648
rect 16623 11645 16635 11679
rect 17310 11676 17316 11688
rect 17271 11648 17316 11676
rect 16577 11639 16635 11645
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 18316 11679 18374 11685
rect 18316 11645 18328 11679
rect 18362 11676 18374 11679
rect 19426 11676 19432 11688
rect 18362 11648 19432 11676
rect 18362 11645 18374 11648
rect 18316 11639 18374 11645
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 19978 11617 19984 11620
rect 19972 11608 19984 11617
rect 14108 11580 19564 11608
rect 19939 11580 19984 11608
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 7156 11512 7205 11540
rect 7156 11500 7162 11512
rect 7193 11509 7205 11512
rect 7239 11540 7251 11543
rect 8846 11540 8852 11552
rect 7239 11512 8852 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 11609 11543 11667 11549
rect 11609 11509 11621 11543
rect 11655 11540 11667 11543
rect 12437 11543 12495 11549
rect 12437 11540 12449 11543
rect 11655 11512 12449 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 12437 11509 12449 11512
rect 12483 11509 12495 11543
rect 12437 11503 12495 11509
rect 13909 11543 13967 11549
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 15286 11540 15292 11552
rect 13955 11512 15292 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 15436 11512 16497 11540
rect 15436 11500 15442 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16485 11503 16543 11509
rect 17497 11543 17555 11549
rect 17497 11509 17509 11543
rect 17543 11540 17555 11543
rect 18138 11540 18144 11552
rect 17543 11512 18144 11540
rect 17543 11509 17555 11512
rect 17497 11503 17555 11509
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 19208 11512 19441 11540
rect 19208 11500 19214 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19536 11540 19564 11580
rect 19972 11571 19984 11580
rect 19978 11568 19984 11571
rect 20036 11568 20042 11620
rect 21085 11543 21143 11549
rect 21085 11540 21097 11543
rect 19536 11512 21097 11540
rect 19429 11503 19487 11509
rect 21085 11509 21097 11512
rect 21131 11509 21143 11543
rect 21085 11503 21143 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 2774 11336 2780 11348
rect 1627 11308 2780 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 4065 11339 4123 11345
rect 4065 11305 4077 11339
rect 4111 11336 4123 11339
rect 4706 11336 4712 11348
rect 4111 11308 4712 11336
rect 4111 11305 4123 11308
rect 4065 11299 4123 11305
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 9030 11336 9036 11348
rect 8991 11308 9036 11336
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 11885 11339 11943 11345
rect 11885 11305 11897 11339
rect 11931 11336 11943 11339
rect 13262 11336 13268 11348
rect 11931 11308 13268 11336
rect 11931 11305 11943 11308
rect 11885 11299 11943 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14608 11308 14933 11336
rect 14608 11296 14614 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 14921 11299 14979 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15746 11336 15752 11348
rect 15707 11308 15752 11336
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 17770 11336 17776 11348
rect 17731 11308 17776 11336
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 18138 11336 18144 11348
rect 18099 11308 18144 11336
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 7009 11271 7067 11277
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 9677 11271 9735 11277
rect 9677 11268 9689 11271
rect 7055 11240 9689 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 9677 11237 9689 11240
rect 9723 11237 9735 11271
rect 12342 11268 12348 11280
rect 9677 11231 9735 11237
rect 9784 11240 10640 11268
rect 12303 11240 12348 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11169 1455 11203
rect 1397 11163 1455 11169
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 3237 11203 3295 11209
rect 1995 11172 3188 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 1412 11132 1440 11163
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1412 11104 2145 11132
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 3160 11064 3188 11172
rect 3237 11169 3249 11203
rect 3283 11200 3295 11203
rect 4154 11200 4160 11212
rect 3283 11172 4160 11200
rect 3283 11169 3295 11172
rect 3237 11163 3295 11169
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 5077 11203 5135 11209
rect 5077 11200 5089 11203
rect 4479 11172 5089 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 5077 11169 5089 11172
rect 5123 11169 5135 11203
rect 5077 11163 5135 11169
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 6914 11200 6920 11212
rect 5767 11172 6920 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 6914 11160 6920 11172
rect 6972 11200 6978 11212
rect 7190 11200 7196 11212
rect 6972 11172 7196 11200
rect 6972 11160 6978 11172
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7926 11209 7932 11212
rect 7920 11200 7932 11209
rect 7300 11172 7932 11200
rect 3326 11132 3332 11144
rect 3287 11104 3332 11132
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 3694 11132 3700 11144
rect 3559 11104 3700 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 3694 11092 3700 11104
rect 3752 11092 3758 11144
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4706 11132 4712 11144
rect 4667 11104 4712 11132
rect 4525 11095 4583 11101
rect 4246 11064 4252 11076
rect 3160 11036 4252 11064
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4540 11064 4568 11095
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 7300 11141 7328 11172
rect 7920 11163 7932 11172
rect 7926 11160 7932 11163
rect 7984 11160 7990 11212
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 9784 11200 9812 11240
rect 10502 11209 10508 11212
rect 10496 11200 10508 11209
rect 8260 11172 9812 11200
rect 10463 11172 10508 11200
rect 8260 11160 8266 11172
rect 10496 11163 10508 11172
rect 10502 11160 10508 11163
rect 10560 11160 10566 11212
rect 10612 11200 10640 11240
rect 12342 11228 12348 11240
rect 12400 11228 12406 11280
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 10612 11172 12265 11200
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 13078 11200 13084 11212
rect 13039 11172 13084 11200
rect 12253 11163 12311 11169
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 13808 11203 13866 11209
rect 13808 11169 13820 11203
rect 13854 11200 13866 11203
rect 15654 11200 15660 11212
rect 13854 11172 14596 11200
rect 15615 11172 15660 11200
rect 13854 11169 13866 11172
rect 13808 11163 13866 11169
rect 14568 11144 14596 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 4816 11104 7113 11132
rect 4816 11076 4844 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11101 7343 11135
rect 7650 11132 7656 11144
rect 7563 11104 7656 11132
rect 7285 11095 7343 11101
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 4798 11064 4804 11076
rect 4540 11036 4804 11064
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 6641 11067 6699 11073
rect 5368 11036 5672 11064
rect 2866 10996 2872 11008
rect 2827 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5368 10996 5396 11036
rect 5534 10996 5540 11008
rect 5132 10968 5396 10996
rect 5495 10968 5540 10996
rect 5132 10956 5138 10968
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 5644 10996 5672 11036
rect 6641 11033 6653 11067
rect 6687 11064 6699 11067
rect 6822 11064 6828 11076
rect 6687 11036 6828 11064
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 7098 10996 7104 11008
rect 5644 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7668 10996 7696 11092
rect 10244 11064 10272 11095
rect 11606 11064 11612 11076
rect 8588 11036 10272 11064
rect 11567 11036 11612 11064
rect 8588 10996 8616 11036
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12452 11064 12480 11095
rect 12124 11036 12480 11064
rect 12124 11024 12130 11036
rect 12710 11024 12716 11076
rect 12768 11064 12774 11076
rect 12897 11067 12955 11073
rect 12897 11064 12909 11067
rect 12768 11036 12909 11064
rect 12768 11024 12774 11036
rect 12897 11033 12909 11036
rect 12943 11064 12955 11067
rect 13556 11064 13584 11095
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 14608 11104 15853 11132
rect 14608 11092 14614 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11132 18475 11135
rect 19426 11132 19432 11144
rect 18463 11104 19432 11132
rect 18463 11101 18475 11104
rect 18417 11095 18475 11101
rect 17586 11064 17592 11076
rect 12943 11036 13584 11064
rect 17547 11036 17592 11064
rect 12943 11033 12955 11036
rect 12897 11027 12955 11033
rect 17586 11024 17592 11036
rect 17644 11064 17650 11076
rect 18248 11064 18276 11095
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 17644 11036 18276 11064
rect 17644 11024 17650 11036
rect 7668 10968 8616 10996
rect 12158 10956 12164 11008
rect 12216 10996 12222 11008
rect 15378 10996 15384 11008
rect 12216 10968 15384 10996
rect 12216 10956 12222 10968
rect 15378 10956 15384 10968
rect 15436 10956 15442 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 1728 10764 2053 10792
rect 1728 10752 1734 10764
rect 2041 10761 2053 10764
rect 2087 10761 2099 10795
rect 2041 10755 2099 10761
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 3384 10764 4077 10792
rect 3384 10752 3390 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 8478 10792 8484 10804
rect 4065 10755 4123 10761
rect 4172 10764 8340 10792
rect 8439 10764 8484 10792
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 4172 10724 4200 10764
rect 3844 10696 4200 10724
rect 3844 10684 3850 10696
rect 7926 10684 7932 10736
rect 7984 10724 7990 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7984 10696 8217 10724
rect 7984 10684 7990 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8312 10724 8340 10764
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 12066 10792 12072 10804
rect 8588 10764 11928 10792
rect 12027 10764 12072 10792
rect 8588 10724 8616 10764
rect 8312 10696 8616 10724
rect 11900 10724 11928 10764
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 12342 10752 12348 10804
rect 12400 10792 12406 10804
rect 14369 10795 14427 10801
rect 12400 10764 14044 10792
rect 12400 10752 12406 10764
rect 12253 10727 12311 10733
rect 12253 10724 12265 10727
rect 11900 10696 12265 10724
rect 8205 10687 8263 10693
rect 12253 10693 12265 10696
rect 12299 10693 12311 10727
rect 12253 10687 12311 10693
rect 2682 10656 2688 10668
rect 2643 10628 2688 10656
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3694 10656 3700 10668
rect 3655 10628 3700 10656
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 5592 10628 6837 10656
rect 5592 10616 5598 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 8220 10656 8248 10687
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8220 10628 9045 10656
rect 6825 10619 6883 10625
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10686 10656 10692 10668
rect 10100 10628 10692 10656
rect 10100 10616 10106 10628
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 14016 10656 14044 10764
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 14550 10792 14556 10804
rect 14415 10764 14556 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 16482 10792 16488 10804
rect 16443 10764 16488 10792
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 15473 10727 15531 10733
rect 15473 10693 15485 10727
rect 15519 10724 15531 10727
rect 15519 10696 16988 10724
rect 15519 10693 15531 10696
rect 15473 10687 15531 10693
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 14016 10628 15945 10656
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 16114 10656 16120 10668
rect 16027 10628 16120 10656
rect 15933 10619 15991 10625
rect 16114 10616 16120 10628
rect 16172 10656 16178 10668
rect 16960 10665 16988 10696
rect 16945 10659 17003 10665
rect 16172 10628 16804 10656
rect 16172 10616 16178 10628
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2866 10588 2872 10600
rect 2547 10560 2872 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 4982 10588 4988 10600
rect 4571 10560 4988 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 8846 10588 8852 10600
rect 8807 10560 8852 10588
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 12158 10588 12164 10600
rect 8956 10560 12164 10588
rect 4062 10480 4068 10532
rect 4120 10520 4126 10532
rect 7098 10529 7104 10532
rect 7092 10520 7104 10529
rect 4120 10492 4568 10520
rect 7059 10492 7104 10520
rect 4120 10480 4126 10492
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2455 10424 3065 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3053 10415 3111 10421
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4430 10452 4436 10464
rect 3568 10424 3613 10452
rect 4391 10424 4436 10452
rect 3568 10412 3574 10424
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 4540 10452 4568 10492
rect 7092 10483 7104 10492
rect 7098 10480 7104 10483
rect 7156 10480 7162 10532
rect 8956 10520 8984 10560
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12768 10560 13001 10588
rect 12768 10548 12774 10560
rect 12989 10557 13001 10560
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 13078 10548 13084 10600
rect 13136 10588 13142 10600
rect 15654 10588 15660 10600
rect 13136 10560 15660 10588
rect 13136 10548 13142 10560
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 7208 10492 8984 10520
rect 10956 10523 11014 10529
rect 7208 10452 7236 10492
rect 10956 10489 10968 10523
rect 11002 10520 11014 10523
rect 11606 10520 11612 10532
rect 11002 10492 11612 10520
rect 11002 10489 11014 10492
rect 10956 10483 11014 10489
rect 11606 10480 11612 10492
rect 11664 10480 11670 10532
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 13256 10523 13314 10529
rect 12299 10492 12480 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 4540 10424 7236 10452
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 11974 10452 11980 10464
rect 8987 10424 11980 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12452 10452 12480 10492
rect 13256 10489 13268 10523
rect 13302 10520 13314 10523
rect 13354 10520 13360 10532
rect 13302 10492 13360 10520
rect 13302 10489 13314 10492
rect 13256 10483 13314 10489
rect 13354 10480 13360 10492
rect 13412 10480 13418 10532
rect 15841 10523 15899 10529
rect 15841 10520 15853 10523
rect 13455 10492 15853 10520
rect 13455 10452 13483 10492
rect 15841 10489 15853 10492
rect 15887 10489 15899 10523
rect 16776 10520 16804 10628
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 17034 10616 17040 10668
rect 17092 10656 17098 10668
rect 17092 10628 17137 10656
rect 17092 10616 17098 10628
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 18012 10628 18061 10656
rect 18012 10616 18018 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 18316 10591 18374 10597
rect 18316 10557 18328 10591
rect 18362 10588 18374 10591
rect 19150 10588 19156 10600
rect 18362 10560 19156 10588
rect 18362 10557 18374 10560
rect 18316 10551 18374 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 16776 10492 19472 10520
rect 15841 10483 15899 10489
rect 16850 10452 16856 10464
rect 12452 10424 13483 10452
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 19444 10461 19472 10492
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10421 19487 10455
rect 19429 10415 19487 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 13078 10248 13084 10260
rect 4028 10220 13084 10248
rect 4028 10208 4034 10220
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13354 10248 13360 10260
rect 13267 10220 13360 10248
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 13722 10248 13728 10260
rect 13679 10220 13728 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 2032 10183 2090 10189
rect 2032 10149 2044 10183
rect 2078 10180 2090 10183
rect 3694 10180 3700 10192
rect 2078 10152 3700 10180
rect 2078 10149 2090 10152
rect 2032 10143 2090 10149
rect 3694 10140 3700 10152
rect 3752 10140 3758 10192
rect 4430 10140 4436 10192
rect 4488 10180 4494 10192
rect 4982 10180 4988 10192
rect 4488 10152 4988 10180
rect 4488 10140 4494 10152
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 5736 10152 6776 10180
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 2314 10112 2320 10124
rect 1811 10084 2320 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 2314 10072 2320 10084
rect 2372 10112 2378 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 2372 10084 4077 10112
rect 2372 10072 2378 10084
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 4332 10115 4390 10121
rect 4332 10081 4344 10115
rect 4378 10112 4390 10115
rect 4706 10112 4712 10124
rect 4378 10084 4712 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 4706 10072 4712 10084
rect 4764 10112 4770 10124
rect 5736 10121 5764 10152
rect 5994 10121 6000 10124
rect 5721 10115 5779 10121
rect 4764 10084 5120 10112
rect 4764 10072 4770 10084
rect 5092 9988 5120 10084
rect 5721 10081 5733 10115
rect 5767 10081 5779 10115
rect 5988 10112 6000 10121
rect 5955 10084 6000 10112
rect 5721 10075 5779 10081
rect 5988 10075 6000 10084
rect 5994 10072 6000 10075
rect 6052 10072 6058 10124
rect 6748 10044 6776 10152
rect 6914 10140 6920 10192
rect 6972 10180 6978 10192
rect 8297 10183 8355 10189
rect 6972 10152 7880 10180
rect 6972 10140 6978 10152
rect 7852 10121 7880 10152
rect 8297 10149 8309 10183
rect 8343 10180 8355 10183
rect 9674 10180 9680 10192
rect 8343 10152 9680 10180
rect 8343 10149 8355 10152
rect 8297 10143 8355 10149
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 12066 10140 12072 10192
rect 12124 10180 12130 10192
rect 12222 10183 12280 10189
rect 12222 10180 12234 10183
rect 12124 10152 12234 10180
rect 12124 10140 12130 10152
rect 12222 10149 12234 10152
rect 12268 10149 12280 10183
rect 13372 10180 13400 10208
rect 13372 10152 14228 10180
rect 12222 10143 12280 10149
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 10318 10112 10324 10124
rect 8435 10084 10324 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 10744 10084 11989 10112
rect 10744 10072 10750 10084
rect 11977 10081 11989 10084
rect 12023 10112 12035 10115
rect 12710 10112 12716 10124
rect 12023 10084 12716 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 13998 10112 14004 10124
rect 13959 10084 14004 10112
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 7650 10044 7656 10056
rect 6748 10016 7656 10044
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 14200 10053 14228 10152
rect 16206 10112 16212 10124
rect 16167 10084 16212 10112
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 16476 10115 16534 10121
rect 16476 10081 16488 10115
rect 16522 10112 16534 10115
rect 17034 10112 17040 10124
rect 16522 10084 17040 10112
rect 16522 10081 16534 10084
rect 16476 10075 16534 10081
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13320 10016 14105 10044
rect 13320 10004 13326 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14185 10047 14243 10053
rect 14185 10013 14197 10047
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 5074 9936 5080 9988
rect 5132 9976 5138 9988
rect 5132 9948 5580 9976
rect 5132 9936 5138 9948
rect 2682 9868 2688 9920
rect 2740 9908 2746 9920
rect 3145 9911 3203 9917
rect 3145 9908 3157 9911
rect 2740 9880 3157 9908
rect 2740 9868 2746 9880
rect 3145 9877 3157 9880
rect 3191 9877 3203 9911
rect 3145 9871 3203 9877
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 3752 9880 5457 9908
rect 3752 9868 3758 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 5552 9908 5580 9948
rect 6656 9948 8064 9976
rect 6656 9908 6684 9948
rect 7098 9908 7104 9920
rect 5552 9880 6684 9908
rect 7059 9880 7104 9908
rect 5445 9871 5503 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 7650 9908 7656 9920
rect 7611 9880 7656 9908
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 7926 9908 7932 9920
rect 7887 9880 7932 9908
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8036 9908 8064 9948
rect 13280 9948 13492 9976
rect 13280 9908 13308 9948
rect 8036 9880 13308 9908
rect 13464 9908 13492 9948
rect 17589 9911 17647 9917
rect 17589 9908 17601 9911
rect 13464 9880 17601 9908
rect 17589 9877 17601 9880
rect 17635 9877 17647 9911
rect 17589 9871 17647 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 3145 9707 3203 9713
rect 3145 9673 3157 9707
rect 3191 9704 3203 9707
rect 3510 9704 3516 9716
rect 3191 9676 3516 9704
rect 3191 9673 3203 9676
rect 3145 9667 3203 9673
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6052 9676 7512 9704
rect 6052 9664 6058 9676
rect 4154 9636 4160 9648
rect 4115 9608 4160 9636
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 4304 9608 5733 9636
rect 4304 9596 4310 9608
rect 5721 9605 5733 9608
rect 5767 9605 5779 9639
rect 5721 9599 5779 9605
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 3835 9540 4813 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 4801 9537 4813 9540
rect 4847 9568 4859 9571
rect 5074 9568 5080 9580
rect 4847 9540 5080 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 7098 9568 7104 9580
rect 6411 9540 7104 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7484 9577 7512 9676
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 17034 9704 17040 9716
rect 8628 9676 9628 9704
rect 16995 9676 17040 9704
rect 8628 9664 8634 9676
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 8588 9568 8616 9664
rect 9600 9636 9628 9676
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 10045 9639 10103 9645
rect 10045 9636 10057 9639
rect 9600 9608 10057 9636
rect 10045 9605 10057 9608
rect 10091 9605 10103 9639
rect 10318 9636 10324 9648
rect 10279 9608 10324 9636
rect 10045 9599 10103 9605
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 10870 9568 10876 9580
rect 7515 9540 8616 9568
rect 10831 9540 10876 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9568 13415 9571
rect 13998 9568 14004 9580
rect 13403 9540 14004 9568
rect 13403 9537 13415 9540
rect 13357 9531 13415 9537
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 16908 9540 17325 9568
rect 16908 9528 16914 9540
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 4706 9500 4712 9512
rect 4264 9472 4712 9500
rect 4264 9444 4292 9472
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 7926 9500 7932 9512
rect 6227 9472 7932 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 8932 9503 8990 9509
rect 8932 9469 8944 9503
rect 8978 9500 8990 9503
rect 10888 9500 10916 9528
rect 8978 9472 10916 9500
rect 15657 9503 15715 9509
rect 8978 9469 8990 9472
rect 8932 9463 8990 9469
rect 15657 9469 15669 9503
rect 15703 9500 15715 9503
rect 16206 9500 16212 9512
rect 15703 9472 16212 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 3513 9435 3571 9441
rect 3513 9401 3525 9435
rect 3559 9432 3571 9435
rect 4246 9432 4252 9444
rect 3559 9404 4252 9432
rect 3559 9401 3571 9404
rect 3513 9395 3571 9401
rect 4246 9392 4252 9404
rect 4304 9392 4310 9444
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9432 4583 9435
rect 5994 9432 6000 9444
rect 4571 9404 6000 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 6135 9404 6868 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 4154 9364 4160 9376
rect 3651 9336 4160 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 5810 9364 5816 9376
rect 4663 9336 5816 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 5810 9324 5816 9336
rect 5868 9364 5874 9376
rect 6178 9364 6184 9376
rect 5868 9336 6184 9364
rect 5868 9324 5874 9336
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6840 9373 6868 9404
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7064 9404 7328 9432
rect 7064 9392 7070 9404
rect 7300 9376 7328 9404
rect 7650 9392 7656 9444
rect 7708 9432 7714 9444
rect 8680 9432 8708 9463
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 7708 9404 8708 9432
rect 10781 9435 10839 9441
rect 7708 9392 7714 9404
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 12250 9432 12256 9444
rect 10827 9404 12256 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 12342 9392 12348 9444
rect 12400 9432 12406 9444
rect 15924 9435 15982 9441
rect 12400 9404 15516 9432
rect 12400 9392 12406 9404
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9333 6883 9367
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 6825 9327 6883 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7340 9336 7385 9364
rect 7340 9324 7346 9336
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 7524 9336 10701 9364
rect 7524 9324 7530 9336
rect 10689 9333 10701 9336
rect 10735 9333 10747 9367
rect 15488 9364 15516 9404
rect 15924 9401 15936 9435
rect 15970 9432 15982 9435
rect 16114 9432 16120 9444
rect 15970 9404 16120 9432
rect 15970 9401 15982 9404
rect 15924 9395 15982 9401
rect 16114 9392 16120 9404
rect 16172 9392 16178 9444
rect 18506 9364 18512 9376
rect 15488 9336 18512 9364
rect 10689 9327 10747 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2038 9160 2044 9172
rect 1995 9132 2044 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 4890 9160 4896 9172
rect 4755 9132 4896 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 4890 9120 4896 9132
rect 4948 9160 4954 9172
rect 5261 9163 5319 9169
rect 5261 9160 5273 9163
rect 4948 9132 5273 9160
rect 4948 9120 4954 9132
rect 5261 9129 5273 9132
rect 5307 9129 5319 9163
rect 5261 9123 5319 9129
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 7190 9160 7196 9172
rect 6411 9132 7196 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 12342 9092 12348 9104
rect 4120 9064 12348 9092
rect 4120 9052 4126 9064
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 1765 9027 1823 9033
rect 1765 9024 1777 9027
rect 1728 8996 1777 9024
rect 1728 8984 1734 8996
rect 1765 8993 1777 8996
rect 1811 8993 1823 9027
rect 1765 8987 1823 8993
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 3660 8996 5181 9024
rect 3660 8984 3666 8996
rect 5169 8993 5181 8996
rect 5215 9024 5227 9027
rect 5718 9024 5724 9036
rect 5215 8996 5724 9024
rect 5215 8993 5227 8996
rect 5169 8987 5227 8993
rect 5718 8984 5724 8996
rect 5776 9024 5782 9036
rect 7466 9024 7472 9036
rect 5776 8996 7472 9024
rect 5776 8984 5782 8996
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8185 9027 8243 9033
rect 8185 9024 8197 9027
rect 7892 8996 8197 9024
rect 7892 8984 7898 8996
rect 8185 8993 8197 8996
rect 8231 8993 8243 9027
rect 8185 8987 8243 8993
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 8812 8996 10057 9024
rect 8812 8984 8818 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4890 8956 4896 8968
rect 4212 8928 4896 8956
rect 4212 8916 4218 8928
rect 4890 8916 4896 8928
rect 4948 8956 4954 8968
rect 5074 8956 5080 8968
rect 4948 8928 5080 8956
rect 4948 8916 4954 8928
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5350 8956 5356 8968
rect 5311 8928 5356 8956
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7650 8956 7656 8968
rect 7248 8928 7656 8956
rect 7248 8916 7254 8928
rect 7650 8916 7656 8928
rect 7708 8956 7714 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 7708 8928 7941 8956
rect 7708 8916 7714 8928
rect 7929 8925 7941 8928
rect 7975 8925 7987 8959
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 7929 8919 7987 8925
rect 8956 8928 10149 8956
rect 4798 8820 4804 8832
rect 4759 8792 4804 8820
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 8956 8820 8984 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10870 8956 10876 8968
rect 10367 8928 10876 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 9309 8891 9367 8897
rect 9309 8857 9321 8891
rect 9355 8888 9367 8891
rect 10336 8888 10364 8919
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 9355 8860 10364 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 5960 8792 8984 8820
rect 5960 8780 5966 8792
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 7892 8588 8585 8616
rect 7892 8576 7898 8588
rect 8573 8585 8585 8588
rect 8619 8585 8631 8619
rect 8573 8579 8631 8585
rect 3510 8508 3516 8560
rect 3568 8548 3574 8560
rect 5350 8548 5356 8560
rect 3568 8520 5356 8548
rect 3568 8508 3574 8520
rect 5350 8508 5356 8520
rect 5408 8548 5414 8560
rect 5408 8520 5764 8548
rect 5408 8508 5414 8520
rect 1670 8480 1676 8492
rect 1631 8452 1676 8480
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 4706 8480 4712 8492
rect 4667 8452 4712 8480
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5736 8489 5764 8520
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 7190 8480 7196 8492
rect 7151 8452 7196 8480
rect 5721 8443 5779 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9180 8452 9413 8480
rect 9180 8440 9186 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 2130 8412 2136 8424
rect 2091 8384 2136 8412
rect 1397 8375 1455 8381
rect 1412 8344 1440 8375
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2400 8415 2458 8421
rect 2400 8381 2412 8415
rect 2446 8412 2458 8415
rect 2682 8412 2688 8424
rect 2446 8384 2688 8412
rect 2446 8381 2458 8384
rect 2400 8375 2458 8381
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8412 4675 8415
rect 4798 8412 4804 8424
rect 4663 8384 4804 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 8754 8412 8760 8424
rect 5552 8384 8760 8412
rect 5552 8356 5580 8384
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 8904 8384 9229 8412
rect 8904 8372 8910 8384
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 11698 8412 11704 8424
rect 9355 8384 11704 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 4525 8347 4583 8353
rect 1412 8316 4476 8344
rect 3510 8276 3516 8288
rect 3471 8248 3516 8276
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 4154 8276 4160 8288
rect 4115 8248 4160 8276
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 4448 8276 4476 8316
rect 4525 8313 4537 8347
rect 4571 8344 4583 8347
rect 5534 8344 5540 8356
rect 4571 8316 5212 8344
rect 5495 8316 5540 8344
rect 4571 8313 4583 8316
rect 4525 8307 4583 8313
rect 4798 8276 4804 8288
rect 4448 8248 4804 8276
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 5184 8285 5212 8316
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5629 8347 5687 8353
rect 5629 8313 5641 8347
rect 5675 8344 5687 8347
rect 5718 8344 5724 8356
rect 5675 8316 5724 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 7460 8347 7518 8353
rect 7460 8313 7472 8347
rect 7506 8344 7518 8347
rect 8202 8344 8208 8356
rect 7506 8316 8208 8344
rect 7506 8313 7518 8316
rect 7460 8307 7518 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 5169 8279 5227 8285
rect 5169 8245 5181 8279
rect 5215 8245 5227 8279
rect 8846 8276 8852 8288
rect 8807 8248 8852 8276
rect 5169 8239 5227 8245
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 9398 8236 9404 8288
rect 9456 8276 9462 8288
rect 17586 8276 17592 8288
rect 9456 8248 17592 8276
rect 9456 8236 9462 8248
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1544 8044 1777 8072
rect 1544 8032 1550 8044
rect 1765 8041 1777 8044
rect 1811 8041 1823 8075
rect 1765 8035 1823 8041
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 4212 8044 4537 8072
rect 4212 8032 4218 8044
rect 4525 8041 4537 8044
rect 4571 8041 4583 8075
rect 4525 8035 4583 8041
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 8754 8072 8760 8084
rect 4948 8044 8760 8072
rect 4948 8032 4954 8044
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8904 8044 8953 8072
rect 8904 8032 8910 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 18601 8075 18659 8081
rect 18601 8041 18613 8075
rect 18647 8072 18659 8075
rect 19702 8072 19708 8084
rect 18647 8044 19708 8072
rect 18647 8041 18659 8044
rect 18601 8035 18659 8041
rect 19702 8032 19708 8044
rect 19760 8032 19766 8084
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 9398 8004 9404 8016
rect 4120 7976 9404 8004
rect 4120 7964 4126 7976
rect 9398 7964 9404 7976
rect 9456 7964 9462 8016
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 2041 7939 2099 7945
rect 2041 7905 2053 7939
rect 2087 7936 2099 7939
rect 2143 7939 2201 7945
rect 2143 7936 2155 7939
rect 2087 7908 2155 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 2143 7905 2155 7908
rect 2189 7905 2201 7939
rect 2143 7899 2201 7905
rect 1596 7868 1624 7899
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4212 7908 4445 7936
rect 4212 7896 4218 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 5436 7939 5494 7945
rect 5436 7936 5448 7939
rect 4433 7899 4491 7905
rect 4724 7908 5448 7936
rect 4724 7877 4752 7908
rect 5436 7905 5448 7908
rect 5482 7936 5494 7939
rect 5994 7936 6000 7948
rect 5482 7908 6000 7936
rect 5482 7905 5494 7908
rect 5436 7899 5494 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 7092 7939 7150 7945
rect 7092 7936 7104 7939
rect 6748 7908 7104 7936
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1596 7840 2329 7868
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 5166 7868 5172 7880
rect 5127 7840 5172 7868
rect 4709 7831 4767 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 6549 7803 6607 7809
rect 6549 7769 6561 7803
rect 6595 7800 6607 7803
rect 6748 7800 6776 7908
rect 7092 7905 7104 7908
rect 7138 7936 7150 7939
rect 8846 7936 8852 7948
rect 7138 7908 8156 7936
rect 8807 7908 8852 7936
rect 7138 7905 7150 7908
rect 7092 7899 7150 7905
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6595 7772 6776 7800
rect 6595 7769 6607 7772
rect 6549 7763 6607 7769
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 2087 7704 4077 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 6730 7732 6736 7744
rect 4304 7704 6736 7732
rect 4304 7692 4310 7704
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 6840 7732 6868 7831
rect 8128 7800 8156 7908
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 18417 7939 18475 7945
rect 18417 7936 18429 7939
rect 8996 7908 18429 7936
rect 8996 7896 9002 7908
rect 18417 7905 18429 7908
rect 18463 7905 18475 7939
rect 18417 7899 18475 7905
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8260 7840 9045 7868
rect 8260 7828 8266 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 9122 7800 9128 7812
rect 8128 7772 9128 7800
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 7190 7732 7196 7744
rect 6840 7704 7196 7732
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 8202 7732 8208 7744
rect 8163 7704 8208 7732
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8478 7732 8484 7744
rect 8439 7704 8484 7732
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5994 7528 6000 7540
rect 4120 7500 5580 7528
rect 5955 7500 6000 7528
rect 4120 7488 4126 7500
rect 5552 7460 5580 7500
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 6788 7500 8401 7528
rect 6788 7488 6794 7500
rect 8389 7497 8401 7500
rect 8435 7497 8447 7531
rect 8389 7491 8447 7497
rect 19153 7531 19211 7537
rect 19153 7497 19165 7531
rect 19199 7528 19211 7531
rect 19334 7528 19340 7540
rect 19199 7500 19340 7528
rect 19199 7497 19211 7500
rect 19153 7491 19211 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 8938 7460 8944 7472
rect 5552 7432 8944 7460
rect 8938 7420 8944 7432
rect 8996 7420 9002 7472
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8202 7392 8208 7404
rect 8159 7364 8208 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 9122 7392 9128 7404
rect 9083 7364 9128 7392
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 2130 7284 2136 7336
rect 2188 7324 2194 7336
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2188 7296 2973 7324
rect 2188 7284 2194 7296
rect 2961 7293 2973 7296
rect 3007 7324 3019 7327
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 3007 7296 4629 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 4617 7293 4629 7296
rect 4663 7324 4675 7327
rect 5166 7324 5172 7336
rect 4663 7296 5172 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 6086 7324 6092 7336
rect 5552 7296 6092 7324
rect 5552 7268 5580 7296
rect 6086 7284 6092 7296
rect 6144 7324 6150 7336
rect 8662 7324 8668 7336
rect 6144 7296 8668 7324
rect 6144 7284 6150 7296
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8812 7296 8953 7324
rect 8812 7284 8818 7296
rect 8941 7293 8953 7296
rect 8987 7293 8999 7327
rect 18966 7324 18972 7336
rect 18927 7296 18972 7324
rect 8941 7287 8999 7293
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 3228 7259 3286 7265
rect 3228 7225 3240 7259
rect 3274 7256 3286 7259
rect 3510 7256 3516 7268
rect 3274 7228 3516 7256
rect 3274 7225 3286 7228
rect 3228 7219 3286 7225
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 4706 7256 4712 7268
rect 4356 7228 4712 7256
rect 4356 7197 4384 7228
rect 4706 7216 4712 7228
rect 4764 7256 4770 7268
rect 4862 7259 4920 7265
rect 4862 7256 4874 7259
rect 4764 7228 4874 7256
rect 4764 7216 4770 7228
rect 4862 7225 4874 7228
rect 4908 7225 4920 7259
rect 4862 7219 4920 7225
rect 5534 7216 5540 7268
rect 5592 7216 5598 7268
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7256 7067 7259
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7055 7228 7849 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 7837 7225 7849 7228
rect 7883 7225 7895 7259
rect 7837 7219 7895 7225
rect 8389 7259 8447 7265
rect 8389 7225 8401 7259
rect 8435 7256 8447 7259
rect 8849 7259 8907 7265
rect 8849 7256 8861 7259
rect 8435 7228 8861 7256
rect 8435 7225 8447 7228
rect 8389 7219 8447 7225
rect 8849 7225 8861 7228
rect 8895 7225 8907 7259
rect 8849 7219 8907 7225
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7157 4399 7191
rect 4341 7151 4399 7157
rect 7469 7191 7527 7197
rect 7469 7157 7481 7191
rect 7515 7188 7527 7191
rect 7558 7188 7564 7200
rect 7515 7160 7564 7188
rect 7515 7157 7527 7160
rect 7469 7151 7527 7157
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 7929 7191 7987 7197
rect 7929 7157 7941 7191
rect 7975 7188 7987 7191
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 7975 7160 8493 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 8481 7157 8493 7160
rect 8527 7157 8539 7191
rect 8481 7151 8539 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 7558 6984 7564 6996
rect 7519 6956 7564 6984
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 8297 6987 8355 6993
rect 8297 6953 8309 6987
rect 8343 6984 8355 6987
rect 8846 6984 8852 6996
rect 8343 6956 8852 6984
rect 8343 6953 8355 6956
rect 8297 6947 8355 6953
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 18966 6916 18972 6928
rect 4120 6888 18972 6916
rect 4120 6876 4126 6888
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 4479 6820 5089 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 8478 6848 8484 6860
rect 7699 6820 8484 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 8662 6848 8668 6860
rect 8623 6820 8668 6848
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 19242 6808 19248 6860
rect 19300 6848 19306 6860
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 19300 6820 19441 6848
rect 19300 6808 19306 6820
rect 19429 6817 19441 6820
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 3936 6752 4537 6780
rect 3936 6740 3942 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4525 6743 4583 6749
rect 4065 6715 4123 6721
rect 4065 6681 4077 6715
rect 4111 6712 4123 6715
rect 4154 6712 4160 6724
rect 4111 6684 4160 6712
rect 4111 6681 4123 6684
rect 4065 6675 4123 6681
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 4540 6712 4568 6743
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 7742 6780 7748 6792
rect 7703 6752 7748 6780
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8754 6780 8760 6792
rect 8715 6752 8760 6780
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6780 8999 6783
rect 9122 6780 9128 6792
rect 8987 6752 9128 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9674 6780 9680 6792
rect 9272 6752 9680 6780
rect 9272 6740 9278 6752
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 7282 6712 7288 6724
rect 4540 6684 7288 6712
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 19610 6712 19616 6724
rect 19571 6684 19616 6712
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 7193 6647 7251 6653
rect 7193 6644 7205 6647
rect 4856 6616 7205 6644
rect 4856 6604 4862 6616
rect 7193 6613 7205 6616
rect 7239 6613 7251 6647
rect 7193 6607 7251 6613
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 19242 6644 19248 6656
rect 9732 6616 19248 6644
rect 9732 6604 9738 6616
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 6178 6440 6184 6452
rect 5868 6412 6184 6440
rect 5868 6400 5874 6412
rect 6178 6400 6184 6412
rect 6236 6440 6242 6452
rect 8754 6440 8760 6452
rect 6236 6412 8760 6440
rect 6236 6400 6242 6412
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 20073 6443 20131 6449
rect 20073 6409 20085 6443
rect 20119 6440 20131 6443
rect 20990 6440 20996 6452
rect 20119 6412 20996 6440
rect 20119 6409 20131 6412
rect 20073 6403 20131 6409
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 19889 6239 19947 6245
rect 19889 6236 19901 6239
rect 4028 6208 19901 6236
rect 4028 6196 4034 6208
rect 19889 6205 19901 6208
rect 19935 6205 19947 6239
rect 19889 6199 19947 6205
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 20441 5899 20499 5905
rect 20441 5865 20453 5899
rect 20487 5896 20499 5899
rect 20806 5896 20812 5908
rect 20487 5868 20812 5896
rect 20487 5865 20499 5868
rect 20441 5859 20499 5865
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 4120 5732 20269 5760
rect 4120 5720 4126 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 20898 5352 20904 5364
rect 20763 5324 20904 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 4120 5120 20545 5148
rect 4120 5108 4126 5120
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4890 4128 4896 4140
rect 4028 4100 4896 4128
rect 4028 4088 4034 4100
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 5626 2564 5632 2576
rect 2832 2536 5632 2564
rect 2832 2524 2838 2536
rect 5626 2524 5632 2536
rect 5684 2524 5690 2576
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 3694 1980 3700 2032
rect 3752 2020 3758 2032
rect 5534 2020 5540 2032
rect 3752 1992 5540 2020
rect 3752 1980 3758 1992
rect 5534 1980 5540 1992
rect 5592 1980 5598 2032
rect 3694 1708 3700 1760
rect 3752 1748 3758 1760
rect 5718 1748 5724 1760
rect 3752 1720 5724 1748
rect 3752 1708 3758 1720
rect 5718 1708 5724 1720
rect 5776 1708 5782 1760
rect 4062 1028 4068 1080
rect 4120 1068 4126 1080
rect 5810 1068 5816 1080
rect 4120 1040 5816 1068
rect 4120 1028 4126 1040
rect 5810 1028 5816 1040
rect 5868 1028 5874 1080
rect 3234 416 3240 468
rect 3292 456 3298 468
rect 4982 456 4988 468
rect 3292 428 4988 456
rect 3292 416 3298 428
rect 4982 416 4988 428
rect 5040 416 5046 468
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2872 20000 2924 20052
rect 5632 20000 5684 20052
rect 9312 20000 9364 20052
rect 12900 20000 12952 20052
rect 13360 20000 13412 20052
rect 15200 20000 15252 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 16120 20000 16172 20052
rect 16580 20000 16632 20052
rect 17040 20000 17092 20052
rect 17500 20000 17552 20052
rect 18420 20000 18472 20052
rect 18880 20000 18932 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 6000 19864 6052 19916
rect 9680 19864 9732 19916
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 12992 19864 13044 19916
rect 13360 19907 13412 19916
rect 13360 19873 13369 19907
rect 13369 19873 13403 19907
rect 13403 19873 13412 19907
rect 13360 19864 13412 19873
rect 14372 19864 14424 19916
rect 15200 19864 15252 19916
rect 16120 19864 16172 19916
rect 16580 19907 16632 19916
rect 16580 19873 16589 19907
rect 16589 19873 16623 19907
rect 16623 19873 16632 19907
rect 16580 19864 16632 19873
rect 17132 19907 17184 19916
rect 17132 19873 17141 19907
rect 17141 19873 17175 19907
rect 17175 19873 17184 19907
rect 17132 19864 17184 19873
rect 17960 19864 18012 19916
rect 18512 19864 18564 19916
rect 18880 19907 18932 19916
rect 18880 19873 18889 19907
rect 18889 19873 18923 19907
rect 18923 19873 18932 19907
rect 18880 19864 18932 19873
rect 4896 19796 4948 19848
rect 5908 19839 5960 19848
rect 5908 19805 5917 19839
rect 5917 19805 5951 19839
rect 5951 19805 5960 19839
rect 5908 19796 5960 19805
rect 9956 19796 10008 19848
rect 10416 19839 10468 19848
rect 2780 19728 2832 19780
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 14280 19728 14332 19780
rect 2228 19660 2280 19712
rect 9772 19703 9824 19712
rect 9772 19669 9781 19703
rect 9781 19669 9815 19703
rect 9815 19669 9824 19703
rect 9772 19660 9824 19669
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3424 19456 3476 19508
rect 1768 19320 1820 19372
rect 17868 19388 17920 19440
rect 18052 19388 18104 19440
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 2872 19252 2924 19304
rect 4344 19252 4396 19304
rect 4804 19252 4856 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 9956 19320 10008 19372
rect 12992 19363 13044 19372
rect 7380 19252 7432 19304
rect 204 19184 256 19236
rect 3148 19184 3200 19236
rect 5908 19184 5960 19236
rect 6828 19184 6880 19236
rect 7288 19184 7340 19236
rect 9680 19252 9732 19304
rect 10048 19295 10100 19304
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 14372 19320 14424 19372
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 17132 19320 17184 19372
rect 18512 19320 18564 19372
rect 10324 19295 10376 19304
rect 10324 19261 10358 19295
rect 10358 19261 10376 19295
rect 10324 19252 10376 19261
rect 12164 19252 12216 19304
rect 13176 19252 13228 19304
rect 13728 19252 13780 19304
rect 14096 19252 14148 19304
rect 15200 19252 15252 19304
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 15752 19252 15804 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 18696 19252 18748 19304
rect 19064 19252 19116 19304
rect 22100 19252 22152 19304
rect 8760 19184 8812 19236
rect 2964 19116 3016 19168
rect 4252 19116 4304 19168
rect 4896 19116 4948 19168
rect 8208 19116 8260 19168
rect 9220 19116 9272 19168
rect 13912 19184 13964 19236
rect 20628 19227 20680 19236
rect 20628 19193 20637 19227
rect 20637 19193 20671 19227
rect 20671 19193 20680 19227
rect 20628 19184 20680 19193
rect 10416 19116 10468 19168
rect 13820 19116 13872 19168
rect 15016 19116 15068 19168
rect 18052 19116 18104 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 1032 18844 1084 18896
rect 2320 18844 2372 18896
rect 1952 18819 2004 18828
rect 1952 18785 1961 18819
rect 1961 18785 1995 18819
rect 1995 18785 2004 18819
rect 1952 18776 2004 18785
rect 2044 18708 2096 18760
rect 2136 18572 2188 18624
rect 4436 18955 4488 18964
rect 4436 18921 4445 18955
rect 4445 18921 4479 18955
rect 4479 18921 4488 18955
rect 4436 18912 4488 18921
rect 5172 18912 5224 18964
rect 6828 18955 6880 18964
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 3148 18844 3200 18896
rect 3332 18819 3384 18828
rect 3332 18785 3341 18819
rect 3341 18785 3375 18819
rect 3375 18785 3384 18819
rect 3332 18776 3384 18785
rect 5908 18844 5960 18896
rect 7104 18844 7156 18896
rect 9772 18776 9824 18828
rect 10416 18819 10468 18828
rect 10416 18785 10450 18819
rect 10450 18785 10468 18819
rect 10416 18776 10468 18785
rect 10784 18776 10836 18828
rect 3516 18751 3568 18760
rect 3516 18717 3525 18751
rect 3525 18717 3559 18751
rect 3559 18717 3568 18751
rect 3516 18708 3568 18717
rect 4252 18708 4304 18760
rect 5080 18708 5132 18760
rect 8116 18751 8168 18760
rect 8116 18717 8125 18751
rect 8125 18717 8159 18751
rect 8159 18717 8168 18751
rect 8116 18708 8168 18717
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 8484 18708 8536 18760
rect 10048 18708 10100 18760
rect 3792 18640 3844 18692
rect 4988 18640 5040 18692
rect 9220 18640 9272 18692
rect 11980 18844 12032 18896
rect 12164 18844 12216 18896
rect 13360 18912 13412 18964
rect 17960 18912 18012 18964
rect 13912 18844 13964 18896
rect 16580 18887 16632 18896
rect 16580 18853 16589 18887
rect 16589 18853 16623 18887
rect 16623 18853 16632 18887
rect 16580 18844 16632 18853
rect 17040 18844 17092 18896
rect 11796 18819 11848 18828
rect 11796 18785 11805 18819
rect 11805 18785 11839 18819
rect 11839 18785 11848 18819
rect 11796 18776 11848 18785
rect 12532 18819 12584 18828
rect 12532 18785 12541 18819
rect 12541 18785 12575 18819
rect 12575 18785 12584 18819
rect 12532 18776 12584 18785
rect 14004 18819 14056 18828
rect 14004 18785 14013 18819
rect 14013 18785 14047 18819
rect 14047 18785 14056 18819
rect 14004 18776 14056 18785
rect 14464 18776 14516 18828
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 16672 18776 16724 18828
rect 14556 18708 14608 18760
rect 15200 18708 15252 18760
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 16488 18708 16540 18760
rect 17960 18776 18012 18828
rect 19064 18887 19116 18896
rect 19064 18853 19073 18887
rect 19073 18853 19107 18887
rect 19107 18853 19116 18887
rect 19064 18844 19116 18853
rect 18880 18708 18932 18760
rect 20628 18640 20680 18692
rect 7104 18572 7156 18624
rect 8760 18572 8812 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18368 2004 18420
rect 8116 18368 8168 18420
rect 8668 18368 8720 18420
rect 9956 18368 10008 18420
rect 10324 18368 10376 18420
rect 15200 18411 15252 18420
rect 15200 18377 15209 18411
rect 15209 18377 15243 18411
rect 15243 18377 15252 18411
rect 15200 18368 15252 18377
rect 572 18300 624 18352
rect 2780 18300 2832 18352
rect 5724 18275 5776 18284
rect 2136 18207 2188 18216
rect 2136 18173 2145 18207
rect 2145 18173 2179 18207
rect 2179 18173 2188 18207
rect 2136 18164 2188 18173
rect 2872 18164 2924 18216
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 5908 18275 5960 18284
rect 5908 18241 5917 18275
rect 5917 18241 5951 18275
rect 5951 18241 5960 18275
rect 5908 18232 5960 18241
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 8944 18232 8996 18284
rect 15844 18275 15896 18284
rect 7104 18207 7156 18216
rect 1676 18096 1728 18148
rect 4252 18096 4304 18148
rect 7104 18173 7113 18207
rect 7113 18173 7147 18207
rect 7147 18173 7156 18207
rect 7104 18164 7156 18173
rect 8852 18164 8904 18216
rect 9680 18164 9732 18216
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 1768 18071 1820 18080
rect 1768 18037 1777 18071
rect 1777 18037 1811 18071
rect 1811 18037 1820 18071
rect 1768 18028 1820 18037
rect 3516 18028 3568 18080
rect 4436 18028 4488 18080
rect 9956 18096 10008 18148
rect 10324 18139 10376 18148
rect 10324 18105 10358 18139
rect 10358 18105 10376 18139
rect 10324 18096 10376 18105
rect 7748 18028 7800 18080
rect 8392 18028 8444 18080
rect 8576 18071 8628 18080
rect 8576 18037 8585 18071
rect 8585 18037 8619 18071
rect 8619 18037 8628 18071
rect 8576 18028 8628 18037
rect 8760 18028 8812 18080
rect 9036 18028 9088 18080
rect 10600 18028 10652 18080
rect 14372 18164 14424 18216
rect 15016 18207 15068 18216
rect 15016 18173 15025 18207
rect 15025 18173 15059 18207
rect 15059 18173 15068 18207
rect 15016 18164 15068 18173
rect 15936 18096 15988 18148
rect 16856 18096 16908 18148
rect 22560 18096 22612 18148
rect 13544 18028 13596 18080
rect 14556 18071 14608 18080
rect 14556 18037 14565 18071
rect 14565 18037 14599 18071
rect 14599 18037 14608 18071
rect 14556 18028 14608 18037
rect 15476 18028 15528 18080
rect 19616 18028 19668 18080
rect 20260 18028 20312 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 3056 17867 3108 17876
rect 3056 17833 3065 17867
rect 3065 17833 3099 17867
rect 3099 17833 3108 17867
rect 3056 17824 3108 17833
rect 3332 17824 3384 17876
rect 5908 17824 5960 17876
rect 15936 17824 15988 17876
rect 17960 17824 18012 17876
rect 9864 17756 9916 17808
rect 14556 17756 14608 17808
rect 2412 17688 2464 17740
rect 6184 17688 6236 17740
rect 7012 17731 7064 17740
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7012 17688 7064 17697
rect 5264 17620 5316 17672
rect 2872 17552 2924 17604
rect 6828 17620 6880 17672
rect 9772 17688 9824 17740
rect 15844 17731 15896 17740
rect 15844 17697 15878 17731
rect 15878 17697 15896 17731
rect 15844 17688 15896 17697
rect 19064 17688 19116 17740
rect 9864 17620 9916 17672
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 13360 17620 13412 17672
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 17960 17620 18012 17672
rect 18512 17620 18564 17672
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 3792 17484 3844 17536
rect 11152 17484 11204 17536
rect 12072 17484 12124 17536
rect 14464 17484 14516 17536
rect 14556 17484 14608 17536
rect 17868 17484 17920 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 5724 17280 5776 17332
rect 5264 17212 5316 17264
rect 8484 17280 8536 17332
rect 10324 17280 10376 17332
rect 11612 17280 11664 17332
rect 12256 17280 12308 17332
rect 12532 17280 12584 17332
rect 14004 17280 14056 17332
rect 15660 17280 15712 17332
rect 15936 17280 15988 17332
rect 17960 17280 18012 17332
rect 19340 17280 19392 17332
rect 19800 17280 19852 17332
rect 2872 17144 2924 17196
rect 6092 17187 6144 17196
rect 6092 17153 6101 17187
rect 6101 17153 6135 17187
rect 6135 17153 6144 17187
rect 6092 17144 6144 17153
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 7288 17144 7340 17196
rect 8392 17144 8444 17196
rect 3792 17076 3844 17128
rect 8024 17076 8076 17128
rect 8852 17076 8904 17128
rect 9496 17076 9548 17128
rect 11888 17144 11940 17196
rect 15660 17144 15712 17196
rect 15844 17144 15896 17196
rect 18604 17187 18656 17196
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 19064 17187 19116 17196
rect 19064 17153 19073 17187
rect 19073 17153 19107 17187
rect 19107 17153 19116 17187
rect 19064 17144 19116 17153
rect 3516 17008 3568 17060
rect 3884 17008 3936 17060
rect 9864 17051 9916 17060
rect 9864 17017 9898 17051
rect 9898 17017 9916 17051
rect 9864 17008 9916 17017
rect 10232 17008 10284 17060
rect 13360 17076 13412 17128
rect 16212 17076 16264 17128
rect 17868 17076 17920 17128
rect 20904 17076 20956 17128
rect 21640 17076 21692 17128
rect 18420 17051 18472 17060
rect 18420 17017 18429 17051
rect 18429 17017 18463 17051
rect 18463 17017 18472 17051
rect 18420 17008 18472 17017
rect 20720 17008 20772 17060
rect 20996 17008 21048 17060
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 4160 16940 4212 16992
rect 5908 16940 5960 16992
rect 6828 16940 6880 16992
rect 8208 16940 8260 16992
rect 9680 16940 9732 16992
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 13268 16940 13320 16992
rect 15844 16983 15896 16992
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 15844 16940 15896 16949
rect 16304 16940 16356 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1492 16643 1544 16652
rect 1492 16609 1501 16643
rect 1501 16609 1535 16643
rect 1535 16609 1544 16643
rect 1492 16600 1544 16609
rect 6184 16736 6236 16788
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 12900 16736 12952 16788
rect 16304 16779 16356 16788
rect 2412 16668 2464 16720
rect 7104 16668 7156 16720
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 4252 16600 4304 16652
rect 5816 16600 5868 16652
rect 7196 16600 7248 16652
rect 8208 16600 8260 16652
rect 12992 16668 13044 16720
rect 16304 16745 16313 16779
rect 16313 16745 16347 16779
rect 16347 16745 16356 16779
rect 16304 16736 16356 16745
rect 16764 16668 16816 16720
rect 18512 16736 18564 16788
rect 18604 16668 18656 16720
rect 3976 16532 4028 16584
rect 1676 16507 1728 16516
rect 1676 16473 1685 16507
rect 1685 16473 1719 16507
rect 1719 16473 1728 16507
rect 1676 16464 1728 16473
rect 2872 16464 2924 16516
rect 7288 16396 7340 16448
rect 8852 16464 8904 16516
rect 8300 16396 8352 16448
rect 10416 16396 10468 16448
rect 12440 16643 12492 16652
rect 12440 16609 12474 16643
rect 12474 16609 12492 16643
rect 11888 16439 11940 16448
rect 11888 16405 11897 16439
rect 11897 16405 11931 16439
rect 11931 16405 11940 16439
rect 11888 16396 11940 16405
rect 12440 16600 12492 16609
rect 12900 16600 12952 16652
rect 13544 16600 13596 16652
rect 14188 16643 14240 16652
rect 14188 16609 14197 16643
rect 14197 16609 14231 16643
rect 14231 16609 14240 16643
rect 14188 16600 14240 16609
rect 17224 16643 17276 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 17224 16609 17258 16643
rect 17258 16609 17276 16643
rect 17224 16600 17276 16609
rect 12900 16396 12952 16448
rect 13084 16396 13136 16448
rect 15568 16464 15620 16516
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 7380 16192 7432 16244
rect 10232 16235 10284 16244
rect 4896 16124 4948 16176
rect 8668 16124 8720 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 5816 16099 5868 16108
rect 4160 15988 4212 16040
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 7748 16056 7800 16108
rect 8208 16056 8260 16108
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 7104 15988 7156 16040
rect 2780 15920 2832 15972
rect 9864 15920 9916 15972
rect 10232 16201 10241 16235
rect 10241 16201 10275 16235
rect 10275 16201 10284 16235
rect 10232 16192 10284 16201
rect 12808 16192 12860 16244
rect 14188 16192 14240 16244
rect 17224 16192 17276 16244
rect 10416 15988 10468 16040
rect 11888 15988 11940 16040
rect 15016 16124 15068 16176
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 14372 16099 14424 16108
rect 14372 16065 14381 16099
rect 14381 16065 14415 16099
rect 14415 16065 14424 16099
rect 14372 16056 14424 16065
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 15568 16056 15620 16108
rect 16028 16099 16080 16108
rect 16028 16065 16037 16099
rect 16037 16065 16071 16099
rect 16071 16065 16080 16099
rect 16028 16056 16080 16065
rect 14464 15988 14516 16040
rect 15108 15988 15160 16040
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 5172 15852 5224 15904
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 6000 15852 6052 15904
rect 7288 15852 7340 15904
rect 11612 15852 11664 15904
rect 12164 15852 12216 15904
rect 12532 15852 12584 15904
rect 16120 15920 16172 15972
rect 16580 15920 16632 15972
rect 13636 15852 13688 15904
rect 16856 15852 16908 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1400 15648 1452 15700
rect 3240 15648 3292 15700
rect 5632 15648 5684 15700
rect 7012 15648 7064 15700
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 10140 15691 10192 15700
rect 10140 15657 10149 15691
rect 10149 15657 10183 15691
rect 10183 15657 10192 15691
rect 10140 15648 10192 15657
rect 12164 15691 12216 15700
rect 12164 15657 12173 15691
rect 12173 15657 12207 15691
rect 12207 15657 12216 15691
rect 12164 15648 12216 15657
rect 13544 15648 13596 15700
rect 14280 15648 14332 15700
rect 1492 15580 1544 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3516 15444 3568 15496
rect 6000 15580 6052 15632
rect 7196 15623 7248 15632
rect 7196 15589 7205 15623
rect 7205 15589 7239 15623
rect 7239 15589 7248 15623
rect 7196 15580 7248 15589
rect 6276 15512 6328 15564
rect 6368 15512 6420 15564
rect 9956 15512 10008 15564
rect 13268 15580 13320 15632
rect 16396 15648 16448 15700
rect 8300 15444 8352 15496
rect 9864 15444 9916 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 5816 15308 5868 15360
rect 7472 15308 7524 15360
rect 12348 15512 12400 15564
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 13820 15512 13872 15564
rect 14464 15512 14516 15564
rect 15016 15512 15068 15564
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 12440 15444 12492 15496
rect 13912 15444 13964 15496
rect 14556 15444 14608 15496
rect 15844 15444 15896 15496
rect 16580 15444 16632 15496
rect 17408 15444 17460 15496
rect 16028 15376 16080 15428
rect 11152 15308 11204 15360
rect 13084 15308 13136 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 5080 15104 5132 15156
rect 5724 15104 5776 15156
rect 6000 15036 6052 15088
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 6276 15011 6328 15020
rect 2780 14968 2832 14977
rect 6276 14977 6285 15011
rect 6285 14977 6319 15011
rect 6319 14977 6328 15011
rect 6276 14968 6328 14977
rect 8852 15104 8904 15156
rect 9864 15147 9916 15156
rect 9864 15113 9873 15147
rect 9873 15113 9907 15147
rect 9907 15113 9916 15147
rect 9864 15104 9916 15113
rect 13176 15104 13228 15156
rect 15660 15147 15712 15156
rect 15660 15113 15669 15147
rect 15669 15113 15703 15147
rect 15703 15113 15712 15147
rect 15660 15104 15712 15113
rect 17408 15147 17460 15156
rect 17408 15113 17417 15147
rect 17417 15113 17451 15147
rect 17451 15113 17460 15147
rect 17408 15104 17460 15113
rect 11612 15011 11664 15020
rect 11612 14977 11621 15011
rect 11621 14977 11655 15011
rect 11655 14977 11664 15011
rect 11612 14968 11664 14977
rect 16028 15011 16080 15020
rect 3976 14900 4028 14952
rect 6552 14900 6604 14952
rect 8300 14900 8352 14952
rect 9680 14900 9732 14952
rect 10232 14900 10284 14952
rect 11060 14900 11112 14952
rect 12348 14900 12400 14952
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 14556 14943 14608 14952
rect 14556 14909 14579 14943
rect 14579 14909 14608 14943
rect 2964 14764 3016 14816
rect 5816 14832 5868 14884
rect 6368 14832 6420 14884
rect 14556 14900 14608 14909
rect 18052 14900 18104 14952
rect 3516 14764 3568 14816
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 7472 14764 7524 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 16948 14832 17000 14884
rect 18512 14832 18564 14884
rect 13544 14764 13596 14773
rect 15568 14764 15620 14816
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 19524 14764 19576 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 4804 14560 4856 14612
rect 7104 14560 7156 14612
rect 14556 14603 14608 14612
rect 14556 14569 14565 14603
rect 14565 14569 14599 14603
rect 14599 14569 14608 14603
rect 14556 14560 14608 14569
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 1400 14492 1452 14544
rect 7012 14492 7064 14544
rect 11612 14492 11664 14544
rect 17960 14492 18012 14544
rect 18696 14492 18748 14544
rect 19524 14492 19576 14544
rect 1952 14424 2004 14476
rect 2504 14424 2556 14476
rect 6000 14467 6052 14476
rect 6000 14433 6009 14467
rect 6009 14433 6043 14467
rect 6043 14433 6052 14467
rect 6000 14424 6052 14433
rect 7472 14424 7524 14476
rect 7748 14424 7800 14476
rect 8300 14424 8352 14476
rect 10232 14424 10284 14476
rect 10416 14467 10468 14476
rect 10416 14433 10425 14467
rect 10425 14433 10459 14467
rect 10459 14433 10468 14467
rect 10416 14424 10468 14433
rect 13084 14424 13136 14476
rect 13268 14424 13320 14476
rect 14372 14424 14424 14476
rect 15108 14424 15160 14476
rect 18052 14467 18104 14476
rect 18052 14433 18061 14467
rect 18061 14433 18095 14467
rect 18095 14433 18104 14467
rect 18052 14424 18104 14433
rect 3332 14399 3384 14408
rect 3332 14365 3341 14399
rect 3341 14365 3375 14399
rect 3375 14365 3384 14399
rect 3332 14356 3384 14365
rect 5540 14399 5592 14408
rect 4160 14288 4212 14340
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 17040 14356 17092 14408
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 17132 14288 17184 14340
rect 2964 14220 3016 14272
rect 6368 14220 6420 14272
rect 11612 14220 11664 14272
rect 18788 14220 18840 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2504 14059 2556 14068
rect 2504 14025 2513 14059
rect 2513 14025 2547 14059
rect 2547 14025 2556 14059
rect 2504 14016 2556 14025
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 5080 14016 5132 14068
rect 9680 14016 9732 14068
rect 11796 14016 11848 14068
rect 13544 14016 13596 14068
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 10416 13923 10468 13932
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 11060 13880 11112 13932
rect 11612 13880 11664 13932
rect 11796 13880 11848 13932
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13360 13880 13412 13932
rect 16028 14016 16080 14068
rect 16304 14016 16356 14068
rect 16948 14016 17000 14068
rect 17500 14016 17552 14068
rect 3332 13812 3384 13864
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 4160 13812 4212 13864
rect 5540 13812 5592 13864
rect 7012 13812 7064 13864
rect 7656 13812 7708 13864
rect 8852 13812 8904 13864
rect 13912 13812 13964 13864
rect 15108 13855 15160 13864
rect 15108 13821 15117 13855
rect 15117 13821 15151 13855
rect 15151 13821 15160 13855
rect 15108 13812 15160 13821
rect 15936 13855 15988 13864
rect 15936 13821 15970 13855
rect 15970 13821 15988 13855
rect 15936 13812 15988 13821
rect 17224 13812 17276 13864
rect 8668 13744 8720 13796
rect 11152 13787 11204 13796
rect 7104 13676 7156 13728
rect 11152 13753 11161 13787
rect 11161 13753 11195 13787
rect 11195 13753 11204 13787
rect 11152 13744 11204 13753
rect 11244 13744 11296 13796
rect 12532 13744 12584 13796
rect 15016 13787 15068 13796
rect 11060 13676 11112 13728
rect 13820 13676 13872 13728
rect 15016 13753 15025 13787
rect 15025 13753 15059 13787
rect 15059 13753 15068 13787
rect 15016 13744 15068 13753
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 18512 13812 18564 13864
rect 17960 13744 18012 13796
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1860 13472 1912 13524
rect 6184 13472 6236 13524
rect 6276 13472 6328 13524
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 4068 13404 4120 13456
rect 11244 13472 11296 13524
rect 13268 13472 13320 13524
rect 13636 13472 13688 13524
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 15752 13472 15804 13524
rect 16672 13515 16724 13524
rect 16672 13481 16681 13515
rect 16681 13481 16715 13515
rect 16715 13481 16724 13515
rect 16672 13472 16724 13481
rect 17132 13515 17184 13524
rect 17132 13481 17141 13515
rect 17141 13481 17175 13515
rect 17175 13481 17184 13515
rect 17132 13472 17184 13481
rect 10784 13447 10836 13456
rect 10784 13413 10793 13447
rect 10793 13413 10827 13447
rect 10827 13413 10836 13447
rect 10784 13404 10836 13413
rect 17040 13447 17092 13456
rect 6000 13336 6052 13388
rect 7748 13336 7800 13388
rect 4712 13268 4764 13320
rect 7012 13200 7064 13252
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 13360 13336 13412 13388
rect 17040 13413 17049 13447
rect 17049 13413 17083 13447
rect 17083 13413 17092 13447
rect 17040 13404 17092 13413
rect 16856 13336 16908 13388
rect 16948 13336 17000 13388
rect 12716 13268 12768 13320
rect 13820 13268 13872 13320
rect 15752 13268 15804 13320
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 16764 13268 16816 13320
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 2596 12928 2648 12980
rect 6000 12928 6052 12980
rect 2872 12860 2924 12912
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 6184 12928 6236 12980
rect 8668 12928 8720 12980
rect 10416 12928 10468 12980
rect 13452 12928 13504 12980
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 11060 12860 11112 12912
rect 13636 12835 13688 12844
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 2964 12724 3016 12776
rect 7656 12724 7708 12776
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 11612 12724 11664 12776
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 12532 12724 12584 12776
rect 15384 12724 15436 12776
rect 15476 12724 15528 12776
rect 17960 12724 18012 12776
rect 18788 12724 18840 12776
rect 5448 12656 5500 12708
rect 9128 12656 9180 12708
rect 16764 12656 16816 12708
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 11980 12631 12032 12640
rect 7288 12588 7340 12597
rect 11980 12597 11989 12631
rect 11989 12597 12023 12631
rect 12023 12597 12032 12631
rect 11980 12588 12032 12597
rect 13544 12631 13596 12640
rect 13544 12597 13553 12631
rect 13553 12597 13587 12631
rect 13587 12597 13596 12631
rect 19432 12631 19484 12640
rect 13544 12588 13596 12597
rect 19432 12597 19441 12631
rect 19441 12597 19475 12631
rect 19475 12597 19484 12631
rect 19432 12588 19484 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 1768 12316 1820 12368
rect 2964 12359 3016 12368
rect 2964 12325 2973 12359
rect 2973 12325 3007 12359
rect 3007 12325 3016 12359
rect 2964 12316 3016 12325
rect 1860 12248 1912 12300
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 8484 12384 8536 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 4068 12316 4120 12368
rect 4160 12248 4212 12300
rect 4712 12316 4764 12368
rect 5540 12316 5592 12368
rect 6552 12316 6604 12368
rect 11980 12384 12032 12436
rect 13544 12384 13596 12436
rect 14004 12384 14056 12436
rect 16764 12427 16816 12436
rect 10416 12316 10468 12368
rect 12532 12359 12584 12368
rect 12532 12325 12541 12359
rect 12541 12325 12575 12359
rect 12575 12325 12584 12359
rect 12532 12316 12584 12325
rect 15660 12359 15712 12368
rect 6828 12248 6880 12300
rect 8484 12248 8536 12300
rect 2320 12112 2372 12164
rect 5540 12180 5592 12232
rect 7104 12180 7156 12232
rect 8208 12223 8260 12232
rect 4252 12044 4304 12096
rect 4712 12044 4764 12096
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 7564 12112 7616 12164
rect 10048 12248 10100 12300
rect 11152 12248 11204 12300
rect 15660 12325 15683 12359
rect 15683 12325 15712 12359
rect 15660 12316 15712 12325
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 16856 12384 16908 12436
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 17776 12316 17828 12368
rect 13544 12248 13596 12300
rect 14464 12291 14516 12300
rect 14464 12257 14473 12291
rect 14473 12257 14507 12291
rect 14507 12257 14516 12291
rect 14464 12248 14516 12257
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10416 12180 10468 12232
rect 13636 12223 13688 12232
rect 12808 12112 12860 12164
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 13820 12180 13872 12232
rect 16672 12248 16724 12300
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 19432 12248 19484 12300
rect 19248 12223 19300 12232
rect 19248 12189 19257 12223
rect 19257 12189 19291 12223
rect 19291 12189 19300 12223
rect 19248 12180 19300 12189
rect 10508 12044 10560 12096
rect 11888 12087 11940 12096
rect 11888 12053 11897 12087
rect 11897 12053 11931 12087
rect 11931 12053 11940 12087
rect 11888 12044 11940 12053
rect 13084 12044 13136 12096
rect 17316 12044 17368 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 2688 11840 2740 11892
rect 7288 11840 7340 11892
rect 9128 11840 9180 11892
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 14096 11840 14148 11892
rect 15660 11840 15712 11892
rect 16120 11883 16172 11892
rect 16120 11849 16129 11883
rect 16129 11849 16163 11883
rect 16163 11849 16172 11883
rect 16120 11840 16172 11849
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 4160 11772 4212 11824
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2320 11636 2372 11688
rect 4068 11636 4120 11688
rect 5448 11704 5500 11756
rect 6644 11704 6696 11756
rect 6736 11636 6788 11688
rect 7104 11704 7156 11756
rect 7564 11636 7616 11688
rect 7656 11636 7708 11688
rect 10508 11704 10560 11756
rect 15476 11772 15528 11824
rect 16212 11772 16264 11824
rect 17960 11772 18012 11824
rect 11612 11704 11664 11756
rect 11888 11704 11940 11756
rect 13636 11704 13688 11756
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 4620 11568 4672 11620
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 5724 11500 5776 11552
rect 6644 11500 6696 11552
rect 6920 11568 6972 11620
rect 8208 11611 8260 11620
rect 8208 11577 8242 11611
rect 8242 11577 8260 11611
rect 8208 11568 8260 11577
rect 9036 11568 9088 11620
rect 14004 11568 14056 11620
rect 14556 11636 14608 11688
rect 15568 11636 15620 11688
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 19432 11636 19484 11688
rect 19984 11611 20036 11620
rect 7104 11500 7156 11552
rect 8852 11500 8904 11552
rect 15292 11500 15344 11552
rect 15384 11500 15436 11552
rect 18144 11500 18196 11552
rect 19156 11500 19208 11552
rect 19984 11577 20018 11611
rect 20018 11577 20036 11611
rect 19984 11568 20036 11577
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2780 11296 2832 11348
rect 4712 11296 4764 11348
rect 9036 11339 9088 11348
rect 9036 11305 9045 11339
rect 9045 11305 9079 11339
rect 9079 11305 9088 11339
rect 9036 11296 9088 11305
rect 13268 11296 13320 11348
rect 14556 11296 14608 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 12348 11271 12400 11280
rect 4160 11160 4212 11212
rect 6920 11160 6972 11212
rect 7196 11160 7248 11212
rect 7932 11203 7984 11212
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 3700 11092 3752 11144
rect 4712 11135 4764 11144
rect 4252 11024 4304 11076
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 7932 11169 7966 11203
rect 7966 11169 7984 11203
rect 7932 11160 7984 11169
rect 8208 11160 8260 11212
rect 10508 11203 10560 11212
rect 10508 11169 10542 11203
rect 10542 11169 10560 11203
rect 10508 11160 10560 11169
rect 12348 11237 12357 11271
rect 12357 11237 12391 11271
rect 12391 11237 12400 11271
rect 12348 11228 12400 11237
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 4804 11024 4856 11076
rect 2872 10999 2924 11008
rect 2872 10965 2881 10999
rect 2881 10965 2915 10999
rect 2915 10965 2924 10999
rect 2872 10956 2924 10965
rect 5080 10956 5132 11008
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 6828 11024 6880 11076
rect 7104 10956 7156 11008
rect 11612 11067 11664 11076
rect 11612 11033 11621 11067
rect 11621 11033 11655 11067
rect 11655 11033 11664 11067
rect 11612 11024 11664 11033
rect 12072 11024 12124 11076
rect 12716 11024 12768 11076
rect 14556 11092 14608 11144
rect 17592 11067 17644 11076
rect 17592 11033 17601 11067
rect 17601 11033 17635 11067
rect 17635 11033 17644 11067
rect 19432 11092 19484 11144
rect 17592 11024 17644 11033
rect 12164 10956 12216 11008
rect 15384 10956 15436 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1676 10752 1728 10804
rect 3332 10752 3384 10804
rect 8484 10795 8536 10804
rect 3792 10684 3844 10736
rect 7932 10684 7984 10736
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 12072 10795 12124 10804
rect 12072 10761 12081 10795
rect 12081 10761 12115 10795
rect 12115 10761 12124 10795
rect 12072 10752 12124 10761
rect 12348 10752 12400 10804
rect 2688 10659 2740 10668
rect 2688 10625 2697 10659
rect 2697 10625 2731 10659
rect 2731 10625 2740 10659
rect 2688 10616 2740 10625
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 5540 10616 5592 10668
rect 10048 10616 10100 10668
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 14556 10752 14608 10804
rect 16488 10795 16540 10804
rect 16488 10761 16497 10795
rect 16497 10761 16531 10795
rect 16531 10761 16540 10795
rect 16488 10752 16540 10761
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 2872 10548 2924 10600
rect 4988 10548 5040 10600
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 4068 10480 4120 10532
rect 7104 10523 7156 10532
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 4436 10455 4488 10464
rect 3516 10412 3568 10421
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 7104 10489 7138 10523
rect 7138 10489 7156 10523
rect 7104 10480 7156 10489
rect 12164 10548 12216 10600
rect 12716 10548 12768 10600
rect 13084 10548 13136 10600
rect 15660 10548 15712 10600
rect 11612 10480 11664 10532
rect 11980 10412 12032 10464
rect 13360 10480 13412 10532
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17960 10616 18012 10668
rect 19156 10548 19208 10600
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 3976 10208 4028 10260
rect 13084 10208 13136 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13728 10208 13780 10260
rect 3700 10140 3752 10192
rect 4436 10140 4488 10192
rect 4988 10140 5040 10192
rect 2320 10072 2372 10124
rect 4712 10072 4764 10124
rect 6000 10115 6052 10124
rect 6000 10081 6034 10115
rect 6034 10081 6052 10115
rect 6000 10072 6052 10081
rect 6920 10140 6972 10192
rect 9680 10140 9732 10192
rect 12072 10140 12124 10192
rect 10324 10072 10376 10124
rect 10692 10072 10744 10124
rect 12716 10072 12768 10124
rect 14004 10115 14056 10124
rect 14004 10081 14013 10115
rect 14013 10081 14047 10115
rect 14047 10081 14056 10115
rect 14004 10072 14056 10081
rect 7656 10004 7708 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 13268 10004 13320 10056
rect 16212 10115 16264 10124
rect 16212 10081 16221 10115
rect 16221 10081 16255 10115
rect 16255 10081 16264 10115
rect 16212 10072 16264 10081
rect 17040 10072 17092 10124
rect 5080 9936 5132 9988
rect 2688 9868 2740 9920
rect 3700 9868 3752 9920
rect 7104 9911 7156 9920
rect 7104 9877 7113 9911
rect 7113 9877 7147 9911
rect 7147 9877 7156 9911
rect 7104 9868 7156 9877
rect 7656 9911 7708 9920
rect 7656 9877 7665 9911
rect 7665 9877 7699 9911
rect 7699 9877 7708 9911
rect 7656 9868 7708 9877
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 3516 9664 3568 9716
rect 6000 9664 6052 9716
rect 4160 9639 4212 9648
rect 4160 9605 4169 9639
rect 4169 9605 4203 9639
rect 4203 9605 4212 9639
rect 4160 9596 4212 9605
rect 4252 9596 4304 9648
rect 5080 9528 5132 9580
rect 7104 9528 7156 9580
rect 8576 9664 8628 9716
rect 17040 9707 17092 9716
rect 17040 9673 17049 9707
rect 17049 9673 17083 9707
rect 17083 9673 17092 9707
rect 17040 9664 17092 9673
rect 10324 9639 10376 9648
rect 10324 9605 10333 9639
rect 10333 9605 10367 9639
rect 10367 9605 10376 9639
rect 10324 9596 10376 9605
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 14004 9528 14056 9580
rect 16856 9528 16908 9580
rect 4712 9460 4764 9512
rect 7932 9460 7984 9512
rect 4252 9392 4304 9444
rect 6000 9392 6052 9444
rect 4160 9324 4212 9376
rect 5816 9324 5868 9376
rect 6184 9324 6236 9376
rect 7012 9392 7064 9444
rect 7656 9392 7708 9444
rect 16212 9460 16264 9512
rect 12256 9392 12308 9444
rect 12348 9392 12400 9444
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 7472 9324 7524 9376
rect 16120 9392 16172 9444
rect 18512 9324 18564 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2044 9120 2096 9172
rect 4896 9120 4948 9172
rect 7196 9120 7248 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 4068 9052 4120 9104
rect 12348 9052 12400 9104
rect 1676 8984 1728 9036
rect 3608 8984 3660 9036
rect 5724 8984 5776 9036
rect 7472 8984 7524 9036
rect 7840 8984 7892 9036
rect 8760 8984 8812 9036
rect 4160 8916 4212 8968
rect 4896 8916 4948 8968
rect 5080 8916 5132 8968
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 7196 8916 7248 8968
rect 7656 8916 7708 8968
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 5908 8780 5960 8832
rect 10876 8916 10928 8968
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 7840 8576 7892 8628
rect 3516 8508 3568 8560
rect 5356 8508 5408 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 9128 8440 9180 8492
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2688 8372 2740 8424
rect 4804 8372 4856 8424
rect 8760 8372 8812 8424
rect 8852 8372 8904 8424
rect 11704 8372 11756 8424
rect 3516 8279 3568 8288
rect 3516 8245 3525 8279
rect 3525 8245 3559 8279
rect 3559 8245 3568 8279
rect 3516 8236 3568 8245
rect 4160 8279 4212 8288
rect 4160 8245 4169 8279
rect 4169 8245 4203 8279
rect 4203 8245 4212 8279
rect 4160 8236 4212 8245
rect 5540 8347 5592 8356
rect 4804 8236 4856 8288
rect 5540 8313 5549 8347
rect 5549 8313 5583 8347
rect 5583 8313 5592 8347
rect 5540 8304 5592 8313
rect 5724 8304 5776 8356
rect 8208 8304 8260 8356
rect 8852 8279 8904 8288
rect 8852 8245 8861 8279
rect 8861 8245 8895 8279
rect 8895 8245 8904 8279
rect 8852 8236 8904 8245
rect 9404 8236 9456 8288
rect 17592 8236 17644 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 1492 8032 1544 8084
rect 4160 8032 4212 8084
rect 4896 8032 4948 8084
rect 8760 8032 8812 8084
rect 8852 8032 8904 8084
rect 19708 8032 19760 8084
rect 4068 7964 4120 8016
rect 9404 7964 9456 8016
rect 4160 7896 4212 7948
rect 6000 7896 6052 7948
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 8852 7939 8904 7948
rect 4252 7692 4304 7744
rect 6736 7692 6788 7744
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 8944 7896 8996 7948
rect 8208 7828 8260 7880
rect 9128 7760 9180 7812
rect 7196 7692 7248 7744
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 4068 7488 4120 7540
rect 6000 7531 6052 7540
rect 6000 7497 6009 7531
rect 6009 7497 6043 7531
rect 6043 7497 6052 7531
rect 6000 7488 6052 7497
rect 6736 7488 6788 7540
rect 19340 7488 19392 7540
rect 8944 7420 8996 7472
rect 8208 7352 8260 7404
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 2136 7284 2188 7336
rect 5172 7284 5224 7336
rect 6092 7284 6144 7336
rect 8668 7284 8720 7336
rect 8760 7284 8812 7336
rect 18972 7327 19024 7336
rect 18972 7293 18981 7327
rect 18981 7293 19015 7327
rect 19015 7293 19024 7327
rect 18972 7284 19024 7293
rect 3516 7216 3568 7268
rect 4712 7216 4764 7268
rect 5540 7216 5592 7268
rect 7564 7148 7616 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 7564 6987 7616 6996
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 8852 6944 8904 6996
rect 4068 6876 4120 6928
rect 18972 6876 19024 6928
rect 8484 6808 8536 6860
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 19248 6808 19300 6860
rect 3884 6740 3936 6792
rect 4712 6783 4764 6792
rect 4160 6672 4212 6724
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 9128 6740 9180 6792
rect 9220 6740 9272 6792
rect 9680 6740 9732 6792
rect 7288 6672 7340 6724
rect 19616 6715 19668 6724
rect 19616 6681 19625 6715
rect 19625 6681 19659 6715
rect 19659 6681 19668 6715
rect 19616 6672 19668 6681
rect 4804 6604 4856 6656
rect 9680 6604 9732 6656
rect 19248 6604 19300 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 5816 6400 5868 6452
rect 6184 6400 6236 6452
rect 8760 6400 8812 6452
rect 20996 6400 21048 6452
rect 3976 6196 4028 6248
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 20812 5856 20864 5908
rect 4068 5720 4120 5772
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 20904 5312 20956 5364
rect 4068 5108 4120 5160
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3976 4088 4028 4140
rect 4896 4088 4948 4140
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2780 2524 2832 2576
rect 5632 2524 5684 2576
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 3700 1980 3752 2032
rect 5540 1980 5592 2032
rect 3700 1708 3752 1760
rect 5724 1708 5776 1760
rect 4068 1028 4120 1080
rect 5816 1028 5868 1080
rect 3240 416 3292 468
rect 4988 416 5040 468
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 1030 22320 1086 22800
rect 1398 22536 1454 22545
rect 1398 22471 1454 22480
rect 216 19242 244 22320
rect 204 19236 256 19242
rect 204 19178 256 19184
rect 584 18358 612 22320
rect 1044 18902 1072 22320
rect 1032 18896 1084 18902
rect 1032 18838 1084 18844
rect 572 18352 624 18358
rect 572 18294 624 18300
rect 1412 15706 1440 22471
rect 1490 22320 1546 22800
rect 1950 22320 2006 22800
rect 2410 22320 2466 22800
rect 2870 22320 2926 22800
rect 3330 22320 3386 22800
rect 3790 22320 3846 22800
rect 4250 22320 4306 22800
rect 4710 22320 4766 22800
rect 5170 22320 5226 22800
rect 5630 22320 5686 22800
rect 6090 22320 6146 22800
rect 6550 22320 6606 22800
rect 7010 22320 7066 22800
rect 7470 22320 7526 22800
rect 7930 22320 7986 22800
rect 8390 22320 8446 22800
rect 8850 22320 8906 22800
rect 9310 22320 9366 22800
rect 9770 22320 9826 22800
rect 10230 22320 10286 22800
rect 10690 22320 10746 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12438 22320 12494 22800
rect 12898 22320 12954 22800
rect 13358 22320 13414 22800
rect 13818 22320 13874 22800
rect 14278 22320 14334 22800
rect 14738 22320 14794 22800
rect 15198 22320 15254 22800
rect 15658 22320 15714 22800
rect 16118 22320 16174 22800
rect 16578 22320 16634 22800
rect 17038 22320 17094 22800
rect 17498 22320 17554 22800
rect 17958 22320 18014 22800
rect 18418 22320 18474 22800
rect 18878 22320 18934 22800
rect 19338 22320 19394 22800
rect 19798 22320 19854 22800
rect 20258 22320 20314 22800
rect 20718 22320 20774 22800
rect 21178 22320 21234 22800
rect 21638 22320 21694 22800
rect 22098 22320 22154 22800
rect 22558 22320 22614 22800
rect 1504 19145 1532 22320
rect 1582 20224 1638 20233
rect 1582 20159 1638 20168
rect 1490 19136 1546 19145
rect 1490 19071 1546 19080
rect 1596 18970 1624 20159
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1780 19378 1808 19858
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1688 18154 1716 19246
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1780 17921 1808 18022
rect 1766 17912 1822 17921
rect 1766 17847 1822 17856
rect 1676 16992 1728 16998
rect 1674 16960 1676 16969
rect 1728 16960 1730 16969
rect 1674 16895 1730 16904
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1504 15638 1532 16594
rect 1674 16552 1730 16561
rect 1674 16487 1676 16496
rect 1728 16487 1730 16496
rect 1676 16458 1728 16464
rect 1766 16008 1822 16017
rect 1766 15943 1822 15952
rect 1492 15632 1544 15638
rect 1492 15574 1544 15580
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 14550 1440 15506
rect 1780 14618 1808 15943
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1400 14544 1452 14550
rect 1400 14486 1452 14492
rect 1490 14104 1546 14113
rect 1490 14039 1546 14048
rect 1504 8090 1532 14039
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1596 12442 1624 13631
rect 1872 13530 1900 19751
rect 1964 18952 1992 22320
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2240 19310 2268 19654
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 1964 18924 2268 18952
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 18426 1992 18770
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1950 18320 2006 18329
rect 1950 18255 2006 18264
rect 1964 17882 1992 18255
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2056 16114 2084 18702
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2148 18222 2176 18566
rect 2240 18329 2268 18924
rect 2332 18902 2360 19858
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2226 18320 2282 18329
rect 2226 18255 2282 18264
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 2424 18057 2452 22320
rect 2884 22250 2912 22320
rect 2884 22222 3280 22250
rect 3054 22128 3110 22137
rect 3054 22063 3110 22072
rect 2962 21584 3018 21593
rect 2962 21519 3018 21528
rect 2870 21176 2926 21185
rect 2870 21111 2926 21120
rect 2778 20632 2834 20641
rect 2778 20567 2834 20576
rect 2792 19786 2820 20567
rect 2884 20058 2912 21111
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2872 19304 2924 19310
rect 2594 19272 2650 19281
rect 2872 19246 2924 19252
rect 2594 19207 2650 19216
rect 2410 18048 2466 18057
rect 2410 17983 2466 17992
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2424 16726 2452 17682
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2516 17377 2544 17478
rect 2502 17368 2558 17377
rect 2502 17303 2558 17312
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2042 14648 2098 14657
rect 2042 14583 2098 14592
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1964 13938 1992 14418
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1780 12374 1808 12718
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1872 11762 1900 12242
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1688 10810 1716 11630
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 2056 9178 2084 14583
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2516 14074 2544 14418
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2608 12986 2636 19207
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2792 18193 2820 18294
rect 2884 18222 2912 19246
rect 2976 19174 3004 21519
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2962 18864 3018 18873
rect 2962 18799 3018 18808
rect 2872 18216 2924 18222
rect 2778 18184 2834 18193
rect 2872 18158 2924 18164
rect 2778 18119 2834 18128
rect 2884 17610 2912 18158
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2884 17202 2912 17546
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16522 2912 17138
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2884 15994 2912 16458
rect 2792 15978 2912 15994
rect 2780 15972 2912 15978
rect 2832 15966 2912 15972
rect 2780 15914 2832 15920
rect 2792 15026 2820 15914
rect 2870 15600 2926 15609
rect 2870 15535 2926 15544
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2778 14784 2834 14793
rect 2778 14719 2834 14728
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2332 11694 2360 12106
rect 2700 11898 2728 12242
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2332 10130 2360 11630
rect 2792 11354 2820 14719
rect 2884 12918 2912 15535
rect 2976 14822 3004 18799
rect 3068 17882 3096 22063
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3160 18902 3188 19178
rect 3252 19009 3280 22222
rect 3344 19530 3372 22320
rect 3344 19514 3464 19530
rect 3344 19508 3476 19514
rect 3344 19502 3424 19508
rect 3424 19450 3476 19456
rect 3238 19000 3294 19009
rect 3238 18935 3294 18944
rect 3148 18896 3200 18902
rect 3148 18838 3200 18844
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3344 17882 3372 18770
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3528 18086 3556 18702
rect 3804 18698 3832 22320
rect 4264 19394 4292 22320
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4264 19366 4384 19394
rect 4356 19310 4384 19366
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 18766 4292 19110
rect 4436 18964 4488 18970
rect 4488 18924 4568 18952
rect 4436 18906 4488 18912
rect 4252 18760 4304 18766
rect 4540 18737 4568 18924
rect 4252 18702 4304 18708
rect 4526 18728 4582 18737
rect 3792 18692 3844 18698
rect 3792 18634 3844 18640
rect 4264 18154 4292 18702
rect 4526 18663 4582 18672
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 3516 18080 3568 18086
rect 4436 18080 4488 18086
rect 3516 18022 3568 18028
rect 4434 18048 4436 18057
rect 4488 18048 4490 18057
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3528 17066 3556 18022
rect 4434 17983 4490 17992
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3804 17134 3832 17478
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3884 17060 3936 17066
rect 3884 17002 3936 17008
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3252 15706 3280 16594
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3528 14822 3556 15438
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2976 13938 3004 14214
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 3344 13870 3372 14350
rect 3528 13870 3556 14758
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2976 12374 3004 12718
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 3238 12200 3294 12209
rect 3238 12135 3294 12144
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8498 1716 8978
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 2136 8424 2188 8430
rect 2332 8412 2360 10066
rect 2700 9926 2728 10610
rect 2884 10606 2912 10950
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 8430 2728 9862
rect 2188 8384 2360 8412
rect 2688 8424 2740 8430
rect 2136 8366 2188 8372
rect 2688 8366 2740 8372
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 2148 7342 2176 8366
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 3252 4321 3280 12135
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3344 10810 3372 11086
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3712 10674 3740 11086
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3436 10266 3464 10406
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3422 10160 3478 10169
rect 3422 10095 3478 10104
rect 3436 9489 3464 10095
rect 3528 9722 3556 10406
rect 3712 10198 3740 10610
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3712 9926 3740 10134
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3422 9480 3478 9489
rect 3422 9415 3478 9424
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3528 8294 3556 8502
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 7274 3556 8230
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3238 4312 3294 4321
rect 3238 4247 3294 4256
rect 2780 2576 2832 2582
rect 2778 2544 2780 2553
rect 2832 2544 2834 2553
rect 2778 2479 2834 2488
rect 3620 649 3648 8978
rect 3804 7585 3832 10678
rect 3896 9081 3924 17002
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3988 15910 4016 16526
rect 4172 16046 4200 16934
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4264 16250 4292 16594
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4724 16114 4752 22320
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3988 14958 4016 15846
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14346 4200 14758
rect 4816 14618 4844 19246
rect 4908 19174 4936 19790
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 5092 18766 5120 19246
rect 5184 18970 5212 22320
rect 5644 20058 5672 22320
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5920 19242 5948 19790
rect 5908 19236 5960 19242
rect 5908 19178 5960 19184
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4172 13870 4200 14282
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4080 12753 4108 13398
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4724 12850 4752 13262
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4724 12374 4752 12786
rect 4068 12368 4120 12374
rect 4066 12336 4068 12345
rect 4712 12368 4764 12374
rect 4120 12336 4122 12345
rect 4250 12336 4306 12345
rect 4066 12271 4122 12280
rect 4160 12300 4212 12306
rect 4250 12271 4306 12280
rect 4710 12336 4712 12345
rect 4764 12336 4766 12345
rect 4710 12271 4766 12280
rect 4160 12242 4212 12248
rect 4172 11830 4200 12242
rect 4264 12102 4292 12271
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4724 11880 4752 12038
rect 4632 11852 4752 11880
rect 4160 11824 4212 11830
rect 4066 11792 4122 11801
rect 4160 11766 4212 11772
rect 4066 11727 4122 11736
rect 4080 11694 4108 11727
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4632 11626 4660 11852
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4632 11234 4660 11562
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4724 11354 4752 11494
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4160 11212 4212 11218
rect 4632 11206 4752 11234
rect 4160 11154 4212 11160
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 3988 10266 4016 10775
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4080 10441 4108 10474
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4172 9654 4200 11154
rect 4724 11150 4752 11206
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4264 9654 4292 11018
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 10198 4476 10406
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4724 10130 4752 10610
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4816 10010 4844 11018
rect 4724 9982 4844 10010
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4724 9518 4752 9982
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4068 9104 4120 9110
rect 3882 9072 3938 9081
rect 4068 9046 4120 9052
rect 3882 9007 3938 9016
rect 4080 8537 4108 9046
rect 4172 8974 4200 9318
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4066 8120 4122 8129
rect 4172 8090 4200 8230
rect 4066 8055 4122 8064
rect 4160 8084 4212 8090
rect 4080 8022 4108 8055
rect 4160 8026 4212 8032
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3790 7576 3846 7585
rect 3790 7511 3846 7520
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4080 7177 4108 7482
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 3884 6792 3936 6798
rect 4080 6769 4108 6870
rect 3884 6734 3936 6740
rect 4066 6760 4122 6769
rect 3896 3505 3924 6734
rect 4172 6730 4200 7890
rect 4264 7750 4292 9386
rect 4908 9178 4936 16118
rect 5000 10606 5028 18634
rect 5920 18290 5948 18838
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5276 17270 5304 17614
rect 5736 17338 5764 18226
rect 5920 17882 5948 18226
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5264 17264 5316 17270
rect 5264 17206 5316 17212
rect 6012 17082 6040 19858
rect 6104 17202 6132 22320
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6196 17202 6224 17682
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6012 17054 6132 17082
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5828 16114 5856 16594
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 5092 14074 5120 15098
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5092 10418 5120 10950
rect 5000 10390 5120 10418
rect 5000 10198 5028 10390
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4066 6695 4122 6704
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5817 4016 6190
rect 3974 5808 4030 5817
rect 3974 5743 4030 5752
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5273 4108 5714
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4865 4108 5102
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3882 3496 3938 3505
rect 3882 3431 3938 3440
rect 3988 2961 4016 4082
rect 4264 3913 4292 7686
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4724 7274 4752 8434
rect 4816 8430 4844 8774
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4724 6798 4752 7210
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4816 6662 4844 8230
rect 4908 8090 4936 8910
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4908 4146 4936 8026
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4250 3904 4306 3913
rect 4250 3839 4306 3848
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 3974 2952 4030 2961
rect 3974 2887 4030 2896
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 3700 2032 3752 2038
rect 3698 2000 3700 2009
rect 3752 2000 3754 2009
rect 3698 1935 3754 1944
rect 3700 1760 3752 1766
rect 3700 1702 3752 1708
rect 3712 1601 3740 1702
rect 3698 1592 3754 1601
rect 3698 1527 3754 1536
rect 4068 1080 4120 1086
rect 4066 1048 4068 1057
rect 4120 1048 4122 1057
rect 4066 983 4122 992
rect 3606 640 3662 649
rect 3606 575 3662 584
rect 5000 474 5028 10134
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5092 9586 5120 9930
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5184 9466 5212 15846
rect 5644 15706 5672 15846
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5736 15162 5764 15846
rect 5828 15366 5856 16050
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 13870 5580 14350
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5460 12102 5488 12650
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5552 12238 5580 12310
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11762 5488 12038
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5552 11014 5580 12174
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10674 5580 10950
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5092 9438 5212 9466
rect 5092 8974 5120 9438
rect 5736 9042 5764 11494
rect 5828 9382 5856 14826
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8566 5396 8910
rect 5920 8838 5948 16934
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6012 15638 6040 15846
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 6012 15094 6040 15574
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 6012 14482 6040 15030
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6012 12986 6040 13330
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9722 6040 10066
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6012 9330 6040 9386
rect 6104 9330 6132 17054
rect 6196 16794 6224 17138
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6288 15026 6316 15506
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6288 13530 6316 14962
rect 6380 14890 6408 15506
rect 6564 14958 6592 22320
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6840 18970 6868 19178
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 7024 18034 7052 22320
rect 7484 19394 7512 22320
rect 7944 20346 7972 22320
rect 7208 19366 7512 19394
rect 7668 20318 7972 20346
rect 7102 19000 7158 19009
rect 7102 18935 7158 18944
rect 7116 18902 7144 18935
rect 7104 18896 7156 18902
rect 7104 18838 7156 18844
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18222 7144 18566
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 6748 18006 7052 18034
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13938 6408 14214
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6380 13546 6408 13874
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6276 13524 6328 13530
rect 6380 13518 6592 13546
rect 6276 13466 6328 13472
rect 6196 12986 6224 13466
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6564 12374 6592 13518
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6656 11558 6684 11698
rect 6748 11694 6776 18006
rect 7208 17898 7236 19366
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 6932 17870 7236 17898
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 16998 6868 17614
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6840 11082 6868 12242
rect 6932 11626 6960 17870
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7024 15706 7052 17682
rect 7300 17202 7328 19178
rect 7392 17218 7420 19246
rect 7288 17196 7340 17202
rect 7392 17190 7512 17218
rect 7288 17138 7340 17144
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 7116 16046 7144 16662
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7116 14618 7144 15982
rect 7208 15638 7236 16594
rect 7300 16454 7328 17138
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15706 7328 15846
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7012 14544 7064 14550
rect 7064 14492 7144 14498
rect 7012 14486 7144 14492
rect 7024 14470 7144 14486
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 13258 7052 13806
rect 7116 13734 7144 14470
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7116 13138 7144 13670
rect 7024 13110 7144 13138
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6932 10198 6960 11154
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 7024 9450 7052 13110
rect 7104 12232 7156 12238
rect 7102 12200 7104 12209
rect 7156 12200 7158 12209
rect 7102 12135 7158 12144
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11762 7144 12038
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7116 11014 7144 11494
rect 7208 11218 7236 13126
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 11898 7328 12582
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7116 9926 7144 10474
rect 7392 10169 7420 16186
rect 7484 15366 7512 17190
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 14482 7512 14758
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7484 13938 7512 14418
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7668 13870 7696 20318
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8220 18766 8248 19110
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8128 18426 8156 18702
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7760 16114 7788 18022
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17218 8248 18702
rect 8404 18086 8432 22320
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8496 17338 8524 18702
rect 8772 18630 8800 19178
rect 8760 18624 8812 18630
rect 8574 18592 8630 18601
rect 8760 18566 8812 18572
rect 8574 18527 8630 18536
rect 8588 18086 8616 18527
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8036 17190 8248 17218
rect 8392 17196 8444 17202
rect 8036 17134 8064 17190
rect 8392 17138 8444 17144
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8220 16658 8248 16934
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 16114 8248 16594
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8312 15502 8340 16390
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8312 14958 8340 15438
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7760 13530 7788 14418
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7760 13394 7788 13466
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7576 11694 7604 12106
rect 7668 11694 7696 12718
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7668 11150 7696 11630
rect 8220 11626 8248 12174
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8206 11248 8262 11257
rect 7932 11212 7984 11218
rect 8206 11183 8208 11192
rect 7932 11154 7984 11160
rect 8260 11183 8262 11192
rect 8208 11154 8260 11160
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7378 10160 7434 10169
rect 7378 10095 7434 10104
rect 7668 10062 7696 11086
rect 7944 10742 7972 11154
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7656 10056 7708 10062
rect 8312 10033 8340 14418
rect 8404 13297 8432 17138
rect 8680 16182 8708 18362
rect 8772 18290 8800 18566
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8864 18222 8892 22320
rect 9324 20058 9352 22320
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9692 19310 9720 19858
rect 9784 19802 9812 22320
rect 9956 19848 10008 19854
rect 9784 19774 9904 19802
rect 9956 19790 10008 19796
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18698 9260 19110
rect 9784 18834 9812 19654
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 8942 18320 8998 18329
rect 8942 18255 8944 18264
rect 8996 18255 8998 18264
rect 8944 18226 8996 18232
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8680 13326 8708 13738
rect 8484 13320 8536 13326
rect 8390 13288 8446 13297
rect 8484 13262 8536 13268
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8390 13223 8446 13232
rect 8496 12442 8524 13262
rect 8680 12986 8708 13262
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8496 10810 8524 12242
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8576 10056 8628 10062
rect 7656 9998 7708 10004
rect 8298 10024 8354 10033
rect 7668 9926 7696 9998
rect 8576 9998 8628 10004
rect 8298 9959 8354 9968
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7116 9586 7144 9862
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7668 9450 7696 9862
rect 7944 9518 7972 9862
rect 8588 9722 8616 9998
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 6012 9302 6132 9330
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5920 8378 5948 8774
rect 5736 8362 5948 8378
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5724 8356 5948 8362
rect 5776 8350 5948 8356
rect 5724 8298 5776 8304
rect 5552 8106 5580 8298
rect 5552 8078 5672 8106
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5184 7342 5212 7822
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5552 2038 5580 7210
rect 5644 2582 5672 8078
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5736 1766 5764 8298
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6012 7546 6040 7890
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6104 7342 6132 9302
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6196 6458 6224 9318
rect 7208 9178 7236 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7208 8498 7236 8910
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 7750 7236 8434
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 6748 7546 6776 7686
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 7300 6730 7328 9318
rect 7484 9042 7512 9318
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7668 8974 7696 9386
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8772 9042 8800 18022
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8864 16522 8892 17070
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8864 16114 8892 16458
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8864 15162 8892 16050
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8864 13870 8892 15098
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 9048 12442 9076 18022
rect 9692 17898 9720 18158
rect 9508 17870 9720 17898
rect 9508 17134 9536 17870
rect 9876 17814 9904 19774
rect 9968 19378 9996 19790
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9954 18864 10010 18873
rect 9954 18799 10010 18808
rect 9968 18426 9996 18799
rect 10060 18766 10088 19246
rect 10244 18884 10272 22320
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10152 18856 10272 18884
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 10060 18222 10088 18702
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9678 17096 9734 17105
rect 9678 17031 9734 17040
rect 9692 16998 9720 17031
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9784 16794 9812 17682
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9876 17066 9904 17614
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9876 15502 9904 15914
rect 9968 15570 9996 18090
rect 10152 15706 10180 18856
rect 10336 18426 10364 19246
rect 10428 19174 10456 19790
rect 10704 19394 10732 22320
rect 10612 19366 10732 19394
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10428 18834 10456 19110
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10336 17678 10364 18090
rect 10612 18086 10640 19366
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10336 17338 10364 17614
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10244 16250 10272 17002
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10428 16046 10456 16390
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9876 15162 9904 15438
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 10244 14958 10272 15438
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 9692 14074 9720 14894
rect 10230 14512 10286 14521
rect 10428 14482 10456 15982
rect 10230 14447 10232 14456
rect 10284 14447 10286 14456
rect 10416 14476 10468 14482
rect 10232 14418 10284 14424
rect 10416 14418 10468 14424
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10428 12986 10456 13874
rect 10796 13462 10824 18770
rect 11058 18184 11114 18193
rect 11058 18119 11114 18128
rect 11072 14958 11100 18119
rect 11164 17542 11192 22320
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 17338 11652 22320
rect 11992 20074 12020 22320
rect 11716 20046 12020 20074
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 15502 11652 15846
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11072 13938 11100 14758
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11164 13802 11192 15302
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11624 15026 11652 15438
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 14550 11652 14962
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11624 13938 11652 14214
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9140 12238 9168 12650
rect 10060 12306 10088 12718
rect 10428 12374 10456 12922
rect 11072 12918 11100 13670
rect 11256 13530 11284 13738
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11624 12782 11652 13874
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11898 9168 12174
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 10606 8892 11494
rect 9048 11354 9076 11562
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 10060 10674 10088 12242
rect 10416 12232 10468 12238
rect 10414 12200 10416 12209
rect 10468 12200 10470 12209
rect 10414 12135 10470 12144
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11762 10548 12038
rect 11164 11898 11192 12242
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 10520 11218 10548 11698
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 11624 11082 11652 11698
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7852 8634 7880 8978
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7852 8514 7880 8570
rect 7760 8486 7880 8514
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 7002 7604 7142
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7760 6798 7788 8486
rect 8772 8430 8800 8978
rect 8864 8430 8892 10542
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9692 9178 9720 10134
rect 10704 10130 10732 10610
rect 11624 10538 11652 11018
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10336 9654 10364 10066
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 10888 8974 10916 9522
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8220 7886 8248 8298
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8864 8090 8892 8230
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7750 8248 7822
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8220 7410 8248 7686
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8496 6866 8524 7686
rect 8772 7342 8800 8026
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8680 6866 8708 7278
rect 8864 7002 8892 7890
rect 8956 7478 8984 7890
rect 9140 7818 9168 8434
rect 11716 8430 11744 20046
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11992 18902 12020 19858
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12176 18902 12204 19246
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 12164 18896 12216 18902
rect 12452 18873 12480 22320
rect 12912 20058 12940 22320
rect 13372 20058 13400 22320
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13004 19378 13032 19858
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 12164 18838 12216 18844
rect 12438 18864 12494 18873
rect 11796 18828 11848 18834
rect 12438 18799 12494 18808
rect 12532 18828 12584 18834
rect 11796 18770 11848 18776
rect 12532 18770 12584 18776
rect 11808 14074 11836 18770
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11900 16454 11928 17138
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 16046 11928 16390
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 8022 9444 8230
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 9140 7410 9168 7754
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 9140 6798 9168 7346
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 8772 6458 8800 6734
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 5724 1760 5776 1766
rect 5724 1702 5776 1708
rect 5828 1086 5856 6394
rect 9232 6225 9260 6734
rect 9692 6662 9720 6734
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 9218 6216 9274 6225
rect 9218 6151 9274 6160
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 5816 1080 5868 1086
rect 5816 1022 5868 1028
rect 11808 626 11836 13874
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11992 12442 12020 12582
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 11762 11928 12038
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12084 11234 12112 17478
rect 12544 17338 12572 18770
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15706 12204 15846
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 11992 11206 12112 11234
rect 11992 10470 12020 11206
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 10810 12112 11018
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 12084 10198 12112 10746
rect 12176 10606 12204 10950
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 12268 9450 12296 17274
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12346 16008 12402 16017
rect 12346 15943 12402 15952
rect 12360 15570 12388 15943
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12452 15502 12480 16594
rect 12820 16250 12848 16934
rect 12912 16794 12940 16934
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12912 16454 12940 16594
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 13004 16402 13032 16662
rect 13084 16448 13136 16454
rect 13004 16396 13084 16402
rect 13004 16390 13136 16396
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12530 16008 12586 16017
rect 12912 15994 12940 16390
rect 13004 16374 13124 16390
rect 13004 16114 13032 16374
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12912 15966 13124 15994
rect 12530 15943 12586 15952
rect 12544 15910 12572 15943
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12360 11286 12388 14894
rect 12544 13802 12572 15506
rect 13096 15366 13124 15966
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13096 14482 13124 15302
rect 13188 15162 13216 19246
rect 13372 18970 13400 19858
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17678 13584 18022
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13372 17134 13400 17614
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 15638 13308 16934
rect 13556 16658 13584 17614
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13544 15700 13596 15706
rect 13648 15688 13676 15846
rect 13596 15660 13676 15688
rect 13544 15642 13596 15648
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 13938 13308 14418
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 13280 13530 13308 13874
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13372 13394 13400 13874
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12544 12374 12572 12718
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12360 10810 12388 11222
rect 12728 11082 12756 13262
rect 13372 12730 13400 13330
rect 13464 12986 13492 14758
rect 13556 14074 13584 14758
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13648 12850 13676 13466
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13372 12702 13676 12730
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13556 12442 13584 12582
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13556 12209 13584 12242
rect 13648 12238 13676 12702
rect 13636 12232 13688 12238
rect 13542 12200 13598 12209
rect 12808 12164 12860 12170
rect 13636 12174 13688 12180
rect 13542 12135 13598 12144
rect 12808 12106 12860 12112
rect 12820 11694 12848 12106
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 13096 11218 13124 12038
rect 13648 11762 13676 12174
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12728 10606 12756 11018
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12728 10130 12756 10542
rect 13096 10266 13124 10542
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 13280 10062 13308 11290
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13372 10266 13400 10474
rect 13740 10266 13768 19246
rect 13832 19174 13860 22320
rect 14292 19786 14320 22320
rect 14752 20244 14780 22320
rect 14752 20216 15056 20244
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14372 19916 14424 19922
rect 14372 19858 14424 19864
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 14384 19378 14412 19858
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13924 18986 13952 19178
rect 13832 18958 13952 18986
rect 13832 15570 13860 18958
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 13734 13860 15506
rect 13924 15502 13952 18838
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14016 17338 14044 18770
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 13870 13952 15438
rect 13912 13864 13964 13870
rect 13964 13812 14044 13818
rect 13912 13806 14044 13812
rect 13924 13790 14044 13806
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13326 13860 13670
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 14016 12442 14044 13790
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13832 11694 13860 12174
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 14016 11626 14044 12378
rect 14108 11898 14136 19246
rect 15028 19174 15056 20216
rect 15212 20058 15240 22320
rect 15672 20058 15700 22320
rect 16132 20058 16160 22320
rect 16592 20058 16620 22320
rect 17052 20058 17080 22320
rect 17512 20058 17540 22320
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17500 20052 17552 20058
rect 17972 20040 18000 22320
rect 18432 20058 18460 22320
rect 18892 20058 18920 22320
rect 17500 19994 17552 20000
rect 17880 20012 18000 20040
rect 18420 20052 18472 20058
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 15212 19310 15240 19858
rect 16132 19378 16160 19858
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 16250 14228 16594
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14292 15706 14320 16526
rect 14384 16114 14412 18158
rect 14476 17542 14504 18770
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 14568 18086 14596 18702
rect 15212 18426 15240 18702
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15016 18216 15068 18222
rect 15014 18184 15016 18193
rect 15068 18184 15070 18193
rect 15014 18119 15070 18128
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14568 17814 14596 18022
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14384 14482 14412 16050
rect 14476 16046 14504 17478
rect 14568 16114 14596 17478
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14476 13530 14504 15506
rect 14568 15502 14596 16050
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15028 15570 15056 16118
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14556 15496 14608 15502
rect 15120 15450 15148 15982
rect 14556 15438 14608 15444
rect 15028 15422 15148 15450
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14568 14618 14596 14894
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 15028 13802 15056 15422
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15120 13870 15148 14418
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14476 12306 14504 13466
rect 15396 12782 15424 19246
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15474 18728 15530 18737
rect 15474 18663 15530 18672
rect 15488 18086 15516 18663
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 14804 15516 18022
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15580 16522 15608 17614
rect 15672 17338 15700 18770
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15580 16114 15608 16458
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15672 15162 15700 17138
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15568 14816 15620 14822
rect 15488 14776 15568 14804
rect 15568 14758 15620 14764
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 15384 12232 15436 12238
rect 15488 12186 15516 12718
rect 15436 12180 15516 12186
rect 15384 12174 15516 12180
rect 15396 12158 15516 12174
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 15488 11830 15516 12158
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15580 11694 15608 14758
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15672 14521 15700 14554
rect 15658 14512 15714 14521
rect 15658 14447 15714 14456
rect 15764 13530 15792 19246
rect 16592 18902 16620 19858
rect 17144 19378 17172 19858
rect 17880 19446 17908 20012
rect 18420 19994 18472 20000
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15856 17746 15884 18226
rect 15948 18154 15976 18702
rect 15936 18148 15988 18154
rect 15936 18090 15988 18096
rect 15948 17882 15976 18090
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15856 17202 15884 17682
rect 15948 17338 15976 17818
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 15502 15884 16934
rect 16224 16674 16252 17070
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16316 16794 16344 16934
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16224 16646 16344 16674
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16040 15434 16068 16050
rect 16316 15994 16344 16646
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16132 15978 16344 15994
rect 16120 15972 16344 15978
rect 16172 15966 16344 15972
rect 16120 15914 16172 15920
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 16040 15026 16068 15370
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 13870 15976 14350
rect 16040 14074 16068 14962
rect 16316 14074 16344 15966
rect 16408 15706 16436 16526
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15672 11898 15700 12310
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 14568 11354 14596 11630
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15304 11354 15332 11494
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14568 10810 14596 11086
rect 15396 11014 15424 11494
rect 15764 11354 15792 13262
rect 16132 11898 16160 13262
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 15672 10606 15700 11154
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 14016 9586 14044 10066
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 16132 9450 16160 10610
rect 16224 10130 16252 11766
rect 16500 10810 16528 18702
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16592 15502 16620 15914
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16684 13530 16712 18770
rect 16776 16726 16804 19246
rect 17972 18970 18000 19858
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 18064 19174 18092 19382
rect 18524 19378 18552 19858
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16868 15910 16896 18090
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 13546 16896 15846
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16960 14074 16988 14826
rect 17052 14618 17080 18838
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17972 17882 18000 18770
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17134 17908 17478
rect 17972 17338 18000 17614
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 18418 17096 18474 17105
rect 18418 17031 18420 17040
rect 18472 17031 18474 17040
rect 18420 17002 18472 17008
rect 18524 16794 18552 17614
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17236 16250 17264 16594
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17420 15162 17448 15438
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16776 13518 16896 13546
rect 16776 13410 16804 13518
rect 16684 13382 16804 13410
rect 16960 13394 16988 14010
rect 17052 13462 17080 14350
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17144 13530 17172 14282
rect 17512 14074 17540 14350
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16856 13388 16908 13394
rect 16684 12306 16712 13382
rect 16856 13330 16908 13336
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16776 12714 16804 13262
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16776 12442 16804 12650
rect 16868 12442 16896 13330
rect 17236 12986 17264 13806
rect 17972 13802 18000 14486
rect 18064 14482 18092 14894
rect 18524 14890 18552 16730
rect 18616 16726 18644 17138
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 18708 14804 18736 19246
rect 18892 18766 18920 19858
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19076 18902 19104 19246
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 19352 18170 19380 22320
rect 19352 18142 19748 18170
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 19076 17202 19104 17682
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 18616 14776 18736 14804
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18616 13818 18644 14776
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18708 13938 18736 14486
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11694 17356 12038
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17788 11354 17816 12310
rect 17972 11830 18000 12718
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9518 16252 10066
rect 16868 9586 16896 10406
rect 17052 10130 17080 10610
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17052 9722 17080 10066
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 12360 9110 12388 9386
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 17604 8294 17632 11018
rect 17972 10674 18000 11766
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 11354 18184 11494
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18524 9382 18552 13806
rect 18616 13790 18736 13818
rect 18708 12442 18736 13790
rect 18800 12782 18828 14214
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 11642 19288 12174
rect 19168 11614 19288 11642
rect 19168 11558 19196 11614
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19168 10606 19196 11494
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 19352 7546 19380 17274
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19536 14550 19564 14758
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 12306 19472 12582
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11694 19472 12242
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19444 11150 19472 11630
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 18984 6934 19012 7278
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19260 6662 19288 6802
rect 19628 6730 19656 18022
rect 19720 8090 19748 18142
rect 19812 17338 19840 22320
rect 20272 18086 20300 22320
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20640 18698 20668 19178
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 20732 17066 20760 22320
rect 21192 17218 21220 22320
rect 20824 17190 21220 17218
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19996 11529 20024 11562
rect 19982 11520 20038 11529
rect 19982 11455 20038 11464
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 20824 5914 20852 17190
rect 21652 17134 21680 22320
rect 22112 19310 22140 22320
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22572 18154 22600 22320
rect 22560 18148 22612 18154
rect 22560 18090 22612 18096
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 20916 5370 20944 17070
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 21008 6458 21036 17002
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 11440 598 11836 626
rect 11440 480 11468 598
rect 3240 468 3292 474
rect 3240 410 3292 416
rect 4988 468 5040 474
rect 4988 410 5040 416
rect 3252 241 3280 410
rect 3238 232 3294 241
rect 3238 167 3294 176
rect 11426 0 11482 480
<< via2 >>
rect 1398 22480 1454 22536
rect 1582 20168 1638 20224
rect 1490 19080 1546 19136
rect 1858 19760 1914 19816
rect 1766 17856 1822 17912
rect 1674 16940 1676 16960
rect 1676 16940 1728 16960
rect 1728 16940 1730 16960
rect 1674 16904 1730 16940
rect 1674 16516 1730 16552
rect 1674 16496 1676 16516
rect 1676 16496 1728 16516
rect 1728 16496 1730 16516
rect 1766 15952 1822 16008
rect 1490 14048 1546 14104
rect 1582 13640 1638 13696
rect 1950 18264 2006 18320
rect 2226 18264 2282 18320
rect 3054 22072 3110 22128
rect 2962 21528 3018 21584
rect 2870 21120 2926 21176
rect 2778 20576 2834 20632
rect 2594 19216 2650 19272
rect 2410 17992 2466 18048
rect 2502 17312 2558 17368
rect 2042 14592 2098 14648
rect 2962 18808 3018 18864
rect 2778 18128 2834 18184
rect 2870 15544 2926 15600
rect 2778 14728 2834 14784
rect 3238 18944 3294 19000
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4526 18672 4582 18728
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4434 18028 4436 18048
rect 4436 18028 4488 18048
rect 4488 18028 4490 18048
rect 4434 17992 4490 18028
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3238 12144 3294 12200
rect 3422 10104 3478 10160
rect 3422 9424 3478 9480
rect 3238 4256 3294 4312
rect 2778 2524 2780 2544
rect 2780 2524 2832 2544
rect 2832 2524 2834 2544
rect 2778 2488 2834 2524
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4066 12688 4122 12744
rect 4066 12316 4068 12336
rect 4068 12316 4120 12336
rect 4120 12316 4122 12336
rect 4066 12280 4122 12316
rect 4250 12280 4306 12336
rect 4710 12316 4712 12336
rect 4712 12316 4764 12336
rect 4764 12316 4766 12336
rect 4710 12280 4766 12316
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 11736 4122 11792
rect 3974 10784 4030 10840
rect 4066 10376 4122 10432
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 3882 9016 3938 9072
rect 4066 8472 4122 8528
rect 4066 8064 4122 8120
rect 3790 7520 3846 7576
rect 4066 7112 4122 7168
rect 4066 6704 4122 6760
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 3974 5752 4030 5808
rect 4066 5208 4122 5264
rect 4066 4800 4122 4856
rect 3882 3440 3938 3496
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4250 3848 4306 3904
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 3974 2896 4030 2952
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 3698 1980 3700 2000
rect 3700 1980 3752 2000
rect 3752 1980 3754 2000
rect 3698 1944 3754 1980
rect 3698 1536 3754 1592
rect 4066 1028 4068 1048
rect 4068 1028 4120 1048
rect 4120 1028 4122 1048
rect 4066 992 4122 1028
rect 3606 584 3662 640
rect 7102 18944 7158 19000
rect 7102 12180 7104 12200
rect 7104 12180 7156 12200
rect 7156 12180 7158 12200
rect 7102 12144 7158 12180
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8574 18536 8630 18592
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8206 11212 8262 11248
rect 8206 11192 8208 11212
rect 8208 11192 8260 11212
rect 8260 11192 8262 11212
rect 7378 10104 7434 10160
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8942 18284 8998 18320
rect 8942 18264 8944 18284
rect 8944 18264 8996 18284
rect 8996 18264 8998 18284
rect 8390 13232 8446 13288
rect 8298 9968 8354 10024
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 9954 18808 10010 18864
rect 9678 17040 9734 17096
rect 10230 14476 10286 14512
rect 10230 14456 10232 14476
rect 10232 14456 10284 14476
rect 10284 14456 10286 14476
rect 11058 18128 11114 18184
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 10414 12180 10416 12200
rect 10416 12180 10468 12200
rect 10468 12180 10470 12200
rect 10414 12144 10470 12180
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 12438 18808 12494 18864
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 9218 6160 9274 6216
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12346 15952 12402 16008
rect 12530 15952 12586 16008
rect 13542 12144 13598 12200
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 15014 18164 15016 18184
rect 15016 18164 15068 18184
rect 15068 18164 15070 18184
rect 15014 18128 15070 18164
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 15474 18672 15530 18728
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 15658 14456 15714 14512
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18418 17060 18474 17096
rect 18418 17040 18420 17060
rect 18420 17040 18472 17060
rect 18472 17040 18474 17060
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 19982 11464 20038 11520
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 3238 176 3294 232
<< metal3 >>
rect 0 22538 480 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 480 22478
rect 1393 22475 1459 22478
rect 0 22130 480 22160
rect 3049 22130 3115 22133
rect 0 22128 3115 22130
rect 0 22072 3054 22128
rect 3110 22072 3115 22128
rect 0 22070 3115 22072
rect 0 22040 480 22070
rect 3049 22067 3115 22070
rect 0 21586 480 21616
rect 2957 21586 3023 21589
rect 0 21584 3023 21586
rect 0 21528 2962 21584
rect 3018 21528 3023 21584
rect 0 21526 3023 21528
rect 0 21496 480 21526
rect 2957 21523 3023 21526
rect 0 21178 480 21208
rect 2865 21178 2931 21181
rect 0 21176 2931 21178
rect 0 21120 2870 21176
rect 2926 21120 2931 21176
rect 0 21118 2931 21120
rect 0 21088 480 21118
rect 2865 21115 2931 21118
rect 0 20634 480 20664
rect 2773 20634 2839 20637
rect 0 20632 2839 20634
rect 0 20576 2778 20632
rect 2834 20576 2839 20632
rect 0 20574 2839 20576
rect 0 20544 480 20574
rect 2773 20571 2839 20574
rect 0 20226 480 20256
rect 1577 20226 1643 20229
rect 0 20224 1643 20226
rect 0 20168 1582 20224
rect 1638 20168 1643 20224
rect 0 20166 1643 20168
rect 0 20136 480 20166
rect 1577 20163 1643 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 480 19758
rect 1853 19755 1919 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 2589 19274 2655 19277
rect 0 19272 2655 19274
rect 0 19216 2594 19272
rect 2650 19216 2655 19272
rect 0 19214 2655 19216
rect 0 19184 480 19214
rect 2589 19211 2655 19214
rect 1485 19138 1551 19141
rect 1485 19136 7482 19138
rect 1485 19080 1490 19136
rect 1546 19080 7482 19136
rect 1485 19078 7482 19080
rect 1485 19075 1551 19078
rect 3233 19002 3299 19005
rect 7097 19002 7163 19005
rect 3233 19000 7163 19002
rect 3233 18944 3238 19000
rect 3294 18944 7102 19000
rect 7158 18944 7163 19000
rect 3233 18942 7163 18944
rect 3233 18939 3299 18942
rect 7097 18939 7163 18942
rect 0 18866 480 18896
rect 2957 18866 3023 18869
rect 0 18864 3023 18866
rect 0 18808 2962 18864
rect 3018 18808 3023 18864
rect 0 18806 3023 18808
rect 0 18776 480 18806
rect 2957 18803 3023 18806
rect 4521 18730 4587 18733
rect 7422 18730 7482 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 9949 18866 10015 18869
rect 12433 18866 12499 18869
rect 9949 18864 12499 18866
rect 9949 18808 9954 18864
rect 10010 18808 12438 18864
rect 12494 18808 12499 18864
rect 9949 18806 12499 18808
rect 9949 18803 10015 18806
rect 12433 18803 12499 18806
rect 15469 18730 15535 18733
rect 4521 18728 4906 18730
rect 4521 18672 4526 18728
rect 4582 18672 4906 18728
rect 4521 18670 4906 18672
rect 7422 18728 15535 18730
rect 7422 18672 15474 18728
rect 15530 18672 15535 18728
rect 7422 18670 15535 18672
rect 4521 18667 4587 18670
rect 4846 18594 4906 18670
rect 15469 18667 15535 18670
rect 8569 18594 8635 18597
rect 4846 18592 8635 18594
rect 4846 18536 8574 18592
rect 8630 18536 8635 18592
rect 4846 18534 8635 18536
rect 8569 18531 8635 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 480 18262
rect 1945 18259 2011 18262
rect 2221 18322 2287 18325
rect 8937 18322 9003 18325
rect 2221 18320 9003 18322
rect 2221 18264 2226 18320
rect 2282 18264 8942 18320
rect 8998 18264 9003 18320
rect 2221 18262 9003 18264
rect 2221 18259 2287 18262
rect 8937 18259 9003 18262
rect 2773 18186 2839 18189
rect 11053 18186 11119 18189
rect 15009 18186 15075 18189
rect 2773 18184 15075 18186
rect 2773 18128 2778 18184
rect 2834 18128 11058 18184
rect 11114 18128 15014 18184
rect 15070 18128 15075 18184
rect 2773 18126 15075 18128
rect 2773 18123 2839 18126
rect 11053 18123 11119 18126
rect 15009 18123 15075 18126
rect 2405 18050 2471 18053
rect 4429 18050 4495 18053
rect 2405 18048 4495 18050
rect 2405 17992 2410 18048
rect 2466 17992 4434 18048
rect 4490 17992 4495 18048
rect 2405 17990 4495 17992
rect 2405 17987 2471 17990
rect 4429 17987 4495 17990
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1761 17914 1827 17917
rect 0 17912 1827 17914
rect 0 17856 1766 17912
rect 1822 17856 1827 17912
rect 0 17854 1827 17856
rect 0 17824 480 17854
rect 1761 17851 1827 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 2497 17370 2563 17373
rect 0 17368 2563 17370
rect 0 17312 2502 17368
rect 2558 17312 2563 17368
rect 0 17310 2563 17312
rect 0 17280 480 17310
rect 2497 17307 2563 17310
rect 9673 17098 9739 17101
rect 18413 17098 18479 17101
rect 9673 17096 18479 17098
rect 9673 17040 9678 17096
rect 9734 17040 18418 17096
rect 18474 17040 18479 17096
rect 9673 17038 18479 17040
rect 9673 17035 9739 17038
rect 18413 17035 18479 17038
rect 0 16962 480 16992
rect 1669 16962 1735 16965
rect 0 16960 1735 16962
rect 0 16904 1674 16960
rect 1730 16904 1735 16960
rect 0 16902 1735 16904
rect 0 16872 480 16902
rect 1669 16899 1735 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 1669 16554 1735 16557
rect 0 16552 1735 16554
rect 0 16496 1674 16552
rect 1730 16496 1735 16552
rect 0 16494 1735 16496
rect 0 16464 480 16494
rect 1669 16491 1735 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1761 16010 1827 16013
rect 0 16008 1827 16010
rect 0 15952 1766 16008
rect 1822 15952 1827 16008
rect 0 15950 1827 15952
rect 0 15920 480 15950
rect 1761 15947 1827 15950
rect 12341 16010 12407 16013
rect 12525 16010 12591 16013
rect 12341 16008 12591 16010
rect 12341 15952 12346 16008
rect 12402 15952 12530 16008
rect 12586 15952 12591 16008
rect 12341 15950 12591 15952
rect 12341 15947 12407 15950
rect 12525 15947 12591 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 2865 15602 2931 15605
rect 0 15600 2931 15602
rect 0 15544 2870 15600
rect 2926 15544 2931 15600
rect 0 15542 2931 15544
rect 0 15512 480 15542
rect 2865 15539 2931 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 0 14998 674 15058
rect 0 14968 480 14998
rect 614 14786 674 14998
rect 2773 14786 2839 14789
rect 614 14784 2839 14786
rect 614 14728 2778 14784
rect 2834 14728 2839 14784
rect 614 14726 2839 14728
rect 2773 14723 2839 14726
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 2037 14650 2103 14653
rect 0 14648 2103 14650
rect 0 14592 2042 14648
rect 2098 14592 2103 14648
rect 0 14590 2103 14592
rect 0 14560 480 14590
rect 2037 14587 2103 14590
rect 10225 14514 10291 14517
rect 15653 14514 15719 14517
rect 10225 14512 15719 14514
rect 10225 14456 10230 14512
rect 10286 14456 15658 14512
rect 15714 14456 15719 14512
rect 10225 14454 15719 14456
rect 10225 14451 10291 14454
rect 15653 14451 15719 14454
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1485 14106 1551 14109
rect 0 14104 1551 14106
rect 0 14048 1490 14104
rect 1546 14048 1551 14104
rect 0 14046 1551 14048
rect 0 14016 480 14046
rect 1485 14043 1551 14046
rect 0 13698 480 13728
rect 1577 13698 1643 13701
rect 0 13696 1643 13698
rect 0 13640 1582 13696
rect 1638 13640 1643 13696
rect 0 13638 1643 13640
rect 0 13608 480 13638
rect 1577 13635 1643 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 8385 13290 8451 13293
rect 0 13288 8451 13290
rect 0 13232 8390 13288
rect 8446 13232 8451 13288
rect 0 13230 8451 13232
rect 0 13200 480 13230
rect 8385 13227 8451 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 480 12686
rect 4061 12683 4127 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 4245 12338 4311 12341
rect 4705 12338 4771 12341
rect 4245 12336 4771 12338
rect 4245 12280 4250 12336
rect 4306 12280 4710 12336
rect 4766 12280 4771 12336
rect 4245 12278 4771 12280
rect 4245 12275 4311 12278
rect 4705 12275 4771 12278
rect 3233 12202 3299 12205
rect 7097 12202 7163 12205
rect 3233 12200 7163 12202
rect 3233 12144 3238 12200
rect 3294 12144 7102 12200
rect 7158 12144 7163 12200
rect 3233 12142 7163 12144
rect 3233 12139 3299 12142
rect 7097 12139 7163 12142
rect 10409 12202 10475 12205
rect 13537 12202 13603 12205
rect 10409 12200 13603 12202
rect 10409 12144 10414 12200
rect 10470 12144 13542 12200
rect 13598 12144 13603 12200
rect 10409 12142 13603 12144
rect 10409 12139 10475 12142
rect 13537 12139 13603 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 480 11734
rect 4061 11731 4127 11734
rect 19977 11522 20043 11525
rect 22320 11522 22800 11552
rect 19977 11520 22800 11522
rect 19977 11464 19982 11520
rect 20038 11464 22800 11520
rect 19977 11462 22800 11464
rect 19977 11459 20043 11462
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 22320 11432 22800 11462
rect 14672 11391 14992 11392
rect 0 11326 4906 11386
rect 0 11296 480 11326
rect 4846 11250 4906 11326
rect 8201 11250 8267 11253
rect 4846 11248 8267 11250
rect 4846 11192 8206 11248
rect 8262 11192 8267 11248
rect 4846 11190 8267 11192
rect 8201 11187 8267 11190
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3969 10842 4035 10845
rect 0 10840 4035 10842
rect 0 10784 3974 10840
rect 4030 10784 4035 10840
rect 0 10782 4035 10784
rect 0 10752 480 10782
rect 3969 10779 4035 10782
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 3417 10162 3483 10165
rect 7373 10162 7439 10165
rect 3417 10160 7439 10162
rect 3417 10104 3422 10160
rect 3478 10104 7378 10160
rect 7434 10104 7439 10160
rect 3417 10102 7439 10104
rect 3417 10099 3483 10102
rect 7373 10099 7439 10102
rect 0 10026 480 10056
rect 8293 10026 8359 10029
rect 0 10024 8359 10026
rect 0 9968 8298 10024
rect 8354 9968 8359 10024
rect 0 9966 8359 9968
rect 0 9936 480 9966
rect 8293 9963 8359 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 0 9482 480 9512
rect 3417 9482 3483 9485
rect 0 9480 3483 9482
rect 0 9424 3422 9480
rect 3478 9424 3483 9480
rect 0 9422 3483 9424
rect 0 9392 480 9422
rect 3417 9419 3483 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 3877 9074 3943 9077
rect 0 9072 3943 9074
rect 0 9016 3882 9072
rect 3938 9016 3943 9072
rect 0 9014 3943 9016
rect 0 8984 480 9014
rect 3877 9011 3943 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 480 8470
rect 4061 8467 4127 8470
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 480 8062
rect 4061 8059 4127 8062
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3785 7578 3851 7581
rect 0 7576 3851 7578
rect 0 7520 3790 7576
rect 3846 7520 3851 7576
rect 0 7518 3851 7520
rect 0 7488 480 7518
rect 3785 7515 3851 7518
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 480 6702
rect 4061 6699 4127 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 480 6248
rect 9213 6218 9279 6221
rect 0 6216 9279 6218
rect 0 6160 9218 6216
rect 9274 6160 9279 6216
rect 0 6158 9279 6160
rect 0 6128 480 6158
rect 9213 6155 9279 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 3969 5810 4035 5813
rect 0 5808 4035 5810
rect 0 5752 3974 5808
rect 4030 5752 4035 5808
rect 0 5750 4035 5752
rect 0 5720 480 5750
rect 3969 5747 4035 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 480 5206
rect 4061 5203 4127 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 480 4798
rect 4061 4795 4127 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 3233 4314 3299 4317
rect 0 4312 3299 4314
rect 0 4256 3238 4312
rect 3294 4256 3299 4312
rect 0 4254 3299 4256
rect 0 4224 480 4254
rect 3233 4251 3299 4254
rect 0 3906 480 3936
rect 4245 3906 4311 3909
rect 0 3904 4311 3906
rect 0 3848 4250 3904
rect 4306 3848 4311 3904
rect 0 3846 4311 3848
rect 0 3816 480 3846
rect 4245 3843 4311 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 0 3498 480 3528
rect 3877 3498 3943 3501
rect 0 3496 3943 3498
rect 0 3440 3882 3496
rect 3938 3440 3943 3496
rect 0 3438 3943 3440
rect 0 3408 480 3438
rect 3877 3435 3943 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 480 2984
rect 3969 2954 4035 2957
rect 0 2952 4035 2954
rect 0 2896 3974 2952
rect 4030 2896 4035 2952
rect 0 2894 4035 2896
rect 0 2864 480 2894
rect 3969 2891 4035 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 2773 2546 2839 2549
rect 0 2544 2839 2546
rect 0 2488 2778 2544
rect 2834 2488 2839 2544
rect 0 2486 2839 2488
rect 0 2456 480 2486
rect 2773 2483 2839 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 3693 2002 3759 2005
rect 0 2000 3759 2002
rect 0 1944 3698 2000
rect 3754 1944 3759 2000
rect 0 1942 3759 1944
rect 0 1912 480 1942
rect 3693 1939 3759 1942
rect 0 1594 480 1624
rect 3693 1594 3759 1597
rect 0 1592 3759 1594
rect 0 1536 3698 1592
rect 3754 1536 3759 1592
rect 0 1534 3759 1536
rect 0 1504 480 1534
rect 3693 1531 3759 1534
rect 0 1050 480 1080
rect 4061 1050 4127 1053
rect 0 1048 4127 1050
rect 0 992 4066 1048
rect 4122 992 4127 1048
rect 0 990 4127 992
rect 0 960 480 990
rect 4061 987 4127 990
rect 0 642 480 672
rect 3601 642 3667 645
rect 0 640 3667 642
rect 0 584 3606 640
rect 3662 584 3667 640
rect 0 582 3667 584
rect 0 552 480 582
rect 3601 579 3667 582
rect 0 234 480 264
rect 3233 234 3299 237
rect 0 232 3299 234
rect 0 176 3238 232
rect 3294 176 3299 232
rect 0 174 3299 176
rect 0 144 480 174
rect 3233 171 3299 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606256979
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606256979
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606256979
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606256979
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606256979
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606256979
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606256979
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606256979
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606256979
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1606256979
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606256979
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1606256979
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1606256979
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606256979
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606256979
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1606256979
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606256979
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1606256979
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1606256979
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606256979
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606256979
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606256979
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1606256979
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1606256979
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1606256979
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1606256979
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606256979
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1606256979
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1606256979
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1606256979
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606256979
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606256979
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606256979
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606256979
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606256979
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1606256979
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606256979
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1606256979
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1606256979
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1606256979
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606256979
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606256979
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606256979
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606256979
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606256979
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606256979
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606256979
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1606256979
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1606256979
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1606256979
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1606256979
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1606256979
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1606256979
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1606256979
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606256979
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606256979
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606256979
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606256979
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606256979
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1606256979
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1606256979
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1606256979
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1606256979
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1606256979
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1606256979
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1606256979
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp 1606256979
transform 1 0 20240 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1606256979
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606256979
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606256979
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606256979
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606256979
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606256979
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606256979
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606256979
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606256979
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606256979
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606256979
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1606256979
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1606256979
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1606256979
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1606256979
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1606256979
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1606256979
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1606256979
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1606256979
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1606256979
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1606256979
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1606256979
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1606256979
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1606256979
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606256979
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606256979
transform 1 0 19872 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1606256979
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_202
timestamp 1606256979
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1606256979
transform 1 0 19136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606256979
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606256979
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606256979
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1606256979
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_46
timestamp 1606256979
transform 1 0 5336 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_58
timestamp 1606256979
transform 1 0 6440 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8280 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7176 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_75
timestamp 1606256979
transform 1 0 8004 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1606256979
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1606256979
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1606256979
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1606256979
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1606256979
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1606256979
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1606256979
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1606256979
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606256979
transform 1 0 19412 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_190
timestamp 1606256979
transform 1 0 18584 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_198
timestamp 1606256979
transform 1 0 19320 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_203
timestamp 1606256979
transform 1 0 19780 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1606256979
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606256979
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2944 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1606256979
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1606256979
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4600 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1606256979
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_54
timestamp 1606256979
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606256979
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606256979
transform 1 0 6992 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8464 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7452 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_67
timestamp 1606256979
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1606256979
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_89
timestamp 1606256979
transform 1 0 9292 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_101
timestamp 1606256979
transform 1 0 10396 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1606256979
transform 1 0 11500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1606256979
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1606256979
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1606256979
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1606256979
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1606256979
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606256979
transform 1 0 18952 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_192
timestamp 1606256979
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_198
timestamp 1606256979
transform 1 0 19320 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_210
timestamp 1606256979
transform 1 0 20424 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_218
timestamp 1606256979
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606256979
transform 1 0 1564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2116 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_9
timestamp 1606256979
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_17
timestamp 1606256979
transform 1 0 2668 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606256979
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp 1606256979
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5152 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1606256979
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8464 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_78
timestamp 1606256979
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1606256979
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1606256979
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1606256979
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1606256979
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1606256979
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1606256979
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_178
timestamp 1606256979
transform 1 0 17480 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1606256979
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606256979
transform 1 0 18400 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_192
timestamp 1606256979
transform 1 0 18768 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1606256979
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1606256979
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2116 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1606256979
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_27
timestamp 1606256979
transform 1 0 3588 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 1606256979
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1606256979
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7176 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1606256979
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1606256979
transform 1 0 9660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1606256979
transform 1 0 10764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1606256979
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606256979
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1606256979
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1606256979
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1606256979
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1606256979
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606256979
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606256979
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606256979
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_11
timestamp 1606256979
transform 1 0 2116 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4784 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1606256979
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606256979
transform 1 0 6348 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_49
timestamp 1606256979
transform 1 0 5612 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_60
timestamp 1606256979
transform 1 0 6624 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7912 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1606256979
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606256979
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_102
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_114
timestamp 1606256979
transform 1 0 11592 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_126
timestamp 1606256979
transform 1 0 12696 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_138
timestamp 1606256979
transform 1 0 13800 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1606256979
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1606256979
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1606256979
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1606256979
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1606256979
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_15
timestamp 1606256979
transform 1 0 2484 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606256979
transform 1 0 3404 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4140 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 3128 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_21
timestamp 1606256979
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_31
timestamp 1606256979
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1606256979
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1606256979
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5704 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_42
timestamp 1606256979
transform 1 0 4968 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1606256979
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_71
timestamp 1606256979
transform 1 0 7636 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_79
timestamp 1606256979
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_66
timestamp 1606256979
transform 1 0 7176 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_70
timestamp 1606256979
transform 1 0 7544 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_83
timestamp 1606256979
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10304 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_98
timestamp 1606256979
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1606256979
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11960 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_109
timestamp 1606256979
transform 1 0 11132 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1606256979
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_123
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1606256979
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1606256979
transform 1 0 11868 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606256979
transform 1 0 13340 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1606256979
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_136
timestamp 1606256979
transform 1 0 13616 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1606256979
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1606256979
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16192 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15640 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_148
timestamp 1606256979
transform 1 0 14720 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1606256979
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 1606256979
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606256979
transform 1 0 17296 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp 1606256979
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1606256979
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1606256979
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1606256979
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1606256979
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_192
timestamp 1606256979
transform 1 0 18768 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_204
timestamp 1606256979
transform 1 0 19872 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1606256979
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1606256979
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1606256979
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1606256979
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_41
timestamp 1606256979
transform 1 0 4876 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1606256979
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1606256979
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10672 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_89
timestamp 1606256979
transform 1 0 9292 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_101
timestamp 1606256979
transform 1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_123
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12972 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_145
timestamp 1606256979
transform 1 0 14444 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15456 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_153
timestamp 1606256979
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_165
timestamp 1606256979
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16468 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_176
timestamp 1606256979
transform 1 0 17296 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1606256979
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_200
timestamp 1606256979
transform 1 0 19504 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1606256979
transform 1 0 20608 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2852 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1932 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1606256979
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1606256979
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1606256979
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1606256979
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606256979
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6624 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 5520 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1606256979
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1606256979
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_59
timestamp 1606256979
transform 1 0 6532 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7636 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1606256979
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10212 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1606256979
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606256979
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_96
timestamp 1606256979
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11868 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_115
timestamp 1606256979
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 12880 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_126
timestamp 1606256979
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_131
timestamp 1606256979
transform 1 0 13156 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1606256979
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_163
timestamp 1606256979
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 17756 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606256979
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1606256979
transform 1 0 17204 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1606256979
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1606256979
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2668 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1656 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_12
timestamp 1606256979
transform 1 0 2208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_16
timestamp 1606256979
transform 1 0 2576 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_33
timestamp 1606256979
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5612 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_44
timestamp 1606256979
transform 1 0 5152 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_48
timestamp 1606256979
transform 1 0 5520 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1606256979
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7912 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_71
timestamp 1606256979
transform 1 0 7636 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606256979
transform 1 0 9660 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_90
timestamp 1606256979
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1606256979
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11132 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1606256979
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1606256979
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14444 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13432 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1606256979
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1606256979
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1606256979
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606256979
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 17112 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1606256979
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_177
timestamp 1606256979
transform 1 0 17388 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606256979
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19688 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1606256979
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1606256979
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1932 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1606256979
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1606256979
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_23
timestamp 1606256979
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5704 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1606256979
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_66
timestamp 1606256979
transform 1 0 7176 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1606256979
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10488 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606256979
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp 1606256979
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12236 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_118
timestamp 1606256979
transform 1 0 11960 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12972 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 14260 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1606256979
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_138
timestamp 1606256979
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1606256979
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606256979
transform 1 0 14536 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15364 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1606256979
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606256979
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17664 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_171
timestamp 1606256979
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1606256979
transform 1 0 17296 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18676 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_189
timestamp 1606256979
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_200
timestamp 1606256979
transform 1 0 19504 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606256979
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606256979
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1606256979
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1932 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1606256979
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606256979
transform 1 0 2300 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606256979
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_17
timestamp 1606256979
transform 1 0 2668 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606256979
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4692 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1606256979
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_33
timestamp 1606256979
transform 1 0 4140 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1606256979
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606256979
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5152 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_55
timestamp 1606256979
transform 1 0 6164 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_60
timestamp 1606256979
transform 1 0 6624 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7912 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 7176 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_71
timestamp 1606256979
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_69
timestamp 1606256979
transform 1 0 7452 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606256979
transform 1 0 9016 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10028 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_90
timestamp 1606256979
transform 1 0 9384 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_96
timestamp 1606256979
transform 1 0 9936 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1606256979
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_89
timestamp 1606256979
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11500 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10764 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1606256979
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606256979
transform 1 0 14076 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12788 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13064 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 14444 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1606256979
transform 1 0 12696 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1606256979
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_144
timestamp 1606256979
transform 1 0 14352 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_143
timestamp 1606256979
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15824 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15640 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1606256979
transform 1 0 15456 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1606256979
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606256979
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16652 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_176
timestamp 1606256979
transform 1 0 17296 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1606256979
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_167
timestamp 1606256979
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606256979
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_200
timestamp 1606256979
transform 1 0 19504 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1606256979
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1606256979
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_212
timestamp 1606256979
transform 1 0 20608 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1748 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_13
timestamp 1606256979
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 3496 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1606256979
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_42
timestamp 1606256979
transform 1 0 4968 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606256979
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8004 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1606256979
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9752 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_91
timestamp 1606256979
transform 1 0 9476 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1606256979
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12604 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1606256979
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1606256979
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1606256979
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15640 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 14628 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1606256979
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1606256979
transform 1 0 17112 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1606256979
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606256979
transform 1 0 19044 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606256979
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_198
timestamp 1606256979
transform 1 0 19320 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_210
timestamp 1606256979
transform 1 0 20424 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1606256979
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606256979
transform 1 0 1564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_9
timestamp 1606256979
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_17
timestamp 1606256979
transform 1 0 2668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606256979
transform 1 0 3312 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_23
timestamp 1606256979
transform 1 0 3220 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_41
timestamp 1606256979
transform 1 0 4876 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606256979
transform 1 0 5520 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5980 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_47
timestamp 1606256979
transform 1 0 5428 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1606256979
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 7636 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1606256979
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_74
timestamp 1606256979
transform 1 0 7912 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10396 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_86
timestamp 1606256979
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1606256979
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 13156 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_129
timestamp 1606256979
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1606256979
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1606256979
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606256979
transform 1 0 16468 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18032 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1606256979
transform 1 0 17020 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_170
timestamp 1606256979
transform 1 0 16744 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_182
timestamp 1606256979
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_200
timestamp 1606256979
transform 1 0 19504 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1606256979
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606256979
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2760 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1932 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1606256979
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_15
timestamp 1606256979
transform 1 0 2484 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_34
timestamp 1606256979
transform 1 0 4232 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5612 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_46
timestamp 1606256979
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1606256979
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8464 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1606256979
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_96
timestamp 1606256979
transform 1 0 9936 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11040 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1606256979
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1606256979
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14260 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13064 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1606256979
transform 1 0 12972 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1606256979
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16008 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_159
timestamp 1606256979
transform 1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18124 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1606256979
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1606256979
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_184
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_201
timestamp 1606256979
transform 1 0 19596 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_213
timestamp 1606256979
transform 1 0 20700 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606256979
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1932 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1606256979
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_15
timestamp 1606256979
transform 1 0 2484 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606256979
transform 1 0 3128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4692 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_21
timestamp 1606256979
transform 1 0 3036 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_25
timestamp 1606256979
transform 1 0 3404 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1606256979
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606256979
transform 1 0 6348 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1606256979
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1606256979
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1606256979
transform 1 0 8004 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8464 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_71
timestamp 1606256979
transform 1 0 7636 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1606256979
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1606256979
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_102
timestamp 1606256979
transform 1 0 10488 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12144 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11040 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_117
timestamp 1606256979
transform 1 0 11868 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 13156 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1606256979
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_134
timestamp 1606256979
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp 1606256979
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15824 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 14628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1606256979
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_169
timestamp 1606256979
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_174
timestamp 1606256979
transform 1 0 17112 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_186
timestamp 1606256979
transform 1 0 18216 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_198
timestamp 1606256979
transform 1 0 19320 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1606256979
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2576 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1840 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1606256979
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1606256979
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4232 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_32
timestamp 1606256979
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5244 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1606256979
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1606256979
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606256979
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_62
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7452 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_68
timestamp 1606256979
transform 1 0 7360 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_78
timestamp 1606256979
transform 1 0 8280 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8832 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10488 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1606256979
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1606256979
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606256979
transform 1 0 13432 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13892 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1606256979
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_137
timestamp 1606256979
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16008 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_148
timestamp 1606256979
transform 1 0 14720 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_160
timestamp 1606256979
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1606256979
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1606256979
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1606256979
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1606256979
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1606256979
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_8
timestamp 1606256979
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606256979
transform 1 0 1472 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606256979
transform 1 0 1472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1606256979
transform 1 0 2576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_16
timestamp 1606256979
transform 1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2852 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_20
timestamp 1606256979
transform 1 0 2944 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3036 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_28
timestamp 1606256979
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1606256979
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_37
timestamp 1606256979
transform 1 0 4508 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606256979
transform 1 0 6624 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4968 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_58
timestamp 1606256979
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1606256979
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_62
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7360 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7084 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_63
timestamp 1606256979
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1606256979
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1606256979
transform 1 0 9752 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9568 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10488 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1606256979
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1606256979
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_101
timestamp 1606256979
transform 1 0 10396 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_84
timestamp 1606256979
transform 1 0 8832 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12144 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1606256979
transform 1 0 11960 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_108
timestamp 1606256979
transform 1 0 11040 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1606256979
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13432 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13800 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1606256979
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1606256979
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_143
timestamp 1606256979
transform 1 0 14260 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15916 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15364 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_147
timestamp 1606256979
transform 1 0 14628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_160
timestamp 1606256979
transform 1 0 15824 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_164
timestamp 1606256979
transform 1 0 16192 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606256979
transform 1 0 16928 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16928 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1606256979
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1606256979
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606256979
transform 1 0 19044 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18584 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606256979
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1606256979
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_206
timestamp 1606256979
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_198
timestamp 1606256979
transform 1 0 19320 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606256979
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_210
timestamp 1606256979
transform 1 0 20424 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_218
timestamp 1606256979
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606256979
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606256979
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606256979
transform 1 0 2300 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1606256979
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1606256979
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606256979
transform 1 0 3404 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1606256979
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1606256979
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5336 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_44
timestamp 1606256979
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_62
timestamp 1606256979
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6992 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_70
timestamp 1606256979
transform 1 0 7544 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_78
timestamp 1606256979
transform 1 0 8280 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606256979
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1606256979
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_114
timestamp 1606256979
transform 1 0 11592 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606256979
transform 1 0 13064 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_126
timestamp 1606256979
transform 1 0 12696 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1606256979
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15548 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606256979
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_154
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1606256979
transform 1 0 17756 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_173
timestamp 1606256979
transform 1 0 17020 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1606256979
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1606256979
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606256979
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606256979
transform 1 0 1564 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2944 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1606256979
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_17
timestamp 1606256979
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_36
timestamp 1606256979
transform 1 0 4416 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1606256979
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5244 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_44
timestamp 1606256979
transform 1 0 5152 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1606256979
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7084 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_71
timestamp 1606256979
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10028 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_86
timestamp 1606256979
transform 1 0 9016 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_94
timestamp 1606256979
transform 1 0 9752 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1606256979
transform 1 0 11500 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1606256979
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_123
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 13156 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15180 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1606256979
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1606256979
transform 1 0 14628 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_162
timestamp 1606256979
transform 1 0 16008 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_174
timestamp 1606256979
transform 1 0 17112 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1606256979
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606256979
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1606256979
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1932 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1606256979
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1606256979
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_19
timestamp 1606256979
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606256979
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_41
timestamp 1606256979
transform 1 0 4876 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5428 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606256979
transform 1 0 7176 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8648 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7636 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_63
timestamp 1606256979
transform 1 0 6900 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_69
timestamp 1606256979
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1606256979
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10120 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1606256979
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1606256979
transform 1 0 10028 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12512 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11776 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1606256979
transform 1 0 11592 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_122
timestamp 1606256979
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_30_130
timestamp 1606256979
transform 1 0 13064 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1606256979
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16284 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1606256979
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18032 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17296 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_171
timestamp 1606256979
transform 1 0 16836 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_175
timestamp 1606256979
transform 1 0 17204 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1606256979
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18768 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1606256979
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_198
timestamp 1606256979
transform 1 0 19320 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1606256979
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606256979
transform 1 0 1656 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_10
timestamp 1606256979
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1606256979
transform 1 0 2760 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3220 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_22
timestamp 1606256979
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 1606256979
transform 1 0 4692 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5060 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606256979
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_62
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7728 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1606256979
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606256979
transform 1 0 9384 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10028 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_88
timestamp 1606256979
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1606256979
transform 1 0 9660 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606256979
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1606256979
transform 1 0 11500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606256979
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12788 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13616 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_133
timestamp 1606256979
transform 1 0 13340 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_142
timestamp 1606256979
transform 1 0 14168 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606256979
transform 1 0 15364 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14628 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15916 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_146
timestamp 1606256979
transform 1 0 14536 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_153
timestamp 1606256979
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_159
timestamp 1606256979
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16744 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_167
timestamp 1606256979
transform 1 0 16468 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_176
timestamp 1606256979
transform 1 0 17296 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1606256979
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606256979
transform 1 0 18768 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 19780 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_190
timestamp 1606256979
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_196
timestamp 1606256979
transform 1 0 19136 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_202
timestamp 1606256979
transform 1 0 19688 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606256979
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606256979
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606256979
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606256979
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1606256979
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1606256979
transform 1 0 2668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606256979
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_25
timestamp 1606256979
transform 1 0 3404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1606256979
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1606256979
transform 1 0 4876 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5244 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_54
timestamp 1606256979
transform 1 0 6072 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8648 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_75
timestamp 1606256979
transform 1 0 8004 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_81
timestamp 1606256979
transform 1 0 8556 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1606256979
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_103
timestamp 1606256979
transform 1 0 10580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606256979
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_115
timestamp 1606256979
transform 1 0 11684 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606256979
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606256979
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606256979
transform 1 0 12788 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13340 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_131
timestamp 1606256979
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1606256979
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1606256979
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606256979
transform 1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606256979
transform 1 0 14628 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_151
timestamp 1606256979
transform 1 0 14996 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1606256979
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_166
timestamp 1606256979
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606256979
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606256979
transform 1 0 17112 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606256979
transform 1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_172
timestamp 1606256979
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1606256979
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1606256979
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606256979
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1606256979
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1606256979
transform 1 0 19228 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_209
timestamp 1606256979
transform 1 0 20332 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal3 s 22320 11432 22800 11552 6 ccff_head
port 0 nsew default input
rlabel metal2 s 11426 0 11482 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 3790 22320 3846 22800 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 8390 22320 8446 22800 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 8850 22320 8906 22800 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 9310 22320 9366 22800 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 9770 22320 9826 22800 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10230 22320 10286 22800 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 10690 22320 10746 22800 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 12438 22320 12494 22800 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 4250 22320 4306 22800 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 5170 22320 5226 22800 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 5630 22320 5686 22800 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 6090 22320 6146 22800 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 6550 22320 6606 22800 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 7010 22320 7066 22800 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 7470 22320 7526 22800 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 7930 22320 7986 22800 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 12898 22320 12954 22800 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 17958 22320 18014 22800 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18418 22320 18474 22800 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 18878 22320 18934 22800 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19338 22320 19394 22800 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 19798 22320 19854 22800 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20258 22320 20314 22800 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 20718 22320 20774 22800 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 21178 22320 21234 22800 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 21638 22320 21694 22800 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 13358 22320 13414 22800 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 13818 22320 13874 22800 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 14278 22320 14334 22800 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 14738 22320 14794 22800 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 15198 22320 15254 22800 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 15658 22320 15714 22800 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 16118 22320 16174 22800 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 16578 22320 16634 22800 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 17038 22320 17094 22800 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_11_
port 82 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_13_
port 83 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_15_
port 84 nsew default input
rlabel metal3 s 0 3816 480 3936 6 left_bottom_grid_pin_17_
port 85 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 86 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 87 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_5_
port 88 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_7_
port 89 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_9_
port 90 nsew default input
rlabel metal2 s 22098 22320 22154 22800 6 prog_clk_0_N_in
port 91 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 92 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_43_
port 93 nsew default input
rlabel metal2 s 1030 22320 1086 22800 6 top_left_grid_pin_44_
port 94 nsew default input
rlabel metal2 s 1490 22320 1546 22800 6 top_left_grid_pin_45_
port 95 nsew default input
rlabel metal2 s 1950 22320 2006 22800 6 top_left_grid_pin_46_
port 96 nsew default input
rlabel metal2 s 2410 22320 2466 22800 6 top_left_grid_pin_47_
port 97 nsew default input
rlabel metal2 s 2870 22320 2926 22800 6 top_left_grid_pin_48_
port 98 nsew default input
rlabel metal2 s 3330 22320 3386 22800 6 top_left_grid_pin_49_
port 99 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 top_right_grid_pin_1_
port 100 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 101 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 102 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
