* NGSPICE file created from sb_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

.subckt sb_1__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_1_
+ left_top_grid_pin_42_ left_top_grid_pin_43_ left_top_grid_pin_44_ left_top_grid_pin_45_
+ left_top_grid_pin_46_ left_top_grid_pin_47_ left_top_grid_pin_48_ left_top_grid_pin_49_
+ prog_clk right_bottom_grid_pin_1_ right_top_grid_pin_42_ right_top_grid_pin_43_
+ right_top_grid_pin_44_ right_top_grid_pin_45_ right_top_grid_pin_46_ right_top_grid_pin_47_
+ right_top_grid_pin_48_ right_top_grid_pin_49_ top_left_grid_pin_34_ top_left_grid_pin_35_
+ top_left_grid_pin_36_ top_left_grid_pin_37_ top_left_grid_pin_38_ top_left_grid_pin_39_
+ top_left_grid_pin_40_ top_left_grid_pin_41_ VPWR VGND
XFILLER_39_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_3__A0 _060_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_38.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A1 mux_left_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_36.mux_l2_in_0__A0 _048_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__124__A _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_062_ _062_/HI _062_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__A1 left_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__119__A _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l3_in_0_ mux_top_track_10.mux_l2_in_1_/X mux_top_track_10.mux_l2_in_0_/X
+ mux_top_track_10.mux_l3_in_0_/S mux_top_track_10.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_28.mux_l2_in_0__A1 mux_top_track_28.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_3__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_114_ _114_/A chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l2_in_1__A1 mux_left_track_33.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l2_in_1_ _035_/HI chanx_left_in[9] mux_top_track_10.mux_l2_in_0_/S
+ mux_top_track_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l3_in_0__S mux_right_track_16.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 right_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_33.mux_l3_in_0__A1 mux_left_track_33.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_2__A0 left_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_2__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_36.mux_l2_in_0__A1 mux_top_track_36.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A mux_left_track_1.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l3_in_1__A0 mux_left_track_9.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ _061_/HI _061_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_30.mux_l2_in_0__S mux_top_track_30.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_2__S mux_left_track_1.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X _081_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ _113_/A chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l4_in_0__A0 mux_left_track_9.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_2__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_10.mux_l2_in_0_ chanx_right_in[19] mux_top_track_10.mux_l1_in_0_/X
+ mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_8.mux_l2_in_3_ _033_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_12.mux_l1_in_1_/S mux_top_track_12.mux_l2_in_0_/S
+ mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A mux_top_track_20.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _073_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_top_track_0.mux_l2_in_3_ _034_/HI chanx_left_in[2] mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_9.mux_l2_in_2__A1 left_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_1__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__S mux_right_track_32.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_10.mux_l2_in_0__A0 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_3__A0 right_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_37_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_1__A1 mux_left_track_9.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S mux_right_track_8.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ _060_/HI _060_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S mux_top_track_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_2__A0 mux_right_track_4.mux_l1_in_5_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ top_left_grid_pin_35_ chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_9.mux_l4_in_0__A1 mux_left_track_9.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_4.mux_l3_in_1__A0 mux_right_track_4.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_25.mux_l2_in_1__S mux_left_track_25.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_10.mux_l3_in_0_/S mux_top_track_12.mux_l1_in_1_/S
+ mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] right_bottom_grid_pin_1_ mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[0] chanx_right_in[2] mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l1_in_0_ chanx_right_in[9] top_left_grid_pin_35_ mux_top_track_10.mux_l1_in_0_/S
+ mux_top_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A0 mux_right_track_4.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_22.mux_l2_in_0_ mux_top_track_22.mux_l1_in_1_/X mux_top_track_22.mux_l1_in_0_/X
+ mux_top_track_22.mux_l2_in_0_/S mux_top_track_22.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0__A1 mux_top_track_10.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A mux_top_track_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 right_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_2__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_18.mux_l1_in_1_/S mux_top_track_18.mux_l2_in_0_/S
+ mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 mux_top_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_22.mux_l1_in_1_ _042_/HI chanx_left_in[17] mux_top_track_22.mux_l1_in_1_/S
+ mux_top_track_22.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_6.mux_l2_in_0__S mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_4.mux_l2_in_2__A1 mux_right_track_4.mux_l1_in_4_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_111_ _111_/A chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__072__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l3_in_1__A1 mux_right_track_4.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__A0 mux_top_track_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_20.mux_l1_in_0__S mux_top_track_20.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_2__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__067__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_1_ right_top_grid_pin_46_ right_top_grid_pin_42_ mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ chanx_right_in[1] top_left_grid_pin_40_ mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A1 mux_right_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_0.mux_l4_in_0__A0 mux_top_track_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X _114_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__080__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_16.mux_l2_in_0_/S mux_top_track_18.mux_l1_in_1_/S
+ mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_14.mux_l1_in_0__A0 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X _117_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_top_track_22.mux_l1_in_0_ chanx_right_in[17] top_left_grid_pin_41_ mux_top_track_22.mux_l1_in_1_/S
+ mux_top_track_22.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__075__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_1.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_34.mux_l2_in_0_ _047_/HI mux_top_track_34.mux_l1_in_0_/X mux_top_track_34.mux_l2_in_0_/S
+ mux_top_track_34.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_110_ _110_/A chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A mux_top_track_6.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_30.mux_l1_in_0_/S mux_top_track_30.mux_l2_in_0_/S
+ mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0__S mux_top_track_12.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l1_in_1__S mux_top_track_18.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__A1 mux_top_track_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X _125_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA__083__A _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_0_ chany_top_in[16] mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 right_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l2_in_0_ top_left_grid_pin_38_ mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_0.mux_l4_in_0__A1 mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__078__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_14.mux_l1_in_0__A1 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__091__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0__A0 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__086__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_38.sky130_fd_sc_hd__buf_4_0_ mux_top_track_38.mux_l2_in_0_/X _106_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_28.mux_l2_in_0_/S mux_top_track_30.mux_l1_in_0_/S
+ mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_34.mux_l1_in_0_ chanx_left_in[7] top_left_grid_pin_39_ mux_top_track_34.mux_l1_in_0_/S
+ mux_top_track_34.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l4_in_0_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_30.mux_l1_in_0__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 right_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 mux_top_track_4.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_36.mux_l1_in_0_/S mux_top_track_36.mux_l2_in_0_/S
+ mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 right_top_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__094__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_32.mux_l2_in_1_/S
+ mux_right_track_32.mux_l3_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_22.mux_l1_in_0__A1 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__S mux_top_track_38.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__089__A _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l4_in_0__S mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X _101_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 top_left_grid_pin_35_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ chanx_left_in[5] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l4_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 right_top_grid_pin_44_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A mux_top_track_12.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X _089_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l3_in_1_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_30.mux_l1_in_0__A1 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_6_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 mux_top_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_1__S mux_top_track_14.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 _038_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 left_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_34.mux_l2_in_0_/S mux_top_track_36.mux_l1_in_0_/S
+ mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_1_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_3__A0 _053_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 mux_top_track_16.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l2_in_3_ _056_/HI left_top_grid_pin_49_ mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l3_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ chanx_left_in[6] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 right_top_grid_pin_45_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l4_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S mux_left_track_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 _043_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_3.mux_l2_in_2_/S mux_left_track_3.mux_l3_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_0_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l1_in_5_ right_bottom_grid_pin_1_ right_top_grid_pin_49_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_5_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 mux_right_track_32.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 mux_top_track_24.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_3__A1 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l4_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A mux_top_track_18.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l3_in_0_/S
+ mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_3.mux_l2_in_2_ left_top_grid_pin_47_ left_top_grid_pin_45_ mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_6.mux_l1_in_3__A0 _051_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_34.mux_l1_in_0__S mux_top_track_34.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_3_ _065_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_1_/S
+ mux_right_track_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_097_ _097_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_2_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_32.mux_l2_in_0__A0 _046_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_top_track_0.mux_l1_in_0_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l1_in_4_ right_top_grid_pin_48_ right_top_grid_pin_47_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_4_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_5.mux_l1_in_5__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l3_in_1_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_6.mux_l1_in_3_/S mux_top_track_6.mux_l2_in_0_/S
+ mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_3.mux_l2_in_1_ left_top_grid_pin_43_ chanx_right_in[13] mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l2_in_3__S mux_left_track_9.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_3__A0 left_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_3__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A mux_left_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_22.mux_l1_in_1_/S mux_top_track_22.mux_l2_in_0_/S
+ mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA__100__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A mux_top_track_30.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_2__A0 mux_left_track_5.mux_l1_in_5_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_096_ chanx_left_in[8] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_1_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_1.mux_l4_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_3__S mux_right_track_24.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A1 mux_top_track_32.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ chanx_right_in[5] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_3_ _061_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_3_ right_top_grid_pin_46_ right_top_grid_pin_45_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_1__A0 mux_left_track_5.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l1_in_1_ _038_/HI chanx_left_in[13] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l4_in_0__A0 mux_left_track_5.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_28.mux_l1_in_0__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_4.mux_l3_in_0_/S mux_top_track_6.mux_l1_in_3_/S
+ mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_3.mux_l2_in_0_ chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/X mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 left_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_20.mux_l2_in_0_/S mux_top_track_22.mux_l1_in_1_/S
+ mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_3__S mux_left_track_17.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_2__A1 mux_left_track_5.mux_l1_in_4_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_095_ chanx_left_in[9] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_38.mux_l2_in_0_/S mux_right_track_0.mux_l1_in_1_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_30.mux_l1_in_0__S mux_top_track_30.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A0 mux_left_track_33.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2__S mux_left_track_1.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ chanx_right_in[6] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X _119_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] right_top_grid_pin_47_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_28.mux_l1_in_0_/S mux_top_track_28.mux_l2_in_0_/S
+ mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_right_track_4.mux_l1_in_2_ right_top_grid_pin_44_ right_top_grid_pin_43_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_1__A1 mux_left_track_5.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A mux_top_track_36.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_38_ mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_24.mux_l2_in_1_/S
+ mux_right_track_24.mux_l3_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_36.mux_l1_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_28.mux_l2_in_0_ _044_/HI mux_top_track_28.mux_l1_in_0_/X mux_top_track_28.mux_l2_in_0_/S
+ mux_top_track_28.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l3_in_0__S mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_30.mux_l2_in_0_ _045_/HI mux_top_track_30.mux_l1_in_0_/X mux_top_track_30.mux_l2_in_0_/S
+ mux_top_track_30.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_5.mux_l4_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_5.mux_l4_in_0__A1 mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_3_ _051_/HI chanx_left_in[6] mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_28.mux_l1_in_0__A1 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__114__A _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_1__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l3_in_1__A0 mux_right_track_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_33.mux_l2_in_0_/S ccff_tail
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_5__S mux_right_track_4.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l2_in_0__S mux_top_track_22.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_3__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l4_in_0__S mux_left_track_3.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l2_in_3__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S mux_top_track_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l4_in_0__A0 mux_right_track_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_094_ chanx_left_in[10] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_9.mux_l3_in_1__S mux_left_track_9.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A1 mux_left_track_33.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__122__A _122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_077_ _077_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l1_in_1_ right_top_grid_pin_43_ chany_top_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_24.mux_l2_in_0_/S mux_top_track_28.mux_l1_in_0_/S
+ mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_1_ right_top_grid_pin_42_ chany_top_in[15] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_1_ mux_top_track_6.mux_l1_in_3_/X mux_top_track_6.mux_l1_in_2_/X
+ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l2_in_1_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_36.mux_l1_in_0__A1 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_34.sky130_fd_sc_hd__buf_4_0_ mux_top_track_34.mux_l2_in_0_/X _108_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A1 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_6__A0 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_2_ chanx_right_in[11] chanx_right_in[6] mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_28.mux_l1_in_0_ chanx_left_in[19] top_left_grid_pin_36_ mux_top_track_28.mux_l1_in_0_/S
+ mux_top_track_28.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_28.sky130_fd_sc_hd__buf_4_0_ mux_top_track_28.mux_l2_in_0_/X _111_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_10.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_1__A1 mux_right_track_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_0_/S
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_top_track_30.mux_l1_in_0_ chanx_left_in[15] top_left_grid_pin_37_ mux_top_track_30.mux_l1_in_0_/S
+ mux_top_track_30.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__125__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ _093_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l4_in_0__A1 mux_right_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_076_ chanx_right_in[8] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X _103_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_16.mux_l3_in_0_/S
+ mux_right_track_24.mux_l1_in_1_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ _059_/HI _059_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X _122_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__S mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_6__A1 left_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_1_ top_left_grid_pin_41_ top_left_grid_pin_39_ mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_3__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 mux_right_track_4.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_092_ chanx_left_in[12] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_38.mux_l1_in_1__A0 _049_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A mux_left_track_3.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A0 _062_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_3__S mux_left_track_1.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_075_ chanx_right_in[9] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_24.mux_l1_in_1__S mux_top_track_24.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l4_in_0__S mux_right_track_2.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_12.mux_l1_in_0__S mux_top_track_12.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l3_in_1__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _097_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 top_left_grid_pin_35_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l3_in_1__S mux_right_track_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l2_in_0__A0 mux_top_track_38.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_058_ _058_/HI _058_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A mux_left_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_14.mux_l1_in_0_/S mux_top_track_14.mux_l2_in_0_/S
+ mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A mux_top_track_22.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X _085_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_10.mux_l3_in_0__S mux_top_track_10.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_091_ chanx_left_in[13] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_38.mux_l1_in_1__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_074_ chanx_right_in[10] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_38.mux_l2_in_0__A1 mux_top_track_38.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_057_ _057_/HI _057_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_35_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A mux_left_track_9.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_109_ _109_/A chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_3_ _059_/HI left_bottom_grid_pin_1_ mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__070__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_3_ _060_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_12.mux_l2_in_0_/S mux_top_track_14.mux_l1_in_0_/S
+ mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_3__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_1__A0 _036_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_6.mux_l2_in_1__S mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_090_ chanx_left_in[14] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A mux_top_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S mux_left_track_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S mux_right_track_0.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_073_ _073_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_28.sky130_fd_sc_hd__buf_4_0__A mux_top_track_28.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_12.mux_l2_in_0__A0 mux_top_track_12.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_16.mux_l2_in_1_/S
+ mux_right_track_16.mux_l3_in_0_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__073__A _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_125_ _125_/A chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_056_ _056_/HI _056_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_20.mux_l1_in_1__S mux_top_track_20.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_3__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__068__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_1.mux_l3_in_1__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_36.mux_l2_in_0__S mux_top_track_36.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_3_ _054_/HI left_top_grid_pin_47_ mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l2_in_2_ left_top_grid_pin_46_ left_top_grid_pin_42_ mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l3_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] right_bottom_grid_pin_1_ mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_20.mux_l1_in_1__A0 _041_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_12.mux_l2_in_0_ mux_top_track_12.mux_l1_in_1_/X mux_top_track_12.mux_l1_in_0_/X
+ mux_top_track_12.mux_l2_in_0_/S mux_top_track_12.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__081__A _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _069_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__076__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_20.mux_l2_in_0__A0 mux_top_track_20.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_12.mux_l1_in_1_ _036_/HI chanx_left_in[10] mux_top_track_12.mux_l1_in_1_/S
+ mux_top_track_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l3_in_0__S mux_right_track_32.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_072_ chanx_right_in[12] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_12.mux_l2_in_0__A1 mux_top_track_12.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l2_in_1_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_3__A0 _040_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_124_ _124_/A chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 mux_top_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A mux_top_track_8.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_32.mux_l1_in_0_/S mux_top_track_32.mux_l2_in_0_/S
+ mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__084__A _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A1 right_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_2_ left_top_grid_pin_43_ chanx_right_in[17] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_1_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__079__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_1_ right_top_grid_pin_48_ right_top_grid_pin_46_ mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_20.mux_l1_in_1__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__S mux_left_track_25.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__092__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_20.mux_l2_in_0__A1 mux_top_track_20.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_12.mux_l1_in_0_ chanx_right_in[10] top_left_grid_pin_36_ mux_top_track_12.mux_l1_in_1_/S
+ mux_top_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__087__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_071_ chanx_right_in[13] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_8.mux_l4_in_0_/S mux_right_track_16.mux_l1_in_3_/S
+ mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_3_ _040_/HI chanx_left_in[4] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_24.mux_l1_in_3_ _063_/HI chanx_left_in[18] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_3__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ _123_/A chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_1_ _043_/HI chanx_left_in[18] mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_30.mux_l2_in_0_/S mux_top_track_32.mux_l1_in_0_/S
+ mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l1_in_1_ chanx_right_in[8] chany_top_in[17] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_106_ _106_/A chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_0_ chany_top_in[18] mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_2__A0 left_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A mux_right_track_16.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__095__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_32.mux_l2_in_0__S mux_top_track_32.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l3_in_1__S mux_right_track_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_2__S mux_left_track_3.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_38.mux_l1_in_1__S mux_top_track_38.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_38.mux_l1_in_1_/S mux_top_track_38.mux_l2_in_0_/S
+ mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_1.mux_l3_in_1__A0 mux_left_track_1.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_30.sky130_fd_sc_hd__buf_4_0_ mux_top_track_30.mux_l2_in_0_/X _110_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_right_track_0.mux_l1_in_1_ right_top_grid_pin_44_ right_top_grid_pin_42_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l4_in_0__A0 mux_left_track_1.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_070_ chanx_right_in[14] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X _113_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l2_in_3__A0 _033_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_2_ chanx_right_in[4] chanx_right_in[3] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[9] right_top_grid_pin_48_ mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__098__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_122_ _122_/A chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[18] top_left_grid_pin_34_ mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_36.mux_l2_in_0_ _048_/HI mux_top_track_36.mux_l1_in_0_/X mux_top_track_36.mux_l2_in_0_/S
+ mux_top_track_36.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X _116_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A mux_right_track_2.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_105_ _105_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_1.mux_l2_in_2__A1 left_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A mux_left_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l4_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l2_in_0__S mux_top_track_18.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A mux_top_track_14.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l3_in_0_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_6.mux_l1_in_2__A0 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X _105_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_36.mux_l2_in_0_/S mux_top_track_38.mux_l1_in_1_/S
+ mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.mux_l3_in_1__A1 mux_left_track_1.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _124_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_6.mux_l2_in_1__A0 mux_top_track_6.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l4_in_0__A1 mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_3__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_41_ top_left_grid_pin_39_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_1_ right_top_grid_pin_44_ chany_top_in[18] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A0 mux_top_track_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A0 _061_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_121_ _121_/A chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l4_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_104_ _104_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_6_ left_bottom_grid_pin_1_ left_top_grid_pin_49_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l3_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_0_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_36.mux_l1_in_0_ chanx_left_in[3] top_left_grid_pin_40_ mux_top_track_36.mux_l1_in_0_/S
+ mux_top_track_36.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l2_in_1__A1 mux_top_track_6.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_1__A0 _039_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 mux_left_track_5.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_22.mux_l1_in_0__S mux_top_track_22.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l3_in_0_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_2.mux_l2_in_2__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_25.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A0 _063_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_3__A0 _056_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_18.mux_l2_in_0__A0 mux_top_track_18.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A1 mux_top_track_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A1 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_120_ _120_/A chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_103_ _103_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l3_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_5_ left_top_grid_pin_48_ left_top_grid_pin_47_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_5_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_5.mux_l1_in_0_/S mux_left_track_5.mux_l2_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_0.mux_l4_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_6__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l4_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0__S mux_top_track_14.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_1__A1 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__101__A _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_1_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_24.mux_l1_in_3__A1 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_3.mux_l2_in_3__A1 left_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_3_ _058_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_0_/S
+ mux_left_track_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_18.mux_l2_in_0__A1 mux_top_track_18.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_24.mux_l1_in_1_/S mux_top_track_24.mux_l2_in_0_/S
+ mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A mux_top_track_32.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_1_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 right_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_033_ _033_/HI _033_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_102_ chanx_left_in[2] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_17.mux_l1_in_1_/S mux_left_track_17.mux_l2_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_4_ left_top_grid_pin_46_ left_top_grid_pin_45_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_4_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_3.mux_l4_in_0_/S mux_left_track_5.mux_l1_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__104__A _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_1_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_34.mux_l2_in_0__A0 _047_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_6.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_17.mux_l1_in_3__A0 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__112__A top_left_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_2_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_22.mux_l2_in_0_/S mux_top_track_24.mux_l1_in_1_/S
+ mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__S mux_right_track_4.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_0.mux_l4_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 right_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_101_ _101_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_9.mux_l4_in_0_/S mux_left_track_17.mux_l1_in_1_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_5.mux_l1_in_3_ left_top_grid_pin_44_ left_top_grid_pin_43_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_5__A0 left_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__120__A _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A mux_top_track_38.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _077_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_34.mux_l2_in_0__A1 mux_top_track_34.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_2__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_3__A0 _055_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_6__S mux_right_track_4.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0__S mux_top_track_10.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_17.mux_l1_in_3__A1 left_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__123__A _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_100_ chanx_left_in[4] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__118__A _118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_42_ chanx_right_in[14] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D mux_top_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_3_ _055_/HI left_top_grid_pin_48_ mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l1_in_5__A1 left_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_2__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_18.mux_l2_in_0_ mux_top_track_18.mux_l1_in_1_/X mux_top_track_18.mux_l1_in_0_/X
+ mux_top_track_18.mux_l2_in_0_/S mux_top_track_18.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_20.mux_l2_in_0_ mux_top_track_20.mux_l1_in_1_/X mux_top_track_20.mux_l1_in_0_/X
+ mux_top_track_20.mux_l2_in_0_/S mux_top_track_20.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l3_in_0_/S
+ mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_4.mux_l4_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_12.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_3__A1 left_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_18.mux_l1_in_1_ _039_/HI chanx_left_in[14] mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_20.mux_l1_in_1_ _041_/HI chanx_left_in[16] mux_top_track_20.mux_l1_in_1_/S
+ mux_top_track_20.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_1__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l3_in_1__A0 mux_right_track_2.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_1_ chanx_right_in[5] chany_top_in[19] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_2_ left_top_grid_pin_44_ chanx_right_in[18] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X _115_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_36.mux_l1_in_0__S mux_top_track_36.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A0 mux_right_track_2.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__S mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_10.mux_l1_in_0_/S mux_top_track_10.mux_l2_in_0_/S
+ mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X _118_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_18.mux_l1_in_0_ chanx_right_in[14] top_left_grid_pin_39_ mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_20.mux_l1_in_0_ chanx_right_in[16] top_left_grid_pin_40_ mux_top_track_20.mux_l1_in_1_/S
+ mux_top_track_20.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_38.mux_l1_in_0__A1 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l2_in_0_ _046_/HI mux_top_track_32.mux_l1_in_0_/X mux_top_track_32.mux_l2_in_0_/S
+ mux_top_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_2__A1 right_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l2_in_3__A0 _059_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_2.mux_l3_in_1__A1 mux_right_track_2.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_1__S mux_top_track_12.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_28.mux_l2_in_0__S mux_top_track_28.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A mux_left_track_5.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l4_in_0__S mux_left_track_9.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_1_ chanx_right_in[9] chany_top_in[16] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_089_ _089_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A1 mux_right_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S mux_right_track_32.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_8.mux_l3_in_0_/S mux_top_track_10.mux_l1_in_0_/S
+ mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l2_in_1_ _052_/HI chanx_left_in[8] mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__A0 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_1_ _064_/HI mux_right_track_32.mux_l1_in_2_/X mux_right_track_32.mux_l2_in_1_/S
+ mux_right_track_32.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_36.sky130_fd_sc_hd__buf_4_0_ mux_top_track_36.mux_l2_in_0_/X _107_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_41_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_16.mux_l1_in_1_/S mux_top_track_16.mux_l2_in_0_/S
+ mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A mux_top_track_24.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_32.mux_l1_in_2_ chanx_left_in[10] right_top_grid_pin_49_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_3__A1 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l1_in_0_ chanx_left_in[11] top_left_grid_pin_38_ mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_10.mux_l2_in_1__A0 _035_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_4__A0 right_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_088_ chanx_left_in[16] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l3_in_0__A0 mux_top_track_10.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A0 _065_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__071__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l3_in_0__S mux_left_track_17.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__S mux_top_track_32.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_0_ chanx_right_in[15] mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__A1 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__066__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_1_/S mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__S mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_14.mux_l2_in_0_/S mux_top_track_16.mux_l1_in_1_/S
+ mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X _121_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l1_in_1_ right_top_grid_pin_45_ chany_top_in[19] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A mux_top_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_10.mux_l2_in_1__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__074__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_4__A1 right_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ chanx_left_in[17] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 mux_top_track_2.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__069__A _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l3_in_0__A1 mux_top_track_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _093_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_20.mux_l1_in_0__A1 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l4_in_0__S mux_left_track_5.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_3__A1 mux_right_track_4.mux_l1_in_6_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__A0 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l4_in_0__S mux_right_track_8.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l1_in_0__S mux_top_track_18.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_3_ _053_/HI left_bottom_grid_pin_1_ mux_left_track_1.mux_l2_in_2_/S
+ mux_left_track_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__082__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__077__A _077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[8] top_left_grid_pin_34_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_32.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_2__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 left_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S mux_left_track_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__090__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_086_ chanx_left_in[18] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 mux_top_track_2.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 left_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_14.mux_l1_in_1__A0 _037_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X _084_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_17_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ _069_/A chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_34.mux_l1_in_0_/S mux_top_track_34.mux_l2_in_0_/S
+ mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_14.mux_l2_in_0__A0 mux_top_track_14.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l2_in_2_ left_top_grid_pin_48_ left_top_grid_pin_46_ mux_left_track_1.mux_l2_in_2_/S
+ mux_left_track_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__093__A _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_3_ _062_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__088__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_22.mux_l1_in_1__A0 _042_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l3_in_1__A0 mux_right_track_8.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__S mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_085_ _085_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 mux_left_track_1.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_1__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l4_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_22.mux_l2_in_0__A0 mux_top_track_22.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S mux_right_track_2.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A mux_top_track_10.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_068_ chanx_right_in[16] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_6.mux_l1_in_1__A0 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l4_in_0__A0 mux_right_track_8.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__096__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_32.mux_l2_in_0_/S mux_top_track_34.mux_l1_in_0_/S
+ mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_14.mux_l2_in_0__A1 mux_top_track_14.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_20.mux_l2_in_0__S mux_top_track_20.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ left_top_grid_pin_44_ mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_2_/S mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_3__S mux_left_track_3.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_3__A0 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l4_in_0__S mux_left_track_1.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_6.mux_l2_in_0__A0 mux_top_track_6.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__S mux_right_track_4.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__S mux_top_track_14.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A1 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_2_ left_top_grid_pin_42_ chanx_right_in[12] mux_left_track_1.mux_l1_in_2_/S
+ mux_left_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] right_top_grid_pin_49_ mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_14.mux_l2_in_0_ mux_top_track_14.mux_l1_in_1_/X mux_top_track_14.mux_l1_in_0_/X
+ mux_top_track_14.mux_l2_in_0_/S mux_top_track_14.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_22.mux_l1_in_1__A1 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_30.mux_l2_in_0__A0 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l3_in_1__A1 mux_right_track_8.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__099__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_084_ _084_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 mux_right_track_16.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_1.mux_l2_in_2_/S mux_left_track_1.mux_l3_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_top_track_14.mux_l1_in_1_ _037_/HI chanx_left_in[12] mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_22.mux_l2_in_0__A1 mux_top_track_22.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ chanx_right_in[17] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l4_in_0__A1 mux_right_track_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_1__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l3_in_0__A0 mux_right_track_16.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_119_ _119_/A chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_2_/S mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_3__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0__A1 mux_top_track_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A mux_top_track_16.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l3_in_0_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_1_ chanx_right_in[2] chany_top_in[14] mux_left_track_1.mux_l1_in_2_/S
+ mux_left_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_2__A0 left_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ right_top_grid_pin_47_ right_top_grid_pin_45_ mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A1 right_top_grid_pin_47_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 mux_right_track_24.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l3_in_0_/X _120_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_30.mux_l2_in_0__A1 mux_top_track_30.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_3.mux_l3_in_1__A0 mux_left_track_3.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_083_ _083_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A1 mux_right_track_16.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_14.mux_l1_in_0_ chanx_right_in[12] top_left_grid_pin_37_ mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_1.mux_l1_in_2_/S mux_left_track_1.mux_l2_in_2_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_3__S mux_top_track_4.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_066_ chanx_right_in[18] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_3.mux_l4_in_0__A0 mux_left_track_3.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A1 mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_3_ _050_/HI chanx_left_in[5] mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l4_in_0_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_118_ _118_/A chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_32.mux_l1_in_2__A0 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_4.mux_l1_in_1_/S mux_top_track_4.mux_l2_in_1_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_24.mux_l1_in_2__A1 right_top_grid_pin_48_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l2_in_1__A0 _064_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_left_track_1.mux_l1_in_2_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_2__A1 left_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_1__S mux_top_track_22.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_4__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0__S mux_top_track_10.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l4_in_0__S mux_right_track_0.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l3_in_1__S mux_left_track_3.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ _057_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_0_/S
+ mux_left_track_33.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_38.mux_l2_in_0__S mux_top_track_38.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_20.mux_l1_in_1_/S mux_top_track_20.mux_l2_in_0_/S
+ mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 mux_right_track_24.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_2__S mux_left_track_9.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l3_in_0__A0 mux_right_track_32.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_3.mux_l3_in_1__A1 mux_left_track_3.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ chanx_right_in[2] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l1_in_1_ right_top_grid_pin_43_ chany_top_in[14] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_2_ left_top_grid_pin_49_ left_top_grid_pin_45_ mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_34.mux_l1_in_0__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l2_in_0_/X _109_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_32.mux_l3_in_0_/S mux_left_track_1.mux_l1_in_2_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 _052_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ _065_/HI _065_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l4_in_0__A1 mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_2_ chanx_right_in[7] chanx_right_in[5] mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ _117_/A chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l1_in_2__S mux_right_track_24.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_32.mux_l1_in_2__A1 right_top_grid_pin_49_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l3_in_0__A0 mux_top_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_38.mux_l2_in_0_ mux_top_track_38.mux_l1_in_1_/X mux_top_track_38.mux_l1_in_0_/X
+ mux_top_track_38.mux_l2_in_0_/S mux_top_track_38.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_1_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2__A0 left_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__A1 mux_right_track_32.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__102__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_0_/S mux_left_track_33.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_38.mux_l1_in_1_ _049_/HI chanx_left_in[1] mux_top_track_38.mux_l1_in_1_/S
+ mux_top_track_38.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_18.mux_l2_in_0_/S mux_top_track_20.mux_l1_in_1_/S
+ mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 mux_left_track_17.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l3_in_0__A1 mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X _104_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_081_ _081_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_33.mux_l1_in_1_ chanx_right_in[10] chany_top_in[15] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_4__A0 left_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_34.mux_l1_in_0__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _123_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_left_track_17.mux_l1_in_2__S mux_left_track_17.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A0 mux_left_track_17.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_064_ _064_/HI _064_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__110__A _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A mux_top_track_34.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_40_ top_left_grid_pin_38_ mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_4.mux_l1_in_3_/S mux_right_track_4.mux_l2_in_1_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ _116_/A chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_3__A0 _058_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_25.mux_l1_in_2__A0 left_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A1 mux_top_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l2_in_1__A0 mux_left_track_25.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_38.mux_l1_in_0_ chanx_right_in[0] top_left_grid_pin_41_ mux_top_track_38.mux_l1_in_1_/S
+ mux_top_track_38.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A1 mux_left_track_17.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A0 mux_left_track_25.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ chanx_right_in[4] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_34.mux_l2_in_0__S mux_top_track_34.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_4__S mux_right_track_4.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_33.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__108__A _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l3_in_1__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_2__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_4__A1 left_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_2__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_17.mux_l3_in_0__A1 mux_left_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_28.mux_l1_in_0__S mux_top_track_28.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ _063_/HI _063_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__A0 left_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_28.mux_l2_in_0__A0 _044_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_2.mux_l4_in_0_/S mux_right_track_4.mux_l1_in_3_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_115_ _115_/A chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_5.mux_l2_in_3__A1 mux_left_track_5.mux_l1_in_6_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA__121__A _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__A0 _057_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__116__A _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 right_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_25.mux_l2_in_1__A1 mux_left_track_25.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A0 mux_left_track_33.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l2_in_1__S mux_top_track_10.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

