magic
tech EFS8A
magscale 1 2
timestamp 1604399647
<< locali >>
rect 8493 4063 8527 4233
rect 3709 2431 3743 2533
<< viali >>
rect 1593 24361 1627 24395
rect 1409 24225 1443 24259
rect 1593 23817 1627 23851
rect 2697 23817 2731 23851
rect 1409 23613 1443 23647
rect 2513 23613 2547 23647
rect 3157 23545 3191 23579
rect 2053 23477 2087 23511
rect 2421 23477 2455 23511
rect 1593 23273 1627 23307
rect 1409 23137 1443 23171
rect 1593 22729 1627 22763
rect 2053 22593 2087 22627
rect 1409 22525 1443 22559
rect 2421 22389 2455 22423
rect 1409 22049 1443 22083
rect 1593 21913 1627 21947
rect 1685 21301 1719 21335
rect 1593 21097 1627 21131
rect 1409 20961 1443 20995
rect 1685 20349 1719 20383
rect 1593 20009 1627 20043
rect 1409 19873 1443 19907
rect 8125 19261 8159 19295
rect 1685 19125 1719 19159
rect 8309 19125 8343 19159
rect 8769 19125 8803 19159
rect 1593 18377 1627 18411
rect 7757 18377 7791 18411
rect 1409 18173 1443 18207
rect 7573 18173 7607 18207
rect 2053 18037 2087 18071
rect 8217 18037 8251 18071
rect 1593 17833 1627 17867
rect 1409 17697 1443 17731
rect 2697 17221 2731 17255
rect 1409 17085 1443 17119
rect 2513 17085 2547 17119
rect 3065 17085 3099 17119
rect 1593 16949 1627 16983
rect 2053 16949 2087 16983
rect 1593 16745 1627 16779
rect 5733 16745 5767 16779
rect 7481 16745 7515 16779
rect 6101 16609 6135 16643
rect 6193 16609 6227 16643
rect 7297 16609 7331 16643
rect 6377 16541 6411 16575
rect 5457 16201 5491 16235
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 6837 16065 6871 16099
rect 5273 15997 5307 16031
rect 5917 15929 5951 15963
rect 5181 15861 5215 15895
rect 7297 15861 7331 15895
rect 1593 15657 1627 15691
rect 6009 15657 6043 15691
rect 6377 15589 6411 15623
rect 1409 15521 1443 15555
rect 6469 15453 6503 15487
rect 6561 15453 6595 15487
rect 4353 15317 4387 15351
rect 7021 15317 7055 15351
rect 5733 15113 5767 15147
rect 8217 15113 8251 15147
rect 1685 15045 1719 15079
rect 2605 15045 2639 15079
rect 2973 15045 3007 15079
rect 4169 15045 4203 15079
rect 6377 15045 6411 15079
rect 3709 14977 3743 15011
rect 4721 14977 4755 15011
rect 6837 14977 6871 15011
rect 2421 14909 2455 14943
rect 4077 14841 4111 14875
rect 4537 14841 4571 14875
rect 7082 14841 7116 14875
rect 4629 14773 4663 14807
rect 6101 14773 6135 14807
rect 1593 14569 1627 14603
rect 4261 14569 4295 14603
rect 6837 14569 6871 14603
rect 7389 14569 7423 14603
rect 5702 14501 5736 14535
rect 1409 14433 1443 14467
rect 5457 14433 5491 14467
rect 1593 14025 1627 14059
rect 6837 14025 6871 14059
rect 5641 13957 5675 13991
rect 6285 13957 6319 13991
rect 2053 13889 2087 13923
rect 4169 13889 4203 13923
rect 7389 13889 7423 13923
rect 1409 13821 1443 13855
rect 2329 13821 2363 13855
rect 3801 13821 3835 13855
rect 4261 13821 4295 13855
rect 4506 13753 4540 13787
rect 7297 13753 7331 13787
rect 6561 13685 6595 13719
rect 7205 13685 7239 13719
rect 1593 13481 1627 13515
rect 2697 13481 2731 13515
rect 5457 13481 5491 13515
rect 7205 13481 7239 13515
rect 6009 13413 6043 13447
rect 6929 13413 6963 13447
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 4344 13345 4378 13379
rect 4077 13277 4111 13311
rect 2329 13141 2363 13175
rect 3893 13141 3927 13175
rect 3341 12937 3375 12971
rect 4813 12937 4847 12971
rect 3801 12869 3835 12903
rect 2697 12801 2731 12835
rect 2881 12801 2915 12835
rect 4353 12801 4387 12835
rect 4169 12733 4203 12767
rect 2145 12665 2179 12699
rect 2605 12665 2639 12699
rect 1685 12597 1719 12631
rect 2237 12597 2271 12631
rect 3709 12597 3743 12631
rect 4261 12597 4295 12631
rect 1593 12393 1627 12427
rect 2329 12393 2363 12427
rect 2973 12393 3007 12427
rect 5457 12393 5491 12427
rect 2605 12325 2639 12359
rect 4344 12325 4378 12359
rect 1409 12257 1443 12291
rect 4077 12257 4111 12291
rect 12256 12257 12290 12291
rect 11989 12189 12023 12223
rect 3893 12053 3927 12087
rect 13369 12053 13403 12087
rect 1593 11849 1627 11883
rect 2145 11849 2179 11883
rect 3709 11849 3743 11883
rect 12081 11849 12115 11883
rect 3801 11713 3835 11747
rect 1961 11645 1995 11679
rect 3341 11577 3375 11611
rect 4068 11577 4102 11611
rect 2513 11509 2547 11543
rect 5181 11509 5215 11543
rect 12725 11509 12759 11543
rect 3801 11305 3835 11339
rect 4353 11305 4387 11339
rect 4445 11169 4479 11203
rect 4712 11169 4746 11203
rect 2973 11101 3007 11135
rect 5825 11033 5859 11067
rect 3617 10761 3651 10795
rect 4813 10761 4847 10795
rect 3801 10693 3835 10727
rect 4445 10625 4479 10659
rect 4169 10557 4203 10591
rect 2421 10421 2455 10455
rect 3341 10421 3375 10455
rect 4261 10421 4295 10455
rect 5273 10421 5307 10455
rect 8861 10421 8895 10455
rect 2421 10217 2455 10251
rect 3893 10217 3927 10251
rect 6101 10217 6135 10251
rect 7757 10217 7791 10251
rect 6193 10149 6227 10183
rect 2789 10081 2823 10115
rect 7849 10081 7883 10115
rect 11233 10081 11267 10115
rect 17224 10081 17258 10115
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 6377 10013 6411 10047
rect 7941 10013 7975 10047
rect 9689 10013 9723 10047
rect 10977 10013 11011 10047
rect 13829 10013 13863 10047
rect 16957 10013 16991 10047
rect 5733 9945 5767 9979
rect 7297 9945 7331 9979
rect 18337 9945 18371 9979
rect 1685 9877 1719 9911
rect 1961 9877 1995 9911
rect 5089 9877 5123 9911
rect 6929 9877 6963 9911
rect 7389 9877 7423 9911
rect 12357 9877 12391 9911
rect 13369 9877 13403 9911
rect 3065 9673 3099 9707
rect 4077 9673 4111 9707
rect 4997 9673 5031 9707
rect 11069 9673 11103 9707
rect 17325 9673 17359 9707
rect 4537 9605 4571 9639
rect 8769 9605 8803 9639
rect 3617 9537 3651 9571
rect 4905 9537 4939 9571
rect 5457 9537 5491 9571
rect 5641 9537 5675 9571
rect 13277 9537 13311 9571
rect 5365 9469 5399 9503
rect 6837 9469 6871 9503
rect 9597 9469 9631 9503
rect 9689 9469 9723 9503
rect 3525 9401 3559 9435
rect 7082 9401 7116 9435
rect 9229 9401 9263 9435
rect 9934 9401 9968 9435
rect 13544 9401 13578 9435
rect 1685 9333 1719 9367
rect 2053 9333 2087 9367
rect 2513 9333 2547 9367
rect 2973 9333 3007 9367
rect 3433 9333 3467 9367
rect 6101 9333 6135 9367
rect 6653 9333 6687 9367
rect 8217 9333 8251 9367
rect 11713 9333 11747 9367
rect 13185 9333 13219 9367
rect 14657 9333 14691 9367
rect 17049 9333 17083 9367
rect 1593 9129 1627 9163
rect 1961 9129 1995 9163
rect 3157 9129 3191 9163
rect 6101 9129 6135 9163
rect 9413 9129 9447 9163
rect 10057 9129 10091 9163
rect 11069 9129 11103 9163
rect 11437 9129 11471 9163
rect 14289 9129 14323 9163
rect 15669 9129 15703 9163
rect 7380 9061 7414 9095
rect 10701 9061 10735 9095
rect 12440 9061 12474 9095
rect 2053 8993 2087 9027
rect 4344 8993 4378 9027
rect 6929 8993 6963 9027
rect 7113 8993 7147 9027
rect 10149 8993 10183 9027
rect 15761 8993 15795 9027
rect 22201 8993 22235 9027
rect 2145 8925 2179 8959
rect 3433 8925 3467 8959
rect 4077 8925 4111 8959
rect 10241 8925 10275 8959
rect 12173 8925 12207 8959
rect 15853 8925 15887 8959
rect 8493 8857 8527 8891
rect 9689 8857 9723 8891
rect 2605 8789 2639 8823
rect 3893 8789 3927 8823
rect 5457 8789 5491 8823
rect 6469 8789 6503 8823
rect 13553 8789 13587 8823
rect 15301 8789 15335 8823
rect 22385 8789 22419 8823
rect 7665 8585 7699 8619
rect 10149 8585 10183 8619
rect 13461 8585 13495 8619
rect 16497 8585 16531 8619
rect 22477 8585 22511 8619
rect 1409 8517 1443 8551
rect 9597 8517 9631 8551
rect 10701 8517 10735 8551
rect 17049 8517 17083 8551
rect 21833 8517 21867 8551
rect 1869 8449 1903 8483
rect 1961 8449 1995 8483
rect 11253 8449 11287 8483
rect 12265 8449 12299 8483
rect 12909 8449 12943 8483
rect 13001 8449 13035 8483
rect 1777 8381 1811 8415
rect 2789 8381 2823 8415
rect 3525 8381 3559 8415
rect 3893 8381 3927 8415
rect 3985 8381 4019 8415
rect 4252 8381 4286 8415
rect 8217 8381 8251 8415
rect 10609 8381 10643 8415
rect 11161 8381 11195 8415
rect 14197 8381 14231 8415
rect 14453 8381 14487 8415
rect 16865 8381 16899 8415
rect 17325 8381 17359 8415
rect 21649 8381 21683 8415
rect 22109 8381 22143 8415
rect 2421 8313 2455 8347
rect 6837 8313 6871 8347
rect 8462 8313 8496 8347
rect 11069 8313 11103 8347
rect 11897 8313 11931 8347
rect 12817 8313 12851 8347
rect 16129 8313 16163 8347
rect 5365 8245 5399 8279
rect 7389 8245 7423 8279
rect 8125 8245 8159 8279
rect 12449 8245 12483 8279
rect 14105 8245 14139 8279
rect 15577 8245 15611 8279
rect 1409 8041 1443 8075
rect 3617 8041 3651 8075
rect 6469 8041 6503 8075
rect 7941 8041 7975 8075
rect 8585 8041 8619 8075
rect 9505 8041 9539 8075
rect 12173 8041 12207 8075
rect 12633 8041 12667 8075
rect 13001 8041 13035 8075
rect 14013 8041 14047 8075
rect 15669 8041 15703 8075
rect 17233 8041 17267 8075
rect 9956 7973 9990 8007
rect 15117 7973 15151 8007
rect 1777 7905 1811 7939
rect 5089 7905 5123 7939
rect 5356 7905 5390 7939
rect 7021 7905 7055 7939
rect 8033 7905 8067 7939
rect 9689 7905 9723 7939
rect 13553 7905 13587 7939
rect 21097 7905 21131 7939
rect 22753 7905 22787 7939
rect 23857 7905 23891 7939
rect 1869 7837 1903 7871
rect 1961 7837 1995 7871
rect 3157 7837 3191 7871
rect 4077 7837 4111 7871
rect 8125 7837 8159 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 15761 7837 15795 7871
rect 15945 7837 15979 7871
rect 17325 7837 17359 7871
rect 17417 7837 17451 7871
rect 18429 7837 18463 7871
rect 2421 7769 2455 7803
rect 7573 7769 7607 7803
rect 14657 7769 14691 7803
rect 16865 7769 16899 7803
rect 2789 7701 2823 7735
rect 4629 7701 4663 7735
rect 4905 7701 4939 7735
rect 7481 7701 7515 7735
rect 8953 7701 8987 7735
rect 11069 7701 11103 7735
rect 13645 7701 13679 7735
rect 15301 7701 15335 7735
rect 18061 7701 18095 7735
rect 18889 7701 18923 7735
rect 21281 7701 21315 7735
rect 22937 7701 22971 7735
rect 24041 7701 24075 7735
rect 1777 7497 1811 7531
rect 3525 7497 3559 7531
rect 5089 7497 5123 7531
rect 7665 7497 7699 7531
rect 7941 7497 7975 7531
rect 9321 7497 9355 7531
rect 12541 7497 12575 7531
rect 13737 7497 13771 7531
rect 14289 7497 14323 7531
rect 15761 7497 15795 7531
rect 16681 7497 16715 7531
rect 17325 7497 17359 7531
rect 21373 7497 21407 7531
rect 22753 7497 22787 7531
rect 7297 7429 7331 7463
rect 11897 7429 11931 7463
rect 16313 7429 16347 7463
rect 17693 7429 17727 7463
rect 24593 7429 24627 7463
rect 2237 7361 2271 7395
rect 2421 7361 2455 7395
rect 4077 7361 4111 7395
rect 5549 7361 5583 7395
rect 5641 7361 5675 7395
rect 6101 7361 6135 7395
rect 8401 7361 8435 7395
rect 8585 7361 8619 7395
rect 9965 7361 9999 7395
rect 10149 7361 10183 7395
rect 11345 7361 11379 7395
rect 13001 7361 13035 7395
rect 13093 7361 13127 7395
rect 14381 7361 14415 7395
rect 3893 7293 3927 7327
rect 4629 7293 4663 7327
rect 9045 7293 9079 7327
rect 9873 7293 9907 7327
rect 12173 7293 12207 7327
rect 18061 7293 18095 7327
rect 20545 7293 20579 7327
rect 21005 7293 21039 7327
rect 23673 7293 23707 7327
rect 24225 7293 24259 7327
rect 6653 7225 6687 7259
rect 8309 7225 8343 7259
rect 12909 7225 12943 7259
rect 14648 7225 14682 7259
rect 18328 7225 18362 7259
rect 1593 7157 1627 7191
rect 2145 7157 2179 7191
rect 2881 7157 2915 7191
rect 3433 7157 3467 7191
rect 3985 7157 4019 7191
rect 4997 7157 5031 7191
rect 5457 7157 5491 7191
rect 9505 7157 9539 7191
rect 10517 7157 10551 7191
rect 10977 7157 11011 7191
rect 16865 7157 16899 7191
rect 19441 7157 19475 7191
rect 20729 7157 20763 7191
rect 23857 7157 23891 7191
rect 2421 6953 2455 6987
rect 3525 6953 3559 6987
rect 5089 6953 5123 6987
rect 7297 6953 7331 6987
rect 7757 6953 7791 6987
rect 10057 6953 10091 6987
rect 12725 6953 12759 6987
rect 15117 6953 15151 6987
rect 16221 6953 16255 6987
rect 16957 6953 16991 6987
rect 18797 6953 18831 6987
rect 8217 6885 8251 6919
rect 9873 6885 9907 6919
rect 15485 6885 15519 6919
rect 2789 6817 2823 6851
rect 5621 6817 5655 6851
rect 10425 6817 10459 6851
rect 11989 6817 12023 6851
rect 13093 6817 13127 6851
rect 13553 6817 13587 6851
rect 17325 6817 17359 6851
rect 17684 6817 17718 6851
rect 22201 6817 22235 6851
rect 23949 6817 23983 6851
rect 1869 6749 1903 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 5365 6749 5399 6783
rect 8309 6749 8343 6783
rect 8493 6749 8527 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 12081 6749 12115 6783
rect 12173 6749 12207 6783
rect 13645 6749 13679 6783
rect 13829 6749 13863 6783
rect 16313 6749 16347 6783
rect 16497 6749 16531 6783
rect 17417 6749 17451 6783
rect 4629 6681 4663 6715
rect 9505 6681 9539 6715
rect 11529 6681 11563 6715
rect 13185 6681 13219 6715
rect 2145 6613 2179 6647
rect 4353 6613 4387 6647
rect 6745 6613 6779 6647
rect 7849 6613 7883 6647
rect 8861 6613 8895 6647
rect 11161 6613 11195 6647
rect 11621 6613 11655 6647
rect 14473 6613 14507 6647
rect 15853 6613 15887 6647
rect 22385 6613 22419 6647
rect 24133 6613 24167 6647
rect 3157 6409 3191 6443
rect 4169 6409 4203 6443
rect 9321 6409 9355 6443
rect 11253 6409 11287 6443
rect 14381 6409 14415 6443
rect 15025 6409 15059 6443
rect 19073 6409 19107 6443
rect 22569 6409 22603 6443
rect 24041 6409 24075 6443
rect 1777 6273 1811 6307
rect 4261 6273 4295 6307
rect 6285 6273 6319 6307
rect 7297 6273 7331 6307
rect 9873 6273 9907 6307
rect 15485 6273 15519 6307
rect 18521 6273 18555 6307
rect 18705 6273 18739 6307
rect 4517 6205 4551 6239
rect 7113 6205 7147 6239
rect 12173 6205 12207 6239
rect 12449 6205 12483 6239
rect 12716 6205 12750 6239
rect 15752 6205 15786 6239
rect 17877 6205 17911 6239
rect 18429 6205 18463 6239
rect 19441 6205 19475 6239
rect 19993 6205 20027 6239
rect 20453 6205 20487 6239
rect 21649 6205 21683 6239
rect 22201 6205 22235 6239
rect 2044 6137 2078 6171
rect 6653 6137 6687 6171
rect 7542 6137 7576 6171
rect 10140 6137 10174 6171
rect 1685 6069 1719 6103
rect 3801 6069 3835 6103
rect 5641 6069 5675 6103
rect 8677 6069 8711 6103
rect 9689 6069 9723 6103
rect 11805 6069 11839 6103
rect 13829 6069 13863 6103
rect 15393 6069 15427 6103
rect 16865 6069 16899 6103
rect 17509 6069 17543 6103
rect 18061 6069 18095 6103
rect 20177 6069 20211 6103
rect 21833 6069 21867 6103
rect 2881 5865 2915 5899
rect 4537 5865 4571 5899
rect 7757 5865 7791 5899
rect 8677 5865 8711 5899
rect 9505 5865 9539 5899
rect 9689 5865 9723 5899
rect 11161 5865 11195 5899
rect 12633 5865 12667 5899
rect 14013 5865 14047 5899
rect 14381 5865 14415 5899
rect 16037 5865 16071 5899
rect 16405 5865 16439 5899
rect 18061 5865 18095 5899
rect 3433 5797 3467 5831
rect 10149 5797 10183 5831
rect 10793 5797 10827 5831
rect 11520 5797 11554 5831
rect 13553 5797 13587 5831
rect 16948 5797 16982 5831
rect 18613 5797 18647 5831
rect 1501 5729 1535 5763
rect 1768 5729 1802 5763
rect 4445 5729 4479 5763
rect 6377 5729 6411 5763
rect 6633 5729 6667 5763
rect 10057 5729 10091 5763
rect 11253 5729 11287 5763
rect 14197 5729 14231 5763
rect 14657 5729 14691 5763
rect 15393 5729 15427 5763
rect 16681 5729 16715 5763
rect 19165 5729 19199 5763
rect 21005 5729 21039 5763
rect 4629 5661 4663 5695
rect 10241 5661 10275 5695
rect 15025 5661 15059 5695
rect 9137 5593 9171 5627
rect 3801 5525 3835 5559
rect 4077 5525 4111 5559
rect 5365 5525 5399 5559
rect 5733 5525 5767 5559
rect 6101 5525 6135 5559
rect 8401 5525 8435 5559
rect 13185 5525 13219 5559
rect 15577 5525 15611 5559
rect 19349 5525 19383 5559
rect 21189 5525 21223 5559
rect 1409 5321 1443 5355
rect 2881 5321 2915 5355
rect 4353 5321 4387 5355
rect 5273 5321 5307 5355
rect 6377 5321 6411 5355
rect 6837 5321 6871 5355
rect 7849 5321 7883 5355
rect 9781 5321 9815 5355
rect 11069 5321 11103 5355
rect 11897 5321 11931 5355
rect 13185 5321 13219 5355
rect 17325 5321 17359 5355
rect 19165 5321 19199 5355
rect 20913 5321 20947 5355
rect 4905 5253 4939 5287
rect 10701 5253 10735 5287
rect 16221 5253 16255 5287
rect 20637 5253 20671 5287
rect 21281 5253 21315 5287
rect 2053 5185 2087 5219
rect 2973 5185 3007 5219
rect 7481 5185 7515 5219
rect 13369 5185 13403 5219
rect 15761 5185 15795 5219
rect 16773 5185 16807 5219
rect 18613 5185 18647 5219
rect 1777 5117 1811 5151
rect 2421 5117 2455 5151
rect 3229 5117 3263 5151
rect 7297 5117 7331 5151
rect 8401 5117 8435 5151
rect 8668 5117 8702 5151
rect 16129 5117 16163 5151
rect 16589 5117 16623 5151
rect 18521 5117 18555 5151
rect 19993 5117 20027 5151
rect 21097 5117 21131 5151
rect 21557 5117 21591 5151
rect 22109 5117 22143 5151
rect 22569 5117 22603 5151
rect 8217 5049 8251 5083
rect 12909 5049 12943 5083
rect 13636 5049 13670 5083
rect 16681 5049 16715 5083
rect 18429 5049 18463 5083
rect 1869 4981 1903 5015
rect 5733 4981 5767 5015
rect 7205 4981 7239 5015
rect 10333 4981 10367 5015
rect 11345 4981 11379 5015
rect 12173 4981 12207 5015
rect 14749 4981 14783 5015
rect 15301 4981 15335 5015
rect 17785 4981 17819 5015
rect 18061 4981 18095 5015
rect 20177 4981 20211 5015
rect 22293 4981 22327 5015
rect 2329 4777 2363 4811
rect 2881 4777 2915 4811
rect 5089 4777 5123 4811
rect 5273 4777 5307 4811
rect 5733 4777 5767 4811
rect 6469 4777 6503 4811
rect 6837 4777 6871 4811
rect 7021 4777 7055 4811
rect 7573 4777 7607 4811
rect 8493 4777 8527 4811
rect 9689 4777 9723 4811
rect 10149 4777 10183 4811
rect 11345 4777 11379 4811
rect 11529 4777 11563 4811
rect 13553 4777 13587 4811
rect 15301 4777 15335 4811
rect 16405 4777 16439 4811
rect 16773 4777 16807 4811
rect 17325 4777 17359 4811
rect 18153 4777 18187 4811
rect 1409 4709 1443 4743
rect 3433 4709 3467 4743
rect 8401 4709 8435 4743
rect 9045 4709 9079 4743
rect 10057 4709 10091 4743
rect 15117 4709 15151 4743
rect 2789 4641 2823 4675
rect 5641 4641 5675 4675
rect 7849 4641 7883 4675
rect 9505 4641 9539 4675
rect 11897 4641 11931 4675
rect 13461 4641 13495 4675
rect 15669 4641 15703 4675
rect 17233 4641 17267 4675
rect 18429 4641 18463 4675
rect 19533 4641 19567 4675
rect 20913 4641 20947 4675
rect 21925 4641 21959 4675
rect 3065 4573 3099 4607
rect 4261 4573 4295 4607
rect 5917 4573 5951 4607
rect 8585 4573 8619 4607
rect 10241 4573 10275 4607
rect 10977 4573 11011 4607
rect 11989 4573 12023 4607
rect 12081 4573 12115 4607
rect 12541 4573 12575 4607
rect 13737 4573 13771 4607
rect 15761 4573 15795 4607
rect 15853 4573 15887 4607
rect 17509 4573 17543 4607
rect 2421 4505 2455 4539
rect 3801 4505 3835 4539
rect 13093 4505 13127 4539
rect 14473 4505 14507 4539
rect 16865 4505 16899 4539
rect 1869 4437 1903 4471
rect 4721 4437 4755 4471
rect 8033 4437 8067 4471
rect 12909 4437 12943 4471
rect 14197 4437 14231 4471
rect 18613 4437 18647 4471
rect 19717 4437 19751 4471
rect 21097 4437 21131 4471
rect 22109 4437 22143 4471
rect 2789 4233 2823 4267
rect 3433 4233 3467 4267
rect 4353 4233 4387 4267
rect 4905 4233 4939 4267
rect 8493 4233 8527 4267
rect 8585 4233 8619 4267
rect 11897 4233 11931 4267
rect 13829 4233 13863 4267
rect 17049 4233 17083 4267
rect 18613 4233 18647 4267
rect 20085 4233 20119 4267
rect 21189 4233 21223 4267
rect 22017 4233 22051 4267
rect 3709 4165 3743 4199
rect 4813 4097 4847 4131
rect 5457 4097 5491 4131
rect 6653 4097 6687 4131
rect 7757 4097 7791 4131
rect 11253 4165 11287 4199
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 14473 4097 14507 4131
rect 17325 4097 17359 4131
rect 1409 4029 1443 4063
rect 7665 4029 7699 4063
rect 8493 4029 8527 4063
rect 8769 4029 8803 4063
rect 9025 4029 9059 4063
rect 10701 4029 10735 4063
rect 11345 4029 11379 4063
rect 13553 4029 13587 4063
rect 14013 4029 14047 4063
rect 14841 4029 14875 4063
rect 15025 4029 15059 4063
rect 15292 4029 15326 4063
rect 18061 4029 18095 4063
rect 18981 4029 19015 4063
rect 19165 4029 19199 4063
rect 20269 4029 20303 4063
rect 21373 4029 21407 4063
rect 22477 4029 22511 4063
rect 22937 4029 22971 4063
rect 1676 3961 1710 3995
rect 5273 3961 5307 3995
rect 6009 3961 6043 3995
rect 7573 3961 7607 3995
rect 12817 3961 12851 3995
rect 19809 3961 19843 3995
rect 20913 3961 20947 3995
rect 3893 3893 3927 3927
rect 5365 3893 5399 3927
rect 7021 3893 7055 3927
rect 7205 3893 7239 3927
rect 8309 3893 8343 3927
rect 10149 3893 10183 3927
rect 11529 3893 11563 3927
rect 12173 3893 12207 3927
rect 12449 3893 12483 3927
rect 14197 3893 14231 3927
rect 16405 3893 16439 3927
rect 17693 3893 17727 3927
rect 18245 3893 18279 3927
rect 19349 3893 19383 3927
rect 20453 3893 20487 3927
rect 21557 3893 21591 3927
rect 22661 3893 22695 3927
rect 2881 3689 2915 3723
rect 3525 3689 3559 3723
rect 4261 3689 4295 3723
rect 4997 3689 5031 3723
rect 5273 3689 5307 3723
rect 6653 3689 6687 3723
rect 9137 3689 9171 3723
rect 10057 3689 10091 3723
rect 11161 3689 11195 3723
rect 13001 3689 13035 3723
rect 13921 3689 13955 3723
rect 15761 3689 15795 3723
rect 18245 3689 18279 3723
rect 19901 3689 19935 3723
rect 21373 3689 21407 3723
rect 1768 3621 1802 3655
rect 5733 3621 5767 3655
rect 7082 3621 7116 3655
rect 10517 3621 10551 3655
rect 11529 3621 11563 3655
rect 11888 3621 11922 3655
rect 13553 3621 13587 3655
rect 14749 3621 14783 3655
rect 20913 3621 20947 3655
rect 1501 3553 1535 3587
rect 5641 3553 5675 3587
rect 6837 3553 6871 3587
rect 10425 3553 10459 3587
rect 11621 3553 11655 3587
rect 14105 3553 14139 3587
rect 15669 3553 15703 3587
rect 17121 3553 17155 3587
rect 19349 3553 19383 3587
rect 23305 3553 23339 3587
rect 5917 3485 5951 3519
rect 9965 3485 9999 3519
rect 10701 3485 10735 3519
rect 15025 3485 15059 3519
rect 15853 3485 15887 3519
rect 16313 3485 16347 3519
rect 16865 3485 16899 3519
rect 8217 3417 8251 3451
rect 8861 3417 8895 3451
rect 3801 3349 3835 3383
rect 6377 3349 6411 3383
rect 14289 3349 14323 3383
rect 15301 3349 15335 3383
rect 16773 3349 16807 3383
rect 18797 3349 18831 3383
rect 19533 3349 19567 3383
rect 23489 3349 23523 3383
rect 1593 3145 1627 3179
rect 1961 3145 1995 3179
rect 2329 3145 2363 3179
rect 3893 3145 3927 3179
rect 4905 3145 4939 3179
rect 4997 3145 5031 3179
rect 6101 3145 6135 3179
rect 9689 3145 9723 3179
rect 10793 3145 10827 3179
rect 12173 3145 12207 3179
rect 15025 3145 15059 3179
rect 16865 3145 16899 3179
rect 17417 3145 17451 3179
rect 19625 3145 19659 3179
rect 20637 3145 20671 3179
rect 7021 3077 7055 3111
rect 8217 3077 8251 3111
rect 11805 3077 11839 3111
rect 15393 3077 15427 3111
rect 21373 3077 21407 3111
rect 23305 3077 23339 3111
rect 2513 3009 2547 3043
rect 5457 3009 5491 3043
rect 5641 3009 5675 3043
rect 7297 3009 7331 3043
rect 8309 3009 8343 3043
rect 10241 3009 10275 3043
rect 11253 3009 11287 3043
rect 11437 3009 11471 3043
rect 12449 3009 12483 3043
rect 15485 3009 15519 3043
rect 18613 3009 18647 3043
rect 19073 3009 19107 3043
rect 20177 3009 20211 3043
rect 2780 2941 2814 2975
rect 4537 2941 4571 2975
rect 6653 2941 6687 2975
rect 8576 2941 8610 2975
rect 12716 2941 12750 2975
rect 20085 2941 20119 2975
rect 21189 2941 21223 2975
rect 21649 2941 21683 2975
rect 22201 2941 22235 2975
rect 22661 2941 22695 2975
rect 24409 2941 24443 2975
rect 24961 2941 24995 2975
rect 5365 2873 5399 2907
rect 14657 2873 14691 2907
rect 15730 2873 15764 2907
rect 17877 2873 17911 2907
rect 18429 2873 18463 2907
rect 19533 2873 19567 2907
rect 19993 2873 20027 2907
rect 7757 2805 7791 2839
rect 10701 2805 10735 2839
rect 11161 2805 11195 2839
rect 13829 2805 13863 2839
rect 18061 2805 18095 2839
rect 18521 2805 18555 2839
rect 22385 2805 22419 2839
rect 24593 2805 24627 2839
rect 1409 2601 1443 2635
rect 1961 2601 1995 2635
rect 2789 2601 2823 2635
rect 5733 2601 5767 2635
rect 6745 2601 6779 2635
rect 8309 2601 8343 2635
rect 9597 2601 9631 2635
rect 10977 2601 11011 2635
rect 12081 2601 12115 2635
rect 12357 2601 12391 2635
rect 14289 2601 14323 2635
rect 16221 2601 16255 2635
rect 16405 2601 16439 2635
rect 18061 2601 18095 2635
rect 18797 2601 18831 2635
rect 19717 2601 19751 2635
rect 20453 2601 20487 2635
rect 24777 2601 24811 2635
rect 3709 2533 3743 2567
rect 3801 2533 3835 2567
rect 7196 2533 7230 2567
rect 16865 2533 16899 2567
rect 21189 2533 21223 2567
rect 23397 2533 23431 2567
rect 3525 2465 3559 2499
rect 4620 2465 4654 2499
rect 6377 2465 6411 2499
rect 6929 2465 6963 2499
rect 9229 2465 9263 2499
rect 9873 2465 9907 2499
rect 11345 2465 11379 2499
rect 12909 2465 12943 2499
rect 13176 2465 13210 2499
rect 14841 2465 14875 2499
rect 16773 2465 16807 2499
rect 18705 2465 18739 2499
rect 19901 2465 19935 2499
rect 20821 2465 20855 2499
rect 22937 2465 22971 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 3709 2397 3743 2431
rect 4353 2397 4387 2431
rect 11437 2397 11471 2431
rect 11621 2397 11655 2431
rect 15301 2397 15335 2431
rect 16957 2397 16991 2431
rect 18981 2397 19015 2431
rect 2421 2329 2455 2363
rect 17693 2329 17727 2363
rect 23121 2329 23155 2363
rect 2237 2261 2271 2295
rect 10057 2261 10091 2295
rect 10425 2261 10459 2295
rect 10793 2261 10827 2295
rect 15853 2261 15887 2295
rect 18337 2261 18371 2295
rect 20085 2261 20119 2295
<< metal1 >>
rect 3326 27072 3332 27124
rect 3384 27112 3390 27124
rect 6270 27112 6276 27124
rect 3384 27084 6276 27112
rect 3384 27072 3390 27084
rect 6270 27072 6276 27084
rect 6328 27072 6334 27124
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2498 24256 2504 24268
rect 1443 24228 2504 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2498 24216 2504 24228
rect 2556 24216 2562 24268
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1486 23808 1492 23860
rect 1544 23848 1550 23860
rect 1581 23851 1639 23857
rect 1581 23848 1593 23851
rect 1544 23820 1593 23848
rect 1544 23808 1550 23820
rect 1581 23817 1593 23820
rect 1627 23817 1639 23851
rect 2682 23848 2688 23860
rect 2643 23820 2688 23848
rect 1581 23811 1639 23817
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 2501 23647 2559 23653
rect 1443 23616 2084 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2056 23520 2084 23616
rect 2501 23613 2513 23647
rect 2547 23613 2559 23647
rect 2501 23607 2559 23613
rect 2516 23576 2544 23607
rect 3142 23576 3148 23588
rect 2516 23548 3148 23576
rect 3142 23536 3148 23548
rect 3200 23536 3206 23588
rect 2038 23508 2044 23520
rect 1999 23480 2044 23508
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2498 23508 2504 23520
rect 2455 23480 2504 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 2498 23468 2504 23480
rect 2556 23468 2562 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1394 23264 1400 23316
rect 1452 23304 1458 23316
rect 1581 23307 1639 23313
rect 1581 23304 1593 23307
rect 1452 23276 1593 23304
rect 1452 23264 1458 23276
rect 1581 23273 1593 23276
rect 1627 23273 1639 23307
rect 1581 23267 1639 23273
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2406 23168 2412 23180
rect 1443 23140 2412 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2406 23128 2412 23140
rect 2464 23128 2470 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 1670 22760 1676 22772
rect 1627 22732 1676 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 1670 22720 1676 22732
rect 1728 22720 1734 22772
rect 2038 22624 2044 22636
rect 1412 22596 2044 22624
rect 1412 22565 1440 22596
rect 2038 22584 2044 22596
rect 2096 22584 2102 22636
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22525 1455 22559
rect 1397 22519 1455 22525
rect 2406 22420 2412 22432
rect 2367 22392 2412 22420
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 1854 22080 1860 22092
rect 1443 22052 1860 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 1854 22040 1860 22052
rect 1912 22040 1918 22092
rect 1578 21944 1584 21956
rect 1539 21916 1584 21944
rect 1578 21904 1584 21916
rect 1636 21904 1642 21956
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1673 21335 1731 21341
rect 1673 21301 1685 21335
rect 1719 21332 1731 21335
rect 1854 21332 1860 21344
rect 1719 21304 1860 21332
rect 1719 21301 1731 21304
rect 1673 21295 1731 21301
rect 1854 21292 1860 21304
rect 1912 21292 1918 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1486 21088 1492 21140
rect 1544 21128 1550 21140
rect 1581 21131 1639 21137
rect 1581 21128 1593 21131
rect 1544 21100 1593 21128
rect 1544 21088 1550 21100
rect 1581 21097 1593 21100
rect 1627 21097 1639 21131
rect 1581 21091 1639 21097
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 1670 20992 1676 21004
rect 1443 20964 1676 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 1670 20952 1676 20964
rect 1728 20952 1734 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1670 20380 1676 20392
rect 1631 20352 1676 20380
rect 1670 20340 1676 20352
rect 1728 20340 1734 20392
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 1670 19904 1676 19916
rect 1443 19876 1676 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 1670 19864 1676 19876
rect 1728 19864 1734 19916
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 8113 19295 8171 19301
rect 8113 19261 8125 19295
rect 8159 19292 8171 19295
rect 8159 19264 8800 19292
rect 8159 19261 8171 19264
rect 8113 19255 8171 19261
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 8294 19156 8300 19168
rect 8255 19128 8300 19156
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8772 19165 8800 19264
rect 11606 19252 11612 19304
rect 11664 19292 11670 19304
rect 12066 19292 12072 19304
rect 11664 19264 12072 19292
rect 11664 19252 11670 19264
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12710 19252 12716 19304
rect 12768 19292 12774 19304
rect 13262 19292 13268 19304
rect 12768 19264 13268 19292
rect 12768 19252 12774 19264
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 8757 19159 8815 19165
rect 8757 19125 8769 19159
rect 8803 19156 8815 19159
rect 9950 19156 9956 19168
rect 8803 19128 9956 19156
rect 8803 19125 8815 19128
rect 8757 19119 8815 19125
rect 9950 19116 9956 19128
rect 10008 19116 10014 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 7742 18408 7748 18420
rect 7703 18380 7748 18408
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 7561 18207 7619 18213
rect 1443 18176 2084 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2056 18077 2084 18176
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 7607 18176 8248 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 8220 18080 8248 18176
rect 2041 18071 2099 18077
rect 2041 18037 2053 18071
rect 2087 18068 2099 18071
rect 2866 18068 2872 18080
rect 2087 18040 2872 18068
rect 2087 18037 2099 18040
rect 2041 18031 2099 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 8202 18068 8208 18080
rect 8163 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1394 17824 1400 17876
rect 1452 17864 1458 17876
rect 1581 17867 1639 17873
rect 1581 17864 1593 17867
rect 1452 17836 1593 17864
rect 1452 17824 1458 17836
rect 1581 17833 1593 17836
rect 1627 17833 1639 17867
rect 1581 17827 1639 17833
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1578 17728 1584 17740
rect 1443 17700 1584 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 2685 17255 2743 17261
rect 2685 17252 2697 17255
rect 1636 17224 2697 17252
rect 1636 17212 1642 17224
rect 2685 17221 2697 17224
rect 2731 17221 2743 17255
rect 2685 17215 2743 17221
rect 14274 17212 14280 17264
rect 14332 17252 14338 17264
rect 14734 17252 14740 17264
rect 14332 17224 14740 17252
rect 14332 17212 14338 17224
rect 14734 17212 14740 17224
rect 14792 17212 14798 17264
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2501 17119 2559 17125
rect 1443 17088 2084 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2056 16992 2084 17088
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 3050 17116 3056 17128
rect 2547 17088 3056 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 1486 16940 1492 16992
rect 1544 16980 1550 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 1544 16952 1593 16980
rect 1544 16940 1550 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 2038 16980 2044 16992
rect 1999 16952 2044 16980
rect 1581 16943 1639 16949
rect 2038 16940 2044 16952
rect 2096 16940 2102 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 5718 16776 5724 16788
rect 5679 16748 5724 16776
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 7466 16776 7472 16788
rect 7427 16748 7472 16776
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 6086 16640 6092 16652
rect 6047 16612 6092 16640
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6546 16640 6552 16652
rect 6227 16612 6552 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 7282 16640 7288 16652
rect 7243 16612 7288 16640
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 6362 16572 6368 16584
rect 6323 16544 6368 16572
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 5442 16232 5448 16244
rect 5403 16204 5448 16232
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6144 16204 6193 16232
rect 6144 16192 6150 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6546 16232 6552 16244
rect 6507 16204 6552 16232
rect 6181 16195 6239 16201
rect 6196 16096 6224 16195
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6196 16068 6837 16096
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 5261 16031 5319 16037
rect 5261 16028 5273 16031
rect 5184 16000 5273 16028
rect 5184 15904 5212 16000
rect 5261 15997 5273 16000
rect 5307 15997 5319 16031
rect 5261 15991 5319 15997
rect 5902 15960 5908 15972
rect 5863 15932 5908 15960
rect 5902 15920 5908 15932
rect 5960 15920 5966 15972
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 7282 15892 7288 15904
rect 7243 15864 7288 15892
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 5997 15691 6055 15697
rect 5997 15657 6009 15691
rect 6043 15688 6055 15691
rect 6546 15688 6552 15700
rect 6043 15660 6552 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 6270 15580 6276 15632
rect 6328 15620 6334 15632
rect 6365 15623 6423 15629
rect 6365 15620 6377 15623
rect 6328 15592 6377 15620
rect 6328 15580 6334 15592
rect 6365 15589 6377 15592
rect 6411 15589 6423 15623
rect 6365 15583 6423 15589
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 6604 15456 6649 15484
rect 6604 15444 6610 15456
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 4614 15348 4620 15360
rect 4387 15320 4620 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 6972 15320 7021 15348
rect 6972 15308 6978 15320
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 6546 15144 6552 15156
rect 5767 15116 6552 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 8168 15116 8217 15144
rect 8168 15104 8174 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 1394 15036 1400 15088
rect 1452 15076 1458 15088
rect 1673 15079 1731 15085
rect 1673 15076 1685 15079
rect 1452 15048 1685 15076
rect 1452 15036 1458 15048
rect 1673 15045 1685 15048
rect 1719 15076 1731 15079
rect 2593 15079 2651 15085
rect 2593 15076 2605 15079
rect 1719 15048 2605 15076
rect 1719 15045 1731 15048
rect 1673 15039 1731 15045
rect 2593 15045 2605 15048
rect 2639 15045 2651 15079
rect 2593 15039 2651 15045
rect 2961 15079 3019 15085
rect 2961 15045 2973 15079
rect 3007 15076 3019 15079
rect 4157 15079 4215 15085
rect 4157 15076 4169 15079
rect 3007 15048 4169 15076
rect 3007 15045 3019 15048
rect 2961 15039 3019 15045
rect 4157 15045 4169 15048
rect 4203 15045 4215 15079
rect 4157 15039 4215 15045
rect 2409 14943 2467 14949
rect 2409 14909 2421 14943
rect 2455 14940 2467 14943
rect 2976 14940 3004 15039
rect 6270 15036 6276 15088
rect 6328 15076 6334 15088
rect 6365 15079 6423 15085
rect 6365 15076 6377 15079
rect 6328 15048 6377 15076
rect 6328 15036 6334 15048
rect 6365 15045 6377 15048
rect 6411 15076 6423 15079
rect 6638 15076 6644 15088
rect 6411 15048 6644 15076
rect 6411 15045 6423 15048
rect 6365 15039 6423 15045
rect 6638 15036 6644 15048
rect 6696 15036 6702 15088
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 15008 3755 15011
rect 4706 15008 4712 15020
rect 3743 14980 4712 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 6822 15008 6828 15020
rect 6783 14980 6828 15008
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 2455 14912 3004 14940
rect 2455 14909 2467 14912
rect 2409 14903 2467 14909
rect 4065 14875 4123 14881
rect 4065 14841 4077 14875
rect 4111 14872 4123 14875
rect 4246 14872 4252 14884
rect 4111 14844 4252 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 4246 14832 4252 14844
rect 4304 14872 4310 14884
rect 4525 14875 4583 14881
rect 4525 14872 4537 14875
rect 4304 14844 4537 14872
rect 4304 14832 4310 14844
rect 4525 14841 4537 14844
rect 4571 14841 4583 14875
rect 4525 14835 4583 14841
rect 6546 14832 6552 14884
rect 6604 14872 6610 14884
rect 7070 14875 7128 14881
rect 7070 14872 7082 14875
rect 6604 14844 7082 14872
rect 6604 14832 6610 14844
rect 7070 14841 7082 14844
rect 7116 14841 7128 14875
rect 7070 14835 7128 14841
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 6089 14807 6147 14813
rect 6089 14773 6101 14807
rect 6135 14804 6147 14807
rect 6454 14804 6460 14816
rect 6135 14776 6460 14804
rect 6135 14773 6147 14776
rect 6089 14767 6147 14773
rect 6454 14764 6460 14776
rect 6512 14804 6518 14816
rect 7190 14804 7196 14816
rect 6512 14776 7196 14804
rect 6512 14764 6518 14776
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 1544 14572 1593 14600
rect 1544 14560 1550 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 4246 14600 4252 14612
rect 4207 14572 4252 14600
rect 1581 14563 1639 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6604 14572 6837 14600
rect 6604 14560 6610 14572
rect 6825 14569 6837 14572
rect 6871 14600 6883 14603
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 6871 14572 7389 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7377 14569 7389 14572
rect 7423 14569 7435 14603
rect 7377 14563 7435 14569
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 5534 14532 5540 14544
rect 4764 14504 5540 14532
rect 4764 14492 4770 14504
rect 5534 14492 5540 14504
rect 5592 14532 5598 14544
rect 5690 14535 5748 14541
rect 5690 14532 5702 14535
rect 5592 14504 5702 14532
rect 5592 14492 5598 14504
rect 5690 14501 5702 14504
rect 5736 14501 5748 14535
rect 5690 14495 5748 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2038 14464 2044 14476
rect 1443 14436 2044 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14464 5503 14467
rect 6730 14464 6736 14476
rect 5491 14436 6736 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 4672 14028 6837 14056
rect 4672 14016 4678 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 5629 13991 5687 13997
rect 5629 13988 5641 13991
rect 5592 13960 5641 13988
rect 5592 13948 5598 13960
rect 5629 13957 5641 13960
rect 5675 13957 5687 13991
rect 5629 13951 5687 13957
rect 6273 13991 6331 13997
rect 6273 13957 6285 13991
rect 6319 13988 6331 13991
rect 6730 13988 6736 14000
rect 6319 13960 6736 13988
rect 6319 13957 6331 13960
rect 6273 13951 6331 13957
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 4154 13920 4160 13932
rect 4067 13892 4160 13920
rect 4154 13880 4160 13892
rect 4212 13920 4218 13932
rect 4212 13892 4292 13920
rect 4212 13880 4218 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 2317 13855 2375 13861
rect 2317 13852 2329 13855
rect 1443 13824 2329 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 2317 13821 2329 13824
rect 2363 13852 2375 13855
rect 2682 13852 2688 13864
rect 2363 13824 2688 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 4264 13861 4292 13892
rect 3789 13855 3847 13861
rect 3789 13821 3801 13855
rect 3835 13852 3847 13855
rect 4249 13855 4307 13861
rect 3835 13824 4200 13852
rect 3835 13821 3847 13824
rect 3789 13815 3847 13821
rect 4172 13784 4200 13824
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 6288 13852 6316 13951
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 4295 13824 6316 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4494 13787 4552 13793
rect 4494 13784 4506 13787
rect 4172 13756 4506 13784
rect 4494 13753 4506 13756
rect 4540 13784 4552 13787
rect 5442 13784 5448 13796
rect 4540 13756 5448 13784
rect 4540 13753 4552 13756
rect 4494 13747 4552 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 7285 13787 7343 13793
rect 7285 13784 7297 13787
rect 6564 13756 7297 13784
rect 6564 13728 6592 13756
rect 7285 13753 7297 13756
rect 7331 13753 7343 13787
rect 7285 13747 7343 13753
rect 6546 13716 6552 13728
rect 6507 13688 6552 13716
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 6972 13688 7205 13716
rect 6972 13676 6978 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1394 13472 1400 13524
rect 1452 13512 1458 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 1452 13484 1593 13512
rect 1452 13472 1458 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 2682 13512 2688 13524
rect 2643 13484 2688 13512
rect 1581 13475 1639 13481
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 5442 13512 5448 13524
rect 5403 13484 5448 13512
rect 5442 13472 5448 13484
rect 5500 13512 5506 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 5500 13484 7205 13512
rect 5500 13472 5506 13484
rect 7193 13481 7205 13484
rect 7239 13512 7251 13515
rect 7374 13512 7380 13524
rect 7239 13484 7380 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 5997 13447 6055 13453
rect 5997 13444 6009 13447
rect 5592 13416 6009 13444
rect 5592 13404 5598 13416
rect 5997 13413 6009 13416
rect 6043 13413 6055 13447
rect 5997 13407 6055 13413
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 6914 13444 6920 13456
rect 6696 13416 6920 13444
rect 6696 13404 6702 13416
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2280 13348 2513 13376
rect 2280 13336 2286 13348
rect 2501 13345 2513 13348
rect 2547 13345 2559 13379
rect 2501 13339 2559 13345
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 4332 13379 4390 13385
rect 4332 13376 4344 13379
rect 3384 13348 4344 13376
rect 3384 13336 3390 13348
rect 4332 13345 4344 13348
rect 4378 13376 4390 13379
rect 5442 13376 5448 13388
rect 4378 13348 5448 13376
rect 4378 13345 4390 13348
rect 4332 13339 4390 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 4062 13308 4068 13320
rect 4023 13280 4068 13308
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 2317 13175 2375 13181
rect 2317 13141 2329 13175
rect 2363 13172 2375 13175
rect 2682 13172 2688 13184
rect 2363 13144 2688 13172
rect 2363 13141 2375 13144
rect 2317 13135 2375 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 3878 13172 3884 13184
rect 3839 13144 3884 13172
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 3326 12968 3332 12980
rect 3287 12940 3332 12968
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4120 12940 4813 12968
rect 4120 12928 4126 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 4801 12931 4859 12937
rect 3789 12903 3847 12909
rect 3789 12900 3801 12903
rect 2700 12872 3801 12900
rect 2700 12844 2728 12872
rect 3789 12869 3801 12872
rect 3835 12869 3847 12903
rect 3789 12863 3847 12869
rect 2682 12832 2688 12844
rect 2643 12804 2688 12832
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3326 12832 3332 12844
rect 2915 12804 3332 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 2314 12724 2320 12776
rect 2372 12764 2378 12776
rect 2884 12764 2912 12795
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4338 12832 4344 12844
rect 3936 12804 4344 12832
rect 3936 12792 3942 12804
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 4154 12764 4160 12776
rect 2372 12736 2912 12764
rect 4115 12736 4160 12764
rect 2372 12724 2378 12736
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 2133 12699 2191 12705
rect 2133 12665 2145 12699
rect 2179 12696 2191 12699
rect 2593 12699 2651 12705
rect 2593 12696 2605 12699
rect 2179 12668 2605 12696
rect 2179 12665 2191 12668
rect 2133 12659 2191 12665
rect 2593 12665 2605 12668
rect 2639 12696 2651 12699
rect 2774 12696 2780 12708
rect 2639 12668 2780 12696
rect 2639 12665 2651 12668
rect 2593 12659 2651 12665
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 3697 12631 3755 12637
rect 3697 12597 3709 12631
rect 3743 12628 3755 12631
rect 4246 12628 4252 12640
rect 3743 12600 4252 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 2314 12424 2320 12436
rect 2275 12396 2320 12424
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2961 12427 3019 12433
rect 2961 12424 2973 12427
rect 2832 12396 2973 12424
rect 2832 12384 2838 12396
rect 2961 12393 2973 12396
rect 3007 12393 3019 12427
rect 2961 12387 3019 12393
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 5166 12424 5172 12436
rect 4304 12396 5172 12424
rect 4304 12384 4310 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5442 12424 5448 12436
rect 5403 12396 5448 12424
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 2222 12316 2228 12368
rect 2280 12356 2286 12368
rect 4338 12365 4344 12368
rect 2593 12359 2651 12365
rect 2593 12356 2605 12359
rect 2280 12328 2605 12356
rect 2280 12316 2286 12328
rect 2593 12325 2605 12328
rect 2639 12325 2651 12359
rect 4332 12356 4344 12365
rect 4299 12328 4344 12356
rect 2593 12319 2651 12325
rect 4332 12319 4344 12328
rect 4338 12316 4344 12319
rect 4396 12316 4402 12368
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1578 12288 1584 12300
rect 1443 12260 1584 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 3970 12288 3976 12300
rect 3752 12260 3976 12288
rect 3752 12248 3758 12260
rect 3970 12248 3976 12260
rect 4028 12288 4034 12300
rect 12250 12297 12256 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 4028 12260 4077 12288
rect 4028 12248 4034 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 12244 12288 12256 12297
rect 12211 12260 12256 12288
rect 4065 12251 4123 12257
rect 12244 12251 12256 12260
rect 12250 12248 12256 12251
rect 12308 12248 12314 12300
rect 11974 12220 11980 12232
rect 11935 12192 11980 12220
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4062 12084 4068 12096
rect 3927 12056 4068 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 12768 12056 13369 12084
rect 12768 12044 12774 12056
rect 13357 12053 13369 12056
rect 13403 12053 13415 12087
rect 13357 12047 13415 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11880 1642 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 1636 11852 2145 11880
rect 1636 11840 1642 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 3694 11880 3700 11892
rect 3655 11852 3700 11880
rect 2133 11843 2191 11849
rect 3694 11840 3700 11852
rect 3752 11840 3758 11892
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 12250 11880 12256 11892
rect 12115 11852 12256 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 3712 11744 3740 11840
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 3712 11716 3801 11744
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 1995 11648 2544 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2516 11549 2544 11648
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 8846 11676 8852 11688
rect 2924 11648 8852 11676
rect 2924 11636 2930 11648
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 4062 11617 4068 11620
rect 3329 11611 3387 11617
rect 3329 11577 3341 11611
rect 3375 11608 3387 11611
rect 4056 11608 4068 11617
rect 3375 11580 4068 11608
rect 3375 11577 3387 11580
rect 3329 11571 3387 11577
rect 4056 11571 4068 11580
rect 4062 11568 4068 11571
rect 4120 11568 4126 11620
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2682 11540 2688 11552
rect 2547 11512 2688 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2682 11500 2688 11512
rect 2740 11500 2746 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 4396 11512 5181 11540
rect 4396 11500 4402 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 5169 11503 5227 11509
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 12713 11543 12771 11549
rect 12713 11540 12725 11543
rect 12032 11512 12725 11540
rect 12032 11500 12038 11512
rect 12713 11509 12725 11512
rect 12759 11540 12771 11543
rect 13170 11540 13176 11552
rect 12759 11512 13176 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3752 11308 3801 11336
rect 3752 11296 3758 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 4338 11336 4344 11348
rect 4299 11308 4344 11336
rect 3789 11299 3847 11305
rect 3804 11200 3832 11299
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 4430 11200 4436 11212
rect 3804 11172 4436 11200
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 4700 11203 4758 11209
rect 4700 11169 4712 11203
rect 4746 11200 4758 11203
rect 4982 11200 4988 11212
rect 4746 11172 4988 11200
rect 4746 11169 4758 11172
rect 4700 11163 4758 11169
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3602 11132 3608 11144
rect 3007 11104 3608 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 5813 11067 5871 11073
rect 5813 11064 5825 11067
rect 5500 11036 5825 11064
rect 5500 11024 5506 11036
rect 5813 11033 5825 11036
rect 5859 11033 5871 11067
rect 5813 11027 5871 11033
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3602 10792 3608 10804
rect 3563 10764 3608 10792
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4488 10764 4813 10792
rect 4488 10752 4494 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 2774 10684 2780 10736
rect 2832 10724 2838 10736
rect 3789 10727 3847 10733
rect 3789 10724 3801 10727
rect 2832 10696 3801 10724
rect 2832 10684 2838 10696
rect 3789 10693 3801 10696
rect 3835 10693 3847 10727
rect 3789 10687 3847 10693
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4120 10628 4445 10656
rect 4120 10616 4126 10628
rect 4433 10625 4445 10628
rect 4479 10656 4491 10659
rect 5442 10656 5448 10668
rect 4479 10628 5448 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 4157 10591 4215 10597
rect 4157 10588 4169 10591
rect 3660 10560 4169 10588
rect 3660 10548 3666 10560
rect 4157 10557 4169 10560
rect 4203 10557 4215 10591
rect 4157 10551 4215 10557
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 1636 10424 2421 10452
rect 1636 10412 1642 10424
rect 2409 10421 2421 10424
rect 2455 10452 2467 10455
rect 2498 10452 2504 10464
rect 2455 10424 2504 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 3329 10455 3387 10461
rect 3329 10421 3341 10455
rect 3375 10452 3387 10455
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 3375 10424 4261 10452
rect 3375 10421 3387 10424
rect 3329 10415 3387 10421
rect 4249 10421 4261 10424
rect 4295 10452 4307 10455
rect 4706 10452 4712 10464
rect 4295 10424 4712 10452
rect 4295 10421 4307 10424
rect 4249 10415 4307 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 5040 10424 5273 10452
rect 5040 10412 5046 10424
rect 5261 10421 5273 10424
rect 5307 10452 5319 10455
rect 5442 10452 5448 10464
rect 5307 10424 5448 10452
rect 5307 10421 5319 10424
rect 5261 10415 5319 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10452 8907 10455
rect 9674 10452 9680 10464
rect 8895 10424 9680 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 3881 10251 3939 10257
rect 3881 10217 3893 10251
rect 3927 10248 3939 10251
rect 4062 10248 4068 10260
rect 3927 10220 4068 10248
rect 3927 10217 3939 10220
rect 3881 10211 3939 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 6086 10248 6092 10260
rect 6047 10220 6092 10248
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7742 10248 7748 10260
rect 7703 10220 7748 10248
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 6181 10183 6239 10189
rect 6181 10149 6193 10183
rect 6227 10180 6239 10183
rect 6362 10180 6368 10192
rect 6227 10152 6368 10180
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 6362 10140 6368 10152
rect 6420 10140 6426 10192
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 2556 10084 2789 10112
rect 2556 10072 2562 10084
rect 2777 10081 2789 10084
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 6696 10084 7849 10112
rect 6696 10072 6702 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 17218 10121 17224 10124
rect 11221 10115 11279 10121
rect 11221 10112 11233 10115
rect 11112 10084 11233 10112
rect 11112 10072 11118 10084
rect 11221 10081 11233 10084
rect 11267 10081 11279 10115
rect 11221 10075 11279 10081
rect 17212 10075 17224 10121
rect 17276 10112 17282 10124
rect 17276 10084 17312 10112
rect 17218 10072 17224 10075
rect 17276 10072 17282 10084
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 7929 10047 7987 10053
rect 6411 10016 6960 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 2976 9976 3004 10007
rect 2832 9948 3004 9976
rect 5721 9979 5779 9985
rect 2832 9936 2838 9948
rect 5721 9945 5733 9979
rect 5767 9976 5779 9979
rect 6822 9976 6828 9988
rect 5767 9948 6828 9976
rect 5767 9945 5779 9948
rect 5721 9939 5779 9945
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 6932 9920 6960 10016
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 9858 10044 9864 10056
rect 9723 10016 9864 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 7285 9979 7343 9985
rect 7285 9945 7297 9979
rect 7331 9976 7343 9979
rect 7944 9976 7972 10007
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10962 10044 10968 10056
rect 10923 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 13814 10044 13820 10056
rect 13775 10016 13820 10044
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 8386 9976 8392 9988
rect 7331 9948 8392 9976
rect 7331 9945 7343 9948
rect 7285 9939 7343 9945
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 18322 9976 18328 9988
rect 18283 9948 18328 9976
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 1670 9908 1676 9920
rect 1631 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 1949 9911 2007 9917
rect 1949 9908 1961 9911
rect 1820 9880 1961 9908
rect 1820 9868 1826 9880
rect 1949 9877 1961 9880
rect 1995 9877 2007 9911
rect 1949 9871 2007 9877
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 5077 9911 5135 9917
rect 5077 9908 5089 9911
rect 4212 9880 5089 9908
rect 4212 9868 4218 9880
rect 5077 9877 5089 9880
rect 5123 9908 5135 9911
rect 5350 9908 5356 9920
rect 5123 9880 5356 9908
rect 5123 9877 5135 9880
rect 5077 9871 5135 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7377 9911 7435 9917
rect 7377 9877 7389 9911
rect 7423 9908 7435 9911
rect 8202 9908 8208 9920
rect 7423 9880 8208 9908
rect 7423 9877 7435 9880
rect 7377 9871 7435 9877
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 11882 9908 11888 9920
rect 11664 9880 11888 9908
rect 11664 9868 11670 9880
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12345 9911 12403 9917
rect 12345 9877 12357 9911
rect 12391 9908 12403 9911
rect 12434 9908 12440 9920
rect 12391 9880 12440 9908
rect 12391 9877 12403 9880
rect 12345 9871 12403 9877
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 13538 9908 13544 9920
rect 13403 9880 13544 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3053 9707 3111 9713
rect 3053 9704 3065 9707
rect 2924 9676 3065 9704
rect 2924 9664 2930 9676
rect 3053 9673 3065 9676
rect 3099 9704 3111 9707
rect 4065 9707 4123 9713
rect 4065 9704 4077 9707
rect 3099 9676 4077 9704
rect 3099 9673 3111 9676
rect 3053 9667 3111 9673
rect 4065 9673 4077 9676
rect 4111 9673 4123 9707
rect 4065 9667 4123 9673
rect 4706 9664 4712 9716
rect 4764 9704 4770 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4764 9676 4997 9704
rect 4764 9664 4770 9676
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 4985 9667 5043 9673
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 7190 9704 7196 9716
rect 6788 9676 7196 9704
rect 6788 9664 6794 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 11054 9704 11060 9716
rect 7800 9676 8248 9704
rect 11015 9676 11060 9704
rect 7800 9664 7806 9676
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 8220 9636 8248 9676
rect 11054 9664 11060 9676
rect 11112 9664 11118 9716
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17313 9707 17371 9713
rect 17313 9704 17325 9707
rect 17276 9676 17325 9704
rect 17276 9664 17282 9676
rect 17313 9673 17325 9676
rect 17359 9673 17371 9707
rect 17313 9667 17371 9673
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 4571 9608 5580 9636
rect 8220 9608 8769 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 5552 9580 5580 9608
rect 8757 9605 8769 9608
rect 8803 9605 8815 9639
rect 17328 9636 17356 9667
rect 18230 9636 18236 9648
rect 17328 9608 18236 9636
rect 8757 9599 8815 9605
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 3602 9568 3608 9580
rect 3563 9540 3608 9568
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5442 9568 5448 9580
rect 4939 9540 5448 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5592 9540 5641 9568
rect 5592 9528 5598 9540
rect 5629 9537 5641 9540
rect 5675 9568 5687 9571
rect 6178 9568 6184 9580
rect 5675 9540 6184 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9568 13323 9571
rect 13311 9540 13400 9568
rect 13311 9537 13323 9540
rect 13265 9531 13323 9537
rect 5350 9500 5356 9512
rect 5311 9472 5356 9500
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 9582 9500 9588 9512
rect 6871 9472 7236 9500
rect 9495 9472 9588 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7208 9444 7236 9472
rect 9582 9460 9588 9472
rect 9640 9500 9646 9512
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 9640 9472 9689 9500
rect 9640 9460 9646 9472
rect 9677 9469 9689 9472
rect 9723 9500 9735 9503
rect 10962 9500 10968 9512
rect 9723 9472 10968 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 13372 9500 13400 9540
rect 14366 9500 14372 9512
rect 13372 9472 14372 9500
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 3513 9435 3571 9441
rect 3513 9432 3525 9435
rect 3200 9404 3525 9432
rect 3200 9392 3206 9404
rect 3513 9401 3525 9404
rect 3559 9401 3571 9435
rect 3513 9395 3571 9401
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7070 9435 7128 9441
rect 7070 9432 7082 9435
rect 6972 9404 7082 9432
rect 6972 9392 6978 9404
rect 7070 9401 7082 9404
rect 7116 9401 7128 9435
rect 7070 9395 7128 9401
rect 7190 9392 7196 9444
rect 7248 9392 7254 9444
rect 9217 9435 9275 9441
rect 9217 9401 9229 9435
rect 9263 9432 9275 9435
rect 9922 9435 9980 9441
rect 9922 9432 9934 9435
rect 9263 9404 9934 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9922 9401 9934 9404
rect 9968 9432 9980 9435
rect 10042 9432 10048 9444
rect 9968 9404 10048 9432
rect 9968 9401 9980 9404
rect 9922 9395 9980 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 1946 9364 1952 9376
rect 1719 9336 1952 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2130 9364 2136 9376
rect 2087 9336 2136 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2501 9367 2559 9373
rect 2501 9333 2513 9367
rect 2547 9364 2559 9367
rect 2682 9364 2688 9376
rect 2547 9336 2688 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 2961 9367 3019 9373
rect 2961 9333 2973 9367
rect 3007 9364 3019 9367
rect 3326 9364 3332 9376
rect 3007 9336 3332 9364
rect 3007 9333 3019 9336
rect 2961 9327 3019 9333
rect 3326 9324 3332 9336
rect 3384 9364 3390 9376
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 3384 9336 3433 9364
rect 3384 9324 3390 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 3421 9327 3479 9333
rect 6089 9367 6147 9373
rect 6089 9333 6101 9367
rect 6135 9364 6147 9367
rect 6362 9364 6368 9376
rect 6135 9336 6368 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6638 9364 6644 9376
rect 6599 9336 6644 9364
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7432 9336 8217 9364
rect 7432 9324 7438 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11020 9336 11713 9364
rect 11020 9324 11026 9336
rect 11701 9333 11713 9336
rect 11747 9364 11759 9367
rect 12158 9364 12164 9376
rect 11747 9336 12164 9364
rect 11747 9333 11759 9336
rect 11701 9327 11759 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 13136 9336 13185 9364
rect 13136 9324 13142 9336
rect 13173 9333 13185 9336
rect 13219 9364 13231 9367
rect 13372 9364 13400 9472
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 13538 9441 13544 9444
rect 13532 9432 13544 9441
rect 13499 9404 13544 9432
rect 13532 9395 13544 9404
rect 13538 9392 13544 9395
rect 13596 9392 13602 9444
rect 13219 9336 13400 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 14332 9336 14657 9364
rect 14332 9324 14338 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 14645 9327 14703 9333
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17037 9367 17095 9373
rect 17037 9364 17049 9367
rect 17000 9336 17049 9364
rect 17000 9324 17006 9336
rect 17037 9333 17049 9336
rect 17083 9364 17095 9367
rect 17494 9364 17500 9376
rect 17083 9336 17500 9364
rect 17083 9333 17095 9336
rect 17037 9327 17095 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2038 9160 2044 9172
rect 1995 9132 2044 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 6086 9160 6092 9172
rect 6047 9132 6092 9160
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 8352 9132 9413 9160
rect 8352 9120 8358 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 7374 9101 7380 9104
rect 7368 9092 7380 9101
rect 7335 9064 7380 9092
rect 7368 9055 7380 9064
rect 7374 9052 7380 9055
rect 7432 9052 7438 9104
rect 2041 9027 2099 9033
rect 2041 8993 2053 9027
rect 2087 9024 2099 9027
rect 2314 9024 2320 9036
rect 2087 8996 2320 9024
rect 2087 8993 2099 8996
rect 2041 8987 2099 8993
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 4332 9027 4390 9033
rect 4332 8993 4344 9027
rect 4378 9024 4390 9027
rect 4614 9024 4620 9036
rect 4378 8996 4620 9024
rect 4378 8993 4390 8996
rect 4332 8987 4390 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 6963 8996 7113 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7101 8993 7113 8996
rect 7147 9024 7159 9027
rect 7190 9024 7196 9036
rect 7147 8996 7196 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 9416 9024 9444 9123
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 9732 9132 10057 9160
rect 9732 9120 9738 9132
rect 10045 9129 10057 9132
rect 10091 9160 10103 9163
rect 10134 9160 10140 9172
rect 10091 9132 10140 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9160 11118 9172
rect 11425 9163 11483 9169
rect 11425 9160 11437 9163
rect 11112 9132 11437 9160
rect 11112 9120 11118 9132
rect 11425 9129 11437 9132
rect 11471 9129 11483 9163
rect 14274 9160 14280 9172
rect 14235 9132 14280 9160
rect 11425 9123 11483 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 15654 9160 15660 9172
rect 15615 9132 15660 9160
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 9824 9064 10701 9092
rect 9824 9052 9830 9064
rect 10689 9061 10701 9064
rect 10735 9092 10747 9095
rect 10962 9092 10968 9104
rect 10735 9064 10968 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 12434 9101 12440 9104
rect 12428 9055 12440 9101
rect 12492 9092 12498 9104
rect 12492 9064 12528 9092
rect 12434 9052 12440 9055
rect 12492 9052 12498 9064
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 9416 8996 10149 9024
rect 10137 8993 10149 8996
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 9024 15807 9027
rect 16114 9024 16120 9036
rect 15795 8996 16120 9024
rect 15795 8993 15807 8996
rect 15749 8987 15807 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 22186 9024 22192 9036
rect 22147 8996 22192 9024
rect 22186 8984 22192 8996
rect 22244 8984 22250 9036
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2866 8956 2872 8968
rect 2188 8928 2872 8956
rect 2188 8916 2194 8928
rect 2866 8916 2872 8928
rect 2924 8956 2930 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 2924 8928 3433 8956
rect 2924 8916 2930 8928
rect 3421 8925 3433 8928
rect 3467 8956 3479 8959
rect 3602 8956 3608 8968
rect 3467 8928 3608 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 4028 8928 4077 8956
rect 4028 8916 4034 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 10042 8916 10048 8968
rect 10100 8956 10106 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 10100 8928 10241 8956
rect 10100 8916 10106 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 12158 8956 12164 8968
rect 12119 8928 12164 8956
rect 10229 8919 10287 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 15838 8956 15844 8968
rect 15799 8928 15844 8956
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 8481 8891 8539 8897
rect 8481 8888 8493 8891
rect 8444 8860 8493 8888
rect 8444 8848 8450 8860
rect 8481 8857 8493 8860
rect 8527 8857 8539 8891
rect 9674 8888 9680 8900
rect 9635 8860 9680 8888
rect 8481 8851 8539 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2593 8823 2651 8829
rect 2593 8820 2605 8823
rect 2280 8792 2605 8820
rect 2280 8780 2286 8792
rect 2593 8789 2605 8792
rect 2639 8789 2651 8823
rect 2593 8783 2651 8789
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 4246 8820 4252 8832
rect 3927 8792 4252 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4246 8780 4252 8792
rect 4304 8820 4310 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 4304 8792 5457 8820
rect 4304 8780 4310 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 6454 8820 6460 8832
rect 6415 8792 6460 8820
rect 5445 8783 5503 8789
rect 6454 8780 6460 8792
rect 6512 8820 6518 8832
rect 6914 8820 6920 8832
rect 6512 8792 6920 8820
rect 6512 8780 6518 8792
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 13538 8820 13544 8832
rect 13499 8792 13544 8820
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 15289 8823 15347 8829
rect 15289 8789 15301 8823
rect 15335 8820 15347 8823
rect 16482 8820 16488 8832
rect 15335 8792 16488 8820
rect 15335 8789 15347 8792
rect 15289 8783 15347 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 22373 8823 22431 8829
rect 22373 8789 22385 8823
rect 22419 8820 22431 8823
rect 23474 8820 23480 8832
rect 22419 8792 23480 8820
rect 22419 8789 22431 8792
rect 22373 8783 22431 8789
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 7374 8576 7380 8628
rect 7432 8616 7438 8628
rect 7653 8619 7711 8625
rect 7653 8616 7665 8619
rect 7432 8588 7665 8616
rect 7432 8576 7438 8588
rect 7653 8585 7665 8588
rect 7699 8616 7711 8619
rect 8110 8616 8116 8628
rect 7699 8588 8116 8616
rect 7699 8585 7711 8588
rect 7653 8579 7711 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 12492 8588 13461 8616
rect 12492 8576 12498 8588
rect 1394 8548 1400 8560
rect 1355 8520 1400 8548
rect 1394 8508 1400 8520
rect 1452 8508 1458 8560
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 9585 8551 9643 8557
rect 9585 8548 9597 8551
rect 9548 8520 9597 8548
rect 9548 8508 9554 8520
rect 9585 8517 9597 8520
rect 9631 8548 9643 8551
rect 10042 8548 10048 8560
rect 9631 8520 10048 8548
rect 9631 8517 9643 8520
rect 9585 8511 9643 8517
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 10689 8551 10747 8557
rect 10689 8517 10701 8551
rect 10735 8548 10747 8551
rect 10735 8520 12940 8548
rect 10735 8517 10747 8520
rect 10689 8511 10747 8517
rect 12912 8492 12940 8520
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 1857 8483 1915 8489
rect 1857 8480 1869 8483
rect 1728 8452 1869 8480
rect 1728 8440 1734 8452
rect 1857 8449 1869 8452
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2004 8452 2049 8480
rect 2004 8440 2010 8452
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 11112 8452 11253 8480
rect 11112 8440 11118 8452
rect 11241 8449 11253 8452
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 12216 8452 12265 8480
rect 12216 8440 12222 8452
rect 12253 8449 12265 8452
rect 12299 8480 12311 8483
rect 12894 8480 12900 8492
rect 12299 8452 12756 8480
rect 12807 8452 12900 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2777 8415 2835 8421
rect 2777 8412 2789 8415
rect 2096 8384 2789 8412
rect 2096 8372 2102 8384
rect 2777 8381 2789 8384
rect 2823 8381 2835 8415
rect 2777 8375 2835 8381
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 3881 8415 3939 8421
rect 3881 8412 3893 8415
rect 3559 8384 3893 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 3881 8381 3893 8384
rect 3927 8412 3939 8415
rect 3970 8412 3976 8424
rect 3927 8384 3976 8412
rect 3927 8381 3939 8384
rect 3881 8375 3939 8381
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 4246 8421 4252 8424
rect 4240 8412 4252 8421
rect 4120 8384 4252 8412
rect 4120 8372 4126 8384
rect 4240 8375 4252 8384
rect 4246 8372 4252 8375
rect 4304 8372 4310 8424
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 10643 8384 11161 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 11149 8381 11161 8384
rect 11195 8412 11207 8415
rect 12342 8412 12348 8424
rect 11195 8384 12348 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 2409 8347 2467 8353
rect 2409 8344 2421 8347
rect 2372 8316 2421 8344
rect 2372 8304 2378 8316
rect 2409 8313 2421 8316
rect 2455 8313 2467 8347
rect 3988 8344 4016 8372
rect 4430 8344 4436 8356
rect 3988 8316 4436 8344
rect 2409 8307 2467 8313
rect 4430 8304 4436 8316
rect 4488 8344 4494 8356
rect 5166 8344 5172 8356
rect 4488 8316 5172 8344
rect 4488 8304 4494 8316
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 6914 8344 6920 8356
rect 6871 8316 6920 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 5350 8276 5356 8288
rect 5311 8248 5356 8276
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 7377 8279 7435 8285
rect 7377 8276 7389 8279
rect 7248 8248 7389 8276
rect 7248 8236 7254 8248
rect 7377 8245 7389 8248
rect 7423 8276 7435 8279
rect 8113 8279 8171 8285
rect 8113 8276 8125 8279
rect 7423 8248 8125 8276
rect 7423 8245 7435 8248
rect 7377 8239 7435 8245
rect 8113 8245 8125 8248
rect 8159 8276 8171 8279
rect 8220 8276 8248 8375
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12728 8412 12756 8452
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13004 8489 13032 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 16485 8619 16543 8625
rect 16485 8616 16497 8619
rect 15712 8588 16497 8616
rect 15712 8576 15718 8588
rect 16485 8585 16497 8588
rect 16531 8585 16543 8619
rect 16485 8579 16543 8585
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 22244 8588 22477 8616
rect 22244 8576 22250 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22465 8579 22523 8585
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 17862 8548 17868 8560
rect 17083 8520 17868 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 17862 8508 17868 8520
rect 17920 8508 17926 8560
rect 21821 8551 21879 8557
rect 21821 8517 21833 8551
rect 21867 8548 21879 8551
rect 22094 8548 22100 8560
rect 21867 8520 22100 8548
rect 21867 8517 21879 8520
rect 21821 8511 21879 8517
rect 22094 8508 22100 8520
rect 22152 8508 22158 8560
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 12728 8384 14197 8412
rect 14185 8381 14197 8384
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 8386 8304 8392 8356
rect 8444 8353 8450 8356
rect 8444 8347 8508 8353
rect 8444 8313 8462 8347
rect 8496 8313 8508 8347
rect 8444 8307 8508 8313
rect 8444 8304 8450 8307
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11057 8347 11115 8353
rect 11057 8344 11069 8347
rect 11020 8316 11069 8344
rect 11020 8304 11026 8316
rect 11057 8313 11069 8316
rect 11103 8313 11115 8347
rect 11057 8307 11115 8313
rect 11885 8347 11943 8353
rect 11885 8313 11897 8347
rect 11931 8344 11943 8347
rect 12066 8344 12072 8356
rect 11931 8316 12072 8344
rect 11931 8313 11943 8316
rect 11885 8307 11943 8313
rect 12066 8304 12072 8316
rect 12124 8344 12130 8356
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 12124 8316 12817 8344
rect 12124 8304 12130 8316
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 12805 8307 12863 8313
rect 8294 8276 8300 8288
rect 8159 8248 8300 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 12437 8279 12495 8285
rect 12437 8245 12449 8279
rect 12483 8276 12495 8279
rect 12526 8276 12532 8288
rect 12483 8248 12532 8276
rect 12483 8245 12495 8248
rect 12437 8239 12495 8245
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 14093 8279 14151 8285
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14200 8276 14228 8375
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14441 8415 14499 8421
rect 14441 8412 14453 8415
rect 14332 8384 14453 8412
rect 14332 8372 14338 8384
rect 14441 8381 14453 8384
rect 14487 8381 14499 8415
rect 16850 8412 16856 8424
rect 16811 8384 16856 8412
rect 14441 8375 14499 8381
rect 16850 8372 16856 8384
rect 16908 8412 16914 8424
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 16908 8384 17325 8412
rect 16908 8372 16914 8384
rect 17313 8381 17325 8384
rect 17359 8381 17371 8415
rect 21634 8412 21640 8424
rect 21595 8384 21640 8412
rect 17313 8375 17371 8381
rect 21634 8372 21640 8384
rect 21692 8412 21698 8424
rect 22097 8415 22155 8421
rect 22097 8412 22109 8415
rect 21692 8384 22109 8412
rect 21692 8372 21698 8384
rect 22097 8381 22109 8384
rect 22143 8381 22155 8415
rect 22097 8375 22155 8381
rect 16114 8344 16120 8356
rect 16075 8316 16120 8344
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 14366 8276 14372 8288
rect 14139 8248 14372 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 15562 8276 15568 8288
rect 15523 8248 15568 8276
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 1762 8072 1768 8084
rect 1443 8044 1768 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 4062 8072 4068 8084
rect 3651 8044 4068 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 6454 8072 6460 8084
rect 6415 8044 6460 8072
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7650 8072 7656 8084
rect 6972 8044 7656 8072
rect 6972 8032 6978 8044
rect 7650 8032 7656 8044
rect 7708 8072 7714 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 7708 8044 7941 8072
rect 7708 8032 7714 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 7929 8035 7987 8041
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8444 8044 8585 8072
rect 8444 8032 8450 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 9490 8072 9496 8084
rect 9451 8044 9496 8072
rect 8573 8035 8631 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 12124 8044 12173 8072
rect 12124 8032 12130 8044
rect 12161 8041 12173 8044
rect 12207 8041 12219 8075
rect 12161 8035 12219 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12492 8044 12633 8072
rect 12492 8032 12498 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12952 8044 13001 8072
rect 12952 8032 12958 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14001 8075 14059 8081
rect 14001 8072 14013 8075
rect 13872 8044 14013 8072
rect 13872 8032 13878 8044
rect 14001 8041 14013 8044
rect 14047 8041 14059 8075
rect 15654 8072 15660 8084
rect 15615 8044 15660 8072
rect 14001 8035 14059 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 17218 8072 17224 8084
rect 17179 8044 17224 8072
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 9582 8004 9588 8016
rect 8352 7976 9588 8004
rect 8352 7964 8358 7976
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 9944 8007 10002 8013
rect 9944 7973 9956 8007
rect 9990 8004 10002 8007
rect 10134 8004 10140 8016
rect 9990 7976 10140 8004
rect 9990 7973 10002 7976
rect 9944 7967 10002 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 15105 8007 15163 8013
rect 15105 7973 15117 8007
rect 15151 8004 15163 8007
rect 15838 8004 15844 8016
rect 15151 7976 15844 8004
rect 15151 7973 15163 7976
rect 15105 7967 15163 7973
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 1762 7936 1768 7948
rect 1723 7908 1768 7936
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5166 7936 5172 7948
rect 5123 7908 5172 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5350 7945 5356 7948
rect 5344 7936 5356 7945
rect 5311 7908 5356 7936
rect 5344 7899 5356 7908
rect 5350 7896 5356 7899
rect 5408 7896 5414 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 6972 7908 7021 7936
rect 6972 7896 6978 7908
rect 7009 7905 7021 7908
rect 7055 7936 7067 7939
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 7055 7908 8033 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 8021 7905 8033 7908
rect 8067 7905 8079 7939
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 8021 7899 8079 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 21082 7936 21088 7948
rect 13587 7908 14320 7936
rect 21043 7908 21088 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 14292 7880 14320 7908
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22738 7936 22744 7948
rect 22152 7908 22744 7936
rect 22152 7896 22158 7908
rect 22738 7896 22744 7908
rect 22796 7896 22802 7948
rect 23842 7936 23848 7948
rect 23803 7908 23848 7936
rect 23842 7896 23848 7908
rect 23900 7896 23906 7948
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1636 7840 1869 7868
rect 1636 7828 1642 7840
rect 1857 7837 1869 7840
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 1964 7800 1992 7831
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2924 7840 3157 7868
rect 2924 7828 2930 7840
rect 3145 7837 3157 7840
rect 3191 7837 3203 7871
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 3145 7831 3203 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 12584 7840 14105 7868
rect 12584 7828 12590 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 14093 7831 14151 7837
rect 2409 7803 2467 7809
rect 2409 7800 2421 7803
rect 1964 7772 2421 7800
rect 2409 7769 2421 7772
rect 2455 7769 2467 7803
rect 7558 7800 7564 7812
rect 7519 7772 7564 7800
rect 2409 7763 2467 7769
rect 2424 7732 2452 7763
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 14108 7800 14136 7831
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 15746 7868 15752 7880
rect 15707 7840 15752 7868
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 15930 7868 15936 7880
rect 15891 7840 15936 7868
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 17310 7868 17316 7880
rect 17271 7840 17316 7868
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 18414 7868 18420 7880
rect 17460 7840 17505 7868
rect 18375 7840 18420 7868
rect 17460 7828 17466 7840
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 14645 7803 14703 7809
rect 14645 7800 14657 7803
rect 14108 7772 14657 7800
rect 14645 7769 14657 7772
rect 14691 7769 14703 7803
rect 14645 7763 14703 7769
rect 16853 7803 16911 7809
rect 16853 7769 16865 7803
rect 16899 7800 16911 7803
rect 17954 7800 17960 7812
rect 16899 7772 17960 7800
rect 16899 7769 16911 7772
rect 16853 7763 16911 7769
rect 17954 7760 17960 7772
rect 18012 7760 18018 7812
rect 2774 7732 2780 7744
rect 2424 7704 2780 7732
rect 2774 7692 2780 7704
rect 2832 7732 2838 7744
rect 4614 7732 4620 7744
rect 2832 7704 2925 7732
rect 4575 7704 4620 7732
rect 2832 7692 2838 7704
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 4890 7732 4896 7744
rect 4851 7704 4896 7732
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 8386 7732 8392 7744
rect 7515 7704 8392 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8938 7732 8944 7744
rect 8899 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 11054 7732 11060 7744
rect 11015 7704 11060 7732
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 13630 7732 13636 7744
rect 13591 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 15286 7732 15292 7744
rect 15247 7704 15292 7732
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 18046 7732 18052 7744
rect 18007 7704 18052 7732
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 18874 7732 18880 7744
rect 18835 7704 18880 7732
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 21269 7735 21327 7741
rect 21269 7701 21281 7735
rect 21315 7732 21327 7735
rect 22094 7732 22100 7744
rect 21315 7704 22100 7732
rect 21315 7701 21327 7704
rect 21269 7695 21327 7701
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22922 7732 22928 7744
rect 22883 7704 22928 7732
rect 22922 7692 22928 7704
rect 22980 7692 22986 7744
rect 24026 7732 24032 7744
rect 23987 7704 24032 7732
rect 24026 7692 24032 7704
rect 24084 7692 24090 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 1765 7531 1823 7537
rect 1765 7528 1777 7531
rect 1728 7500 1777 7528
rect 1728 7488 1734 7500
rect 1765 7497 1777 7500
rect 1811 7497 1823 7531
rect 1765 7491 1823 7497
rect 3513 7531 3571 7537
rect 3513 7497 3525 7531
rect 3559 7528 3571 7531
rect 4890 7528 4896 7540
rect 3559 7500 4896 7528
rect 3559 7497 3571 7500
rect 3513 7491 3571 7497
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 7650 7528 7656 7540
rect 7611 7500 7656 7528
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 9306 7528 9312 7540
rect 9267 7500 9312 7528
rect 9306 7488 9312 7500
rect 9364 7528 9370 7540
rect 9364 7500 9996 7528
rect 9364 7488 9370 7500
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2774 7392 2780 7404
rect 2455 7364 2780 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2774 7352 2780 7364
rect 2832 7392 2838 7404
rect 2958 7392 2964 7404
rect 2832 7364 2964 7392
rect 2832 7352 2838 7364
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 4028 7364 4077 7392
rect 4028 7352 4034 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4908 7392 4936 7488
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 7285 7463 7343 7469
rect 7285 7460 7297 7463
rect 6972 7432 7297 7460
rect 6972 7420 6978 7432
rect 7285 7429 7297 7432
rect 7331 7460 7343 7463
rect 7331 7432 8616 7460
rect 7331 7429 7343 7432
rect 7285 7423 7343 7429
rect 8588 7404 8616 7432
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 4908 7364 5549 7392
rect 4065 7355 4123 7361
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 6089 7395 6147 7401
rect 6089 7392 6101 7395
rect 5675 7364 6101 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6089 7361 6101 7364
rect 6135 7361 6147 7395
rect 8386 7392 8392 7404
rect 8347 7364 8392 7392
rect 6089 7355 6147 7361
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3568 7296 3893 7324
rect 3568 7284 3574 7296
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7324 4675 7327
rect 5350 7324 5356 7336
rect 4663 7296 5356 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 5350 7284 5356 7296
rect 5408 7324 5414 7336
rect 5644 7324 5672 7355
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8570 7392 8576 7404
rect 8531 7364 8576 7392
rect 8570 7352 8576 7364
rect 8628 7352 8634 7404
rect 9968 7401 9996 7500
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 12250 7528 12256 7540
rect 11756 7500 12256 7528
rect 11756 7488 11762 7500
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12526 7528 12532 7540
rect 12487 7500 12532 7528
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 13725 7531 13783 7537
rect 13725 7497 13737 7531
rect 13771 7528 13783 7531
rect 13814 7528 13820 7540
rect 13771 7500 13820 7528
rect 13771 7497 13783 7500
rect 13725 7491 13783 7497
rect 13814 7488 13820 7500
rect 13872 7488 13878 7540
rect 14277 7531 14335 7537
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 14366 7528 14372 7540
rect 14323 7500 14372 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 14366 7488 14372 7500
rect 14424 7528 14430 7540
rect 15470 7528 15476 7540
rect 14424 7500 15476 7528
rect 14424 7488 14430 7500
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15749 7531 15807 7537
rect 15749 7497 15761 7531
rect 15795 7528 15807 7531
rect 15838 7528 15844 7540
rect 15795 7500 15844 7528
rect 15795 7497 15807 7500
rect 15749 7491 15807 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 15988 7500 16681 7528
rect 15988 7488 15994 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 17310 7528 17316 7540
rect 17271 7500 17316 7528
rect 16669 7491 16727 7497
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 21361 7531 21419 7537
rect 21361 7528 21373 7531
rect 21140 7500 21373 7528
rect 21140 7488 21146 7500
rect 21361 7497 21373 7500
rect 21407 7497 21419 7531
rect 22738 7528 22744 7540
rect 22699 7500 22744 7528
rect 21361 7491 21419 7497
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 13538 7460 13544 7472
rect 11931 7432 13544 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 10134 7392 10140 7404
rect 10047 7364 10140 7392
rect 9953 7355 10011 7361
rect 10134 7352 10140 7364
rect 10192 7392 10198 7404
rect 10962 7392 10968 7404
rect 10192 7364 10968 7392
rect 10192 7352 10198 7364
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 12986 7392 12992 7404
rect 12947 7364 12992 7392
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13096 7401 13124 7432
rect 13538 7420 13544 7432
rect 13596 7420 13602 7472
rect 14384 7401 14412 7488
rect 15654 7420 15660 7472
rect 15712 7460 15718 7472
rect 16301 7463 16359 7469
rect 16301 7460 16313 7463
rect 15712 7432 16313 7460
rect 15712 7420 15718 7432
rect 16301 7429 16313 7432
rect 16347 7429 16359 7463
rect 16301 7423 16359 7429
rect 17218 7420 17224 7472
rect 17276 7460 17282 7472
rect 17681 7463 17739 7469
rect 17681 7460 17693 7463
rect 17276 7432 17693 7460
rect 17276 7420 17282 7432
rect 17681 7429 17693 7432
rect 17727 7429 17739 7463
rect 17681 7423 17739 7429
rect 23842 7420 23848 7472
rect 23900 7460 23906 7472
rect 24581 7463 24639 7469
rect 24581 7460 24593 7463
rect 23900 7432 24593 7460
rect 23900 7420 23906 7432
rect 24581 7429 24593 7432
rect 24627 7429 24639 7463
rect 24581 7423 24639 7429
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 14369 7395 14427 7401
rect 14369 7361 14381 7395
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 5408 7296 5672 7324
rect 9033 7327 9091 7333
rect 5408 7284 5414 7296
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9858 7324 9864 7336
rect 9079 7296 9864 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 12158 7324 12164 7336
rect 12119 7296 12164 7324
rect 12158 7284 12164 7296
rect 12216 7324 12222 7336
rect 13004 7324 13032 7352
rect 12216 7296 13032 7324
rect 12216 7284 12222 7296
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 18046 7324 18052 7336
rect 17552 7296 18052 7324
rect 17552 7284 17558 7296
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 20530 7324 20536 7336
rect 20491 7296 20536 7324
rect 20530 7284 20536 7296
rect 20588 7324 20594 7336
rect 20993 7327 21051 7333
rect 20993 7324 21005 7327
rect 20588 7296 21005 7324
rect 20588 7284 20594 7296
rect 20993 7293 21005 7296
rect 21039 7293 21051 7327
rect 20993 7287 21051 7293
rect 23474 7284 23480 7336
rect 23532 7324 23538 7336
rect 23661 7327 23719 7333
rect 23661 7324 23673 7327
rect 23532 7296 23673 7324
rect 23532 7284 23538 7296
rect 23661 7293 23673 7296
rect 23707 7324 23719 7327
rect 24213 7327 24271 7333
rect 24213 7324 24225 7327
rect 23707 7296 24225 7324
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 24213 7293 24225 7296
rect 24259 7293 24271 7327
rect 24213 7287 24271 7293
rect 6641 7259 6699 7265
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 8297 7259 8355 7265
rect 8297 7256 8309 7259
rect 6687 7228 8309 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 8297 7225 8309 7228
rect 8343 7256 8355 7259
rect 8343 7228 9536 7256
rect 8343 7225 8355 7228
rect 8297 7219 8355 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 2130 7188 2136 7200
rect 2091 7160 2136 7188
rect 2130 7148 2136 7160
rect 2188 7148 2194 7200
rect 2406 7148 2412 7200
rect 2464 7188 2470 7200
rect 2869 7191 2927 7197
rect 2869 7188 2881 7191
rect 2464 7160 2881 7188
rect 2464 7148 2470 7160
rect 2869 7157 2881 7160
rect 2915 7188 2927 7191
rect 3142 7188 3148 7200
rect 2915 7160 3148 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 3970 7188 3976 7200
rect 3467 7160 3976 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4985 7191 5043 7197
rect 4985 7157 4997 7191
rect 5031 7188 5043 7191
rect 5166 7188 5172 7200
rect 5031 7160 5172 7188
rect 5031 7157 5043 7160
rect 4985 7151 5043 7157
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5442 7188 5448 7200
rect 5403 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 9508 7197 9536 7228
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 12897 7259 12955 7265
rect 12897 7256 12909 7259
rect 12860 7228 12909 7256
rect 12860 7216 12866 7228
rect 12897 7225 12909 7228
rect 12943 7225 12955 7259
rect 12897 7219 12955 7225
rect 14636 7259 14694 7265
rect 14636 7225 14648 7259
rect 14682 7256 14694 7259
rect 14826 7256 14832 7268
rect 14682 7228 14832 7256
rect 14682 7225 14694 7228
rect 14636 7219 14694 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 18316 7259 18374 7265
rect 18316 7225 18328 7259
rect 18362 7256 18374 7259
rect 18874 7256 18880 7268
rect 18362 7228 18880 7256
rect 18362 7225 18374 7228
rect 18316 7219 18374 7225
rect 18874 7216 18880 7228
rect 18932 7216 18938 7268
rect 9493 7191 9551 7197
rect 9493 7157 9505 7191
rect 9539 7157 9551 7191
rect 9493 7151 9551 7157
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10505 7191 10563 7197
rect 10505 7188 10517 7191
rect 9824 7160 10517 7188
rect 9824 7148 9830 7160
rect 10505 7157 10517 7160
rect 10551 7157 10563 7191
rect 10962 7188 10968 7200
rect 10923 7160 10968 7188
rect 10505 7151 10563 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 16850 7188 16856 7200
rect 16811 7160 16856 7188
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 19426 7188 19432 7200
rect 19387 7160 19432 7188
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 20714 7188 20720 7200
rect 20675 7160 20720 7188
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 23842 7188 23848 7200
rect 23803 7160 23848 7188
rect 23842 7148 23848 7160
rect 23900 7148 23906 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 2188 6956 2421 6984
rect 2188 6944 2194 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 3510 6984 3516 6996
rect 3471 6956 3516 6984
rect 2409 6947 2467 6953
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1857 6783 1915 6789
rect 1857 6780 1869 6783
rect 1728 6752 1869 6780
rect 1728 6740 1734 6752
rect 1857 6749 1869 6752
rect 1903 6780 1915 6783
rect 1903 6752 2360 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 1912 6616 2145 6644
rect 1912 6604 1918 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 2332 6644 2360 6752
rect 2424 6712 2452 6947
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 5077 6987 5135 6993
rect 5077 6984 5089 6987
rect 4120 6956 5089 6984
rect 4120 6944 4126 6956
rect 5077 6953 5089 6956
rect 5123 6984 5135 6987
rect 5442 6984 5448 6996
rect 5123 6956 5448 6984
rect 5123 6953 5135 6956
rect 5077 6947 5135 6953
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 7248 6956 7297 6984
rect 7248 6944 7254 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 7745 6987 7803 6993
rect 7745 6953 7757 6987
rect 7791 6984 7803 6987
rect 8110 6984 8116 6996
rect 7791 6956 8116 6984
rect 7791 6953 7803 6956
rect 7745 6947 7803 6953
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 8444 6956 10057 6984
rect 8444 6944 8450 6956
rect 10045 6953 10057 6956
rect 10091 6953 10103 6987
rect 10045 6947 10103 6953
rect 12713 6987 12771 6993
rect 12713 6953 12725 6987
rect 12759 6984 12771 6987
rect 12802 6984 12808 6996
rect 12759 6956 12808 6984
rect 12759 6953 12771 6956
rect 12713 6947 12771 6953
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15746 6984 15752 6996
rect 15151 6956 15752 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 8202 6916 8208 6928
rect 8163 6888 8208 6916
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9861 6919 9919 6925
rect 9861 6916 9873 6919
rect 9824 6888 9873 6916
rect 9824 6876 9830 6888
rect 9861 6885 9873 6888
rect 9907 6885 9919 6919
rect 9861 6879 9919 6885
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 3878 6848 3884 6860
rect 2823 6820 3884 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5609 6851 5667 6857
rect 5609 6848 5621 6851
rect 5500 6820 5621 6848
rect 5500 6808 5506 6820
rect 5609 6817 5621 6820
rect 5655 6817 5667 6851
rect 5609 6811 5667 6817
rect 6748 6820 8524 6848
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 2869 6783 2927 6789
rect 2869 6780 2881 6783
rect 2556 6752 2881 6780
rect 2556 6740 2562 6752
rect 2869 6749 2881 6752
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3142 6780 3148 6792
rect 3099 6752 3148 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 5166 6740 5172 6792
rect 5224 6780 5230 6792
rect 5353 6783 5411 6789
rect 5353 6780 5365 6783
rect 5224 6752 5365 6780
rect 5224 6740 5230 6752
rect 5353 6749 5365 6752
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 4617 6715 4675 6721
rect 4617 6712 4629 6715
rect 2424 6684 4629 6712
rect 4617 6681 4629 6684
rect 4663 6681 4675 6715
rect 4617 6675 4675 6681
rect 3234 6644 3240 6656
rect 2332 6616 3240 6644
rect 2133 6607 2191 6613
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 4338 6644 4344 6656
rect 4299 6616 4344 6644
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 5368 6644 5396 6743
rect 6270 6644 6276 6656
rect 5368 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 6748 6653 6776 6820
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 6972 6752 8309 6780
rect 6972 6740 6978 6752
rect 8297 6749 8309 6752
rect 8343 6780 8355 6783
rect 8386 6780 8392 6792
rect 8343 6752 8392 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8496 6789 8524 6820
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10413 6851 10471 6857
rect 10413 6848 10425 6851
rect 9732 6820 10425 6848
rect 9732 6808 9738 6820
rect 10413 6817 10425 6820
rect 10459 6817 10471 6851
rect 10870 6848 10876 6860
rect 10413 6811 10471 6817
rect 10520 6820 10876 6848
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6780 8539 6783
rect 8570 6780 8576 6792
rect 8527 6752 8576 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 10520 6789 10548 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 13078 6848 13084 6860
rect 13039 6820 13084 6848
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 13538 6848 13544 6860
rect 13499 6820 13544 6848
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 9364 6752 10517 6780
rect 9364 6740 9370 6752
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10962 6780 10968 6792
rect 10735 6752 10968 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 9490 6712 9496 6724
rect 9403 6684 9496 6712
rect 9490 6672 9496 6684
rect 9548 6712 9554 6724
rect 10704 6712 10732 6743
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 11204 6752 12081 6780
rect 11204 6740 11210 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12161 6743 12219 6749
rect 9548 6684 10732 6712
rect 9548 6672 9554 6684
rect 10778 6672 10784 6724
rect 10836 6712 10842 6724
rect 11517 6715 11575 6721
rect 11517 6712 11529 6715
rect 10836 6684 11529 6712
rect 10836 6672 10842 6684
rect 11517 6681 11529 6684
rect 11563 6712 11575 6715
rect 12176 6712 12204 6743
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 13630 6780 13636 6792
rect 12492 6752 13636 6780
rect 12492 6740 12498 6752
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13814 6780 13820 6792
rect 13775 6752 13820 6780
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 11563 6684 12204 6712
rect 13173 6715 13231 6721
rect 11563 6681 11575 6684
rect 11517 6675 11575 6681
rect 13173 6681 13185 6715
rect 13219 6712 13231 6715
rect 15120 6712 15148 6947
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 16206 6984 16212 6996
rect 16167 6956 16212 6984
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 16942 6984 16948 6996
rect 16855 6956 16948 6984
rect 16942 6944 16948 6956
rect 17000 6984 17006 6996
rect 17402 6984 17408 6996
rect 17000 6956 17408 6984
rect 17000 6944 17006 6956
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 18785 6987 18843 6993
rect 18785 6953 18797 6987
rect 18831 6984 18843 6987
rect 18874 6984 18880 6996
rect 18831 6956 18880 6984
rect 18831 6953 18843 6956
rect 18785 6947 18843 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 15470 6916 15476 6928
rect 15431 6888 15476 6916
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 16500 6820 17325 6848
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16500 6789 16528 6820
rect 17313 6817 17325 6820
rect 17359 6848 17371 6851
rect 17672 6851 17730 6857
rect 17672 6848 17684 6851
rect 17359 6820 17684 6848
rect 17359 6817 17371 6820
rect 17313 6811 17371 6817
rect 17672 6817 17684 6820
rect 17718 6848 17730 6851
rect 18046 6848 18052 6860
rect 17718 6820 18052 6848
rect 17718 6817 17730 6820
rect 17672 6811 17730 6817
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 22094 6808 22100 6860
rect 22152 6848 22158 6860
rect 22189 6851 22247 6857
rect 22189 6848 22201 6851
rect 22152 6820 22201 6848
rect 22152 6808 22158 6820
rect 22189 6817 22201 6820
rect 22235 6848 22247 6851
rect 22554 6848 22560 6860
rect 22235 6820 22560 6848
rect 22235 6817 22247 6820
rect 22189 6811 22247 6817
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6848 23995 6851
rect 24026 6848 24032 6860
rect 23983 6820 24032 6848
rect 23983 6817 23995 6820
rect 23937 6811 23995 6817
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 15988 6752 16313 6780
rect 15988 6740 15994 6752
rect 16301 6749 16313 6752
rect 16347 6749 16359 6783
rect 16301 6743 16359 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 17402 6780 17408 6792
rect 17363 6752 17408 6780
rect 16485 6743 16543 6749
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 13219 6684 15148 6712
rect 13219 6681 13231 6684
rect 13173 6675 13231 6681
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6512 6616 6745 6644
rect 6512 6604 6518 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 7834 6644 7840 6656
rect 7795 6616 7840 6644
rect 6733 6607 6791 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8849 6647 8907 6653
rect 8849 6644 8861 6647
rect 8352 6616 8861 6644
rect 8352 6604 8358 6616
rect 8849 6613 8861 6616
rect 8895 6613 8907 6647
rect 8849 6607 8907 6613
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6644 11207 6647
rect 11238 6644 11244 6656
rect 11195 6616 11244 6644
rect 11195 6613 11207 6616
rect 11149 6607 11207 6613
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11606 6644 11612 6656
rect 11567 6616 11612 6644
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 14461 6647 14519 6653
rect 14461 6613 14473 6647
rect 14507 6644 14519 6647
rect 14826 6644 14832 6656
rect 14507 6616 14832 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15838 6644 15844 6656
rect 15799 6616 15844 6644
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 22370 6644 22376 6656
rect 22331 6616 22376 6644
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 24118 6644 24124 6656
rect 24079 6616 24124 6644
rect 24118 6604 24124 6616
rect 24176 6604 24182 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3145 6443 3203 6449
rect 3145 6440 3157 6443
rect 3108 6412 3157 6440
rect 3108 6400 3114 6412
rect 3145 6409 3157 6412
rect 3191 6409 3203 6443
rect 3145 6403 3203 6409
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 5166 6440 5172 6452
rect 4203 6412 5172 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1728 6276 1777 6304
rect 1728 6264 1734 6276
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 3234 6264 3240 6316
rect 3292 6304 3298 6316
rect 4264 6313 4292 6412
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 9306 6440 9312 6452
rect 9267 6412 9312 6440
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 11241 6443 11299 6449
rect 11241 6409 11253 6443
rect 11287 6440 11299 6443
rect 11514 6440 11520 6452
rect 11287 6412 11520 6440
rect 11287 6409 11299 6412
rect 11241 6403 11299 6409
rect 11514 6400 11520 6412
rect 11572 6440 11578 6452
rect 13814 6440 13820 6452
rect 11572 6412 13820 6440
rect 11572 6400 11578 6412
rect 13814 6400 13820 6412
rect 13872 6440 13878 6452
rect 14369 6443 14427 6449
rect 14369 6440 14381 6443
rect 13872 6412 14381 6440
rect 13872 6400 13878 6412
rect 14369 6409 14381 6412
rect 14415 6409 14427 6443
rect 14369 6403 14427 6409
rect 15013 6443 15071 6449
rect 15013 6409 15025 6443
rect 15059 6440 15071 6443
rect 15746 6440 15752 6452
rect 15059 6412 15752 6440
rect 15059 6409 15071 6412
rect 15013 6403 15071 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 18874 6400 18880 6452
rect 18932 6440 18938 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18932 6412 19073 6440
rect 18932 6400 18938 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 22554 6440 22560 6452
rect 22515 6412 22560 6440
rect 19061 6403 19119 6409
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 24026 6440 24032 6452
rect 23987 6412 24032 6440
rect 24026 6400 24032 6412
rect 24084 6400 24090 6452
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 3292 6276 4261 6304
rect 3292 6264 3298 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 6270 6304 6276 6316
rect 6183 6276 6276 6304
rect 4249 6267 4307 6273
rect 6270 6264 6276 6276
rect 6328 6304 6334 6316
rect 7190 6304 7196 6316
rect 6328 6276 7196 6304
rect 6328 6264 6334 6276
rect 7190 6264 7196 6276
rect 7248 6304 7254 6316
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7248 6276 7297 6304
rect 7248 6264 7254 6276
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 9858 6304 9864 6316
rect 9819 6276 9864 6304
rect 7285 6267 7343 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 15470 6304 15476 6316
rect 15431 6276 15476 6304
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 18506 6304 18512 6316
rect 18467 6276 18512 6304
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 18892 6304 18920 6400
rect 18739 6276 18920 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 842 6196 848 6248
rect 900 6236 906 6248
rect 900 6208 4292 6236
rect 900 6196 906 6208
rect 2032 6171 2090 6177
rect 2032 6137 2044 6171
rect 2078 6168 2090 6171
rect 2866 6168 2872 6180
rect 2078 6140 2872 6168
rect 2078 6137 2090 6140
rect 2032 6131 2090 6137
rect 2866 6128 2872 6140
rect 2924 6128 2930 6180
rect 4264 6168 4292 6208
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4505 6239 4563 6245
rect 4505 6236 4517 6239
rect 4396 6208 4517 6236
rect 4396 6196 4402 6208
rect 4505 6205 4517 6208
rect 4551 6205 4563 6239
rect 6362 6236 6368 6248
rect 6275 6208 6368 6236
rect 4505 6199 4563 6205
rect 6362 6196 6368 6208
rect 6420 6236 6426 6248
rect 6914 6236 6920 6248
rect 6420 6208 6920 6236
rect 6420 6196 6426 6208
rect 6914 6196 6920 6208
rect 6972 6236 6978 6248
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 6972 6208 7113 6236
rect 6972 6196 6978 6208
rect 7101 6205 7113 6208
rect 7147 6205 7159 6239
rect 9876 6236 9904 6264
rect 10962 6236 10968 6248
rect 9876 6208 10968 6236
rect 7101 6199 7159 6205
rect 10962 6196 10968 6208
rect 11020 6236 11026 6248
rect 11882 6236 11888 6248
rect 11020 6208 11888 6236
rect 11020 6196 11026 6208
rect 11882 6196 11888 6208
rect 11940 6236 11946 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11940 6208 12173 6236
rect 11940 6196 11946 6208
rect 12161 6205 12173 6208
rect 12207 6236 12219 6239
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12207 6208 12449 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 12704 6239 12762 6245
rect 12704 6205 12716 6239
rect 12750 6236 12762 6239
rect 13078 6236 13084 6248
rect 12750 6208 13084 6236
rect 12750 6205 12762 6208
rect 12704 6199 12762 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 15746 6245 15752 6248
rect 15740 6236 15752 6245
rect 15707 6208 15752 6236
rect 15740 6199 15752 6208
rect 15746 6196 15752 6199
rect 15804 6196 15810 6248
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 18414 6236 18420 6248
rect 17911 6208 18420 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 18524 6236 18552 6264
rect 19429 6239 19487 6245
rect 19429 6236 19441 6239
rect 18524 6208 19441 6236
rect 19429 6205 19441 6208
rect 19475 6205 19487 6239
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 19429 6199 19487 6205
rect 19978 6196 19984 6208
rect 20036 6236 20042 6248
rect 20441 6239 20499 6245
rect 20441 6236 20453 6239
rect 20036 6208 20453 6236
rect 20036 6196 20042 6208
rect 20441 6205 20453 6208
rect 20487 6205 20499 6239
rect 20441 6199 20499 6205
rect 20714 6196 20720 6248
rect 20772 6236 20778 6248
rect 21637 6239 21695 6245
rect 21637 6236 21649 6239
rect 20772 6208 21649 6236
rect 20772 6196 20778 6208
rect 21637 6205 21649 6208
rect 21683 6236 21695 6239
rect 22189 6239 22247 6245
rect 22189 6236 22201 6239
rect 21683 6208 22201 6236
rect 21683 6205 21695 6208
rect 21637 6199 21695 6205
rect 22189 6205 22201 6208
rect 22235 6205 22247 6239
rect 22189 6199 22247 6205
rect 6380 6168 6408 6196
rect 4264 6140 6408 6168
rect 6641 6171 6699 6177
rect 6641 6137 6653 6171
rect 6687 6168 6699 6171
rect 7530 6171 7588 6177
rect 7530 6168 7542 6171
rect 6687 6140 7542 6168
rect 6687 6137 6699 6140
rect 6641 6131 6699 6137
rect 7530 6137 7542 6140
rect 7576 6168 7588 6171
rect 7742 6168 7748 6180
rect 7576 6140 7748 6168
rect 7576 6137 7588 6140
rect 7530 6131 7588 6137
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 10128 6171 10186 6177
rect 10128 6137 10140 6171
rect 10174 6168 10186 6171
rect 10778 6168 10784 6180
rect 10174 6140 10784 6168
rect 10174 6137 10186 6140
rect 10128 6131 10186 6137
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 18322 6168 18328 6180
rect 17512 6140 18328 6168
rect 17512 6112 17540 6140
rect 18322 6128 18328 6140
rect 18380 6128 18386 6180
rect 1673 6103 1731 6109
rect 1673 6069 1685 6103
rect 1719 6100 1731 6103
rect 2498 6100 2504 6112
rect 1719 6072 2504 6100
rect 1719 6069 1731 6072
rect 1673 6063 1731 6069
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 3878 6100 3884 6112
rect 3835 6072 3884 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 5408 6072 5641 6100
rect 5408 6060 5414 6072
rect 5629 6069 5641 6072
rect 5675 6069 5687 6103
rect 8662 6100 8668 6112
rect 8623 6072 8668 6100
rect 5629 6063 5687 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 9674 6100 9680 6112
rect 9635 6072 9680 6100
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11388 6072 11805 6100
rect 11388 6060 11394 6072
rect 11793 6069 11805 6072
rect 11839 6100 11851 6103
rect 11974 6100 11980 6112
rect 11839 6072 11980 6100
rect 11839 6069 11851 6072
rect 11793 6063 11851 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 15381 6103 15439 6109
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 15930 6100 15936 6112
rect 15427 6072 15936 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16853 6103 16911 6109
rect 16853 6069 16865 6103
rect 16899 6100 16911 6103
rect 16942 6100 16948 6112
rect 16899 6072 16948 6100
rect 16899 6069 16911 6072
rect 16853 6063 16911 6069
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 17494 6100 17500 6112
rect 17455 6072 17500 6100
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6100 18107 6103
rect 19242 6100 19248 6112
rect 18095 6072 19248 6100
rect 18095 6069 18107 6072
rect 18049 6063 18107 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 20162 6100 20168 6112
rect 20123 6072 20168 6100
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 21821 6103 21879 6109
rect 21821 6069 21833 6103
rect 21867 6100 21879 6103
rect 21910 6100 21916 6112
rect 21867 6072 21916 6100
rect 21867 6069 21879 6072
rect 21821 6063 21879 6069
rect 21910 6060 21916 6072
rect 21968 6060 21974 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2866 5896 2872 5908
rect 2827 5868 2872 5896
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4212 5868 4537 5896
rect 4212 5856 4218 5868
rect 4525 5865 4537 5868
rect 4571 5896 4583 5899
rect 4890 5896 4896 5908
rect 4571 5868 4896 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 7742 5896 7748 5908
rect 7703 5868 7748 5896
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8628 5868 8677 5896
rect 8628 5856 8634 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 9490 5896 9496 5908
rect 9451 5868 9496 5896
rect 8665 5859 8723 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 11146 5896 11152 5908
rect 9723 5868 11152 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 12621 5899 12679 5905
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 13078 5896 13084 5908
rect 12667 5868 13084 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13998 5896 14004 5908
rect 13959 5868 14004 5896
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14366 5896 14372 5908
rect 14327 5868 14372 5896
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 16025 5899 16083 5905
rect 16025 5865 16037 5899
rect 16071 5896 16083 5899
rect 16206 5896 16212 5908
rect 16071 5868 16212 5896
rect 16071 5865 16083 5868
rect 16025 5859 16083 5865
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 16393 5899 16451 5905
rect 16393 5865 16405 5899
rect 16439 5896 16451 5899
rect 18046 5896 18052 5908
rect 16439 5868 18052 5896
rect 16439 5865 16451 5868
rect 16393 5859 16451 5865
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 1670 5788 1676 5840
rect 1728 5788 1734 5840
rect 1946 5788 1952 5840
rect 2004 5828 2010 5840
rect 2774 5828 2780 5840
rect 2004 5800 2780 5828
rect 2004 5788 2010 5800
rect 2774 5788 2780 5800
rect 2832 5828 2838 5840
rect 3421 5831 3479 5837
rect 3421 5828 3433 5831
rect 2832 5800 3433 5828
rect 2832 5788 2838 5800
rect 3421 5797 3433 5800
rect 3467 5797 3479 5831
rect 3421 5791 3479 5797
rect 10137 5831 10195 5837
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 10226 5828 10232 5840
rect 10183 5800 10232 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 10778 5828 10784 5840
rect 10739 5800 10784 5828
rect 10778 5788 10784 5800
rect 10836 5788 10842 5840
rect 11514 5837 11520 5840
rect 11508 5828 11520 5837
rect 11475 5800 11520 5828
rect 11508 5791 11520 5800
rect 11514 5788 11520 5791
rect 11572 5788 11578 5840
rect 12158 5788 12164 5840
rect 12216 5828 12222 5840
rect 13538 5828 13544 5840
rect 12216 5800 13544 5828
rect 12216 5788 12222 5800
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 16942 5837 16948 5840
rect 16936 5828 16948 5837
rect 16903 5800 16948 5828
rect 16936 5791 16948 5800
rect 16942 5788 16948 5791
rect 17000 5788 17006 5840
rect 17954 5788 17960 5840
rect 18012 5828 18018 5840
rect 18506 5828 18512 5840
rect 18012 5800 18512 5828
rect 18012 5788 18018 5800
rect 18506 5788 18512 5800
rect 18564 5828 18570 5840
rect 18601 5831 18659 5837
rect 18601 5828 18613 5831
rect 18564 5800 18613 5828
rect 18564 5788 18570 5800
rect 18601 5797 18613 5800
rect 18647 5797 18659 5831
rect 18601 5791 18659 5797
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 1688 5760 1716 5788
rect 1535 5732 1716 5760
rect 1756 5763 1814 5769
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 1756 5729 1768 5763
rect 1802 5760 1814 5763
rect 1964 5760 1992 5788
rect 1802 5732 1992 5760
rect 4433 5763 4491 5769
rect 1802 5729 1814 5732
rect 1756 5723 1814 5729
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 4706 5760 4712 5772
rect 4479 5732 4712 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 6328 5732 6377 5760
rect 6328 5720 6334 5732
rect 6365 5729 6377 5732
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6621 5763 6679 5769
rect 6621 5760 6633 5763
rect 6512 5732 6633 5760
rect 6512 5720 6518 5732
rect 6621 5729 6633 5732
rect 6667 5729 6679 5763
rect 6621 5723 6679 5729
rect 7006 5720 7012 5772
rect 7064 5760 7070 5772
rect 7190 5760 7196 5772
rect 7064 5732 7196 5760
rect 7064 5720 7070 5732
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10962 5720 10968 5772
rect 11020 5760 11026 5772
rect 11241 5763 11299 5769
rect 11241 5760 11253 5763
rect 11020 5732 11253 5760
rect 11020 5720 11026 5732
rect 11241 5729 11253 5732
rect 11287 5729 11299 5763
rect 14182 5760 14188 5772
rect 14143 5732 14188 5760
rect 11241 5723 11299 5729
rect 14182 5720 14188 5732
rect 14240 5760 14246 5772
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 14240 5732 14657 5760
rect 14240 5720 14246 5732
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 15381 5763 15439 5769
rect 15381 5729 15393 5763
rect 15427 5729 15439 5763
rect 15381 5723 15439 5729
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 4632 5624 4660 5655
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 10229 5695 10287 5701
rect 8720 5664 10088 5692
rect 8720 5652 8726 5664
rect 4396 5596 4660 5624
rect 9125 5627 9183 5633
rect 4396 5584 4402 5596
rect 9125 5593 9137 5627
rect 9171 5624 9183 5627
rect 9582 5624 9588 5636
rect 9171 5596 9588 5624
rect 9171 5593 9183 5596
rect 9125 5587 9183 5593
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 10060 5624 10088 5664
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 15010 5692 15016 5704
rect 14971 5664 15016 5692
rect 10229 5655 10287 5661
rect 10244 5624 10272 5655
rect 15010 5652 15016 5664
rect 15068 5692 15074 5704
rect 15396 5692 15424 5723
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 15528 5732 16681 5760
rect 15528 5720 15534 5732
rect 16669 5729 16681 5732
rect 16715 5760 16727 5763
rect 17494 5760 17500 5772
rect 16715 5732 17500 5760
rect 16715 5729 16727 5732
rect 16669 5723 16727 5729
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 19150 5760 19156 5772
rect 19111 5732 19156 5760
rect 19150 5720 19156 5732
rect 19208 5720 19214 5772
rect 20162 5720 20168 5772
rect 20220 5760 20226 5772
rect 20898 5760 20904 5772
rect 20220 5732 20904 5760
rect 20220 5720 20226 5732
rect 20898 5720 20904 5732
rect 20956 5760 20962 5772
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20956 5732 21005 5760
rect 20956 5720 20962 5732
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 15068 5664 15424 5692
rect 15068 5652 15074 5664
rect 11054 5624 11060 5636
rect 10060 5596 11060 5624
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 2924 5528 3801 5556
rect 2924 5516 2930 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 3789 5519 3847 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 5350 5556 5356 5568
rect 4212 5528 5356 5556
rect 4212 5516 4218 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5500 5528 5733 5556
rect 5500 5516 5506 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 6086 5556 6092 5568
rect 6047 5528 6092 5556
rect 5721 5519 5779 5525
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8386 5556 8392 5568
rect 8260 5528 8392 5556
rect 8260 5516 8266 5528
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 13173 5559 13231 5565
rect 13173 5556 13185 5559
rect 12492 5528 13185 5556
rect 12492 5516 12498 5528
rect 13173 5525 13185 5528
rect 13219 5525 13231 5559
rect 13173 5519 13231 5525
rect 15565 5559 15623 5565
rect 15565 5525 15577 5559
rect 15611 5556 15623 5559
rect 15838 5556 15844 5568
rect 15611 5528 15844 5556
rect 15611 5525 15623 5528
rect 15565 5519 15623 5525
rect 15838 5516 15844 5528
rect 15896 5516 15902 5568
rect 19334 5556 19340 5568
rect 19295 5528 19340 5556
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 21174 5556 21180 5568
rect 21135 5528 21180 5556
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 2222 5352 2228 5364
rect 1443 5324 2228 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3234 5352 3240 5364
rect 2915 5324 3240 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 2406 5284 2412 5296
rect 2056 5256 2412 5284
rect 2056 5225 2084 5256
rect 2406 5244 2412 5256
rect 2464 5244 2470 5296
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 2976 5225 3004 5324
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 4338 5352 4344 5364
rect 4299 5324 4344 5352
rect 4338 5312 4344 5324
rect 4396 5352 4402 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 4396 5324 5273 5352
rect 4396 5312 4402 5324
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6328 5324 6377 5352
rect 6328 5312 6334 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6822 5352 6828 5364
rect 6783 5324 6828 5352
rect 6365 5315 6423 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7800 5324 7849 5352
rect 7800 5312 7806 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10778 5352 10784 5364
rect 9815 5324 10784 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11606 5312 11612 5364
rect 11664 5352 11670 5364
rect 11882 5352 11888 5364
rect 11664 5324 11888 5352
rect 11664 5312 11670 5324
rect 11882 5312 11888 5324
rect 11940 5352 11946 5364
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 11940 5324 13185 5352
rect 11940 5312 11946 5324
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 13173 5315 13231 5321
rect 17313 5355 17371 5361
rect 17313 5321 17325 5355
rect 17359 5352 17371 5355
rect 17494 5352 17500 5364
rect 17359 5324 17500 5352
rect 17359 5321 17371 5324
rect 17313 5315 17371 5321
rect 4890 5284 4896 5296
rect 4851 5256 4896 5284
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2648 5188 2973 5216
rect 2648 5176 2654 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 7760 5216 7788 5312
rect 10042 5244 10048 5296
rect 10100 5284 10106 5296
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 10100 5256 10701 5284
rect 10100 5244 10106 5256
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 10689 5247 10747 5253
rect 7515 5188 7788 5216
rect 13188 5216 13216 5315
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 19150 5352 19156 5364
rect 19111 5324 19156 5352
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 20898 5352 20904 5364
rect 20859 5324 20904 5352
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 16206 5284 16212 5296
rect 16167 5256 16212 5284
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 20625 5287 20683 5293
rect 20625 5253 20637 5287
rect 20671 5284 20683 5287
rect 21269 5287 21327 5293
rect 21269 5284 21281 5287
rect 20671 5256 21281 5284
rect 20671 5253 20683 5256
rect 20625 5247 20683 5253
rect 21269 5253 21281 5256
rect 21315 5253 21327 5287
rect 21269 5247 21327 5253
rect 13357 5219 13415 5225
rect 13357 5216 13369 5219
rect 13188 5188 13369 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 13357 5185 13369 5188
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5216 15807 5219
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 15795 5188 16773 5216
rect 15795 5185 15807 5188
rect 15749 5179 15807 5185
rect 16761 5185 16773 5188
rect 16807 5216 16819 5219
rect 16942 5216 16948 5228
rect 16807 5188 16948 5216
rect 16807 5185 16819 5188
rect 16761 5179 16819 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 18598 5216 18604 5228
rect 18559 5188 18604 5216
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1452 5120 1777 5148
rect 1452 5108 1458 5120
rect 1765 5117 1777 5120
rect 1811 5148 1823 5151
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 1811 5120 2421 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3217 5151 3275 5157
rect 3217 5148 3229 5151
rect 3108 5120 3229 5148
rect 3108 5108 3114 5120
rect 3217 5117 3229 5120
rect 3263 5117 3275 5151
rect 3217 5111 3275 5117
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5148 7343 5151
rect 7834 5148 7840 5160
rect 7331 5120 7840 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 8662 5157 8668 5160
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5117 8447 5151
rect 8656 5148 8668 5157
rect 8623 5120 8668 5148
rect 8389 5111 8447 5117
rect 8656 5111 8668 5120
rect 6270 5040 6276 5092
rect 6328 5080 6334 5092
rect 6730 5080 6736 5092
rect 6328 5052 6736 5080
rect 6328 5040 6334 5052
rect 6730 5040 6736 5052
rect 6788 5080 6794 5092
rect 8205 5083 8263 5089
rect 8205 5080 8217 5083
rect 6788 5052 8217 5080
rect 6788 5040 6794 5052
rect 8205 5049 8217 5052
rect 8251 5080 8263 5083
rect 8404 5080 8432 5111
rect 8662 5108 8668 5111
rect 8720 5108 8726 5160
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 16577 5151 16635 5157
rect 16577 5148 16589 5151
rect 16163 5120 16589 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 16577 5117 16589 5120
rect 16623 5148 16635 5151
rect 16850 5148 16856 5160
rect 16623 5120 16856 5148
rect 16623 5117 16635 5120
rect 16577 5111 16635 5117
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 18506 5148 18512 5160
rect 18467 5120 18512 5148
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5148 20039 5151
rect 20640 5148 20668 5247
rect 21082 5148 21088 5160
rect 20027 5120 20668 5148
rect 21043 5120 21088 5148
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 21082 5108 21088 5120
rect 21140 5148 21146 5160
rect 21545 5151 21603 5157
rect 21545 5148 21557 5151
rect 21140 5120 21557 5148
rect 21140 5108 21146 5120
rect 21545 5117 21557 5120
rect 21591 5117 21603 5151
rect 21545 5111 21603 5117
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22557 5151 22615 5157
rect 22557 5148 22569 5151
rect 22152 5120 22569 5148
rect 22152 5108 22158 5120
rect 22557 5117 22569 5120
rect 22603 5117 22615 5151
rect 22557 5111 22615 5117
rect 8251 5052 8432 5080
rect 8251 5049 8263 5052
rect 8205 5043 8263 5049
rect 8404 5024 8432 5052
rect 10226 5040 10232 5092
rect 10284 5040 10290 5092
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 13624 5083 13682 5089
rect 13624 5080 13636 5083
rect 12943 5052 13636 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 13624 5049 13636 5052
rect 13670 5080 13682 5083
rect 13722 5080 13728 5092
rect 13670 5052 13728 5080
rect 13670 5049 13682 5052
rect 13624 5043 13682 5049
rect 13722 5040 13728 5052
rect 13780 5040 13786 5092
rect 16482 5040 16488 5092
rect 16540 5080 16546 5092
rect 16669 5083 16727 5089
rect 16669 5080 16681 5083
rect 16540 5052 16681 5080
rect 16540 5040 16546 5052
rect 16669 5049 16681 5052
rect 16715 5049 16727 5083
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 16669 5043 16727 5049
rect 17788 5052 18429 5080
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1820 4984 1869 5012
rect 1820 4972 1826 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 6822 5012 6828 5024
rect 5767 4984 6828 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 6822 4972 6828 4984
rect 6880 5012 6886 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6880 4984 7205 5012
rect 6880 4972 6886 4984
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7193 4975 7251 4981
rect 8386 4972 8392 5024
rect 8444 4972 8450 5024
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 10244 5012 10272 5040
rect 17788 5024 17816 5052
rect 18417 5049 18429 5052
rect 18463 5049 18475 5083
rect 18417 5043 18475 5049
rect 10321 5015 10379 5021
rect 10321 5012 10333 5015
rect 10100 4984 10333 5012
rect 10100 4972 10106 4984
rect 10321 4981 10333 4984
rect 10367 4981 10379 5015
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 10321 4975 10379 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 12158 5012 12164 5024
rect 12119 4984 12164 5012
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 14737 5015 14795 5021
rect 14737 4981 14749 5015
rect 14783 5012 14795 5015
rect 14826 5012 14832 5024
rect 14783 4984 14832 5012
rect 14783 4981 14795 4984
rect 14737 4975 14795 4981
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 15286 5012 15292 5024
rect 15247 4984 15292 5012
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 20162 5012 20168 5024
rect 20123 4984 20168 5012
rect 20162 4972 20168 4984
rect 20220 4972 20226 5024
rect 22278 5012 22284 5024
rect 22239 4984 22284 5012
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2590 4808 2596 4820
rect 2363 4780 2596 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 4062 4808 4068 4820
rect 2915 4780 4068 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 4062 4768 4068 4780
rect 4120 4808 4126 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 4120 4780 5089 4808
rect 4120 4768 4126 4780
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 5077 4771 5135 4777
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 6086 4808 6092 4820
rect 5767 4780 6092 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 6454 4808 6460 4820
rect 6415 4780 6460 4808
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 6822 4808 6828 4820
rect 6783 4780 6828 4808
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7834 4808 7840 4820
rect 7607 4780 7840 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 8938 4808 8944 4820
rect 8527 4780 8944 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 8938 4768 8944 4780
rect 8996 4808 9002 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 8996 4780 9689 4808
rect 8996 4768 9002 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 10134 4808 10140 4820
rect 10095 4780 10140 4808
rect 9677 4771 9735 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11422 4808 11428 4820
rect 11379 4780 11428 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11517 4811 11575 4817
rect 11517 4777 11529 4811
rect 11563 4808 11575 4811
rect 13538 4808 13544 4820
rect 11563 4780 13544 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 15286 4808 15292 4820
rect 15247 4780 15292 4808
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 16393 4811 16451 4817
rect 16393 4777 16405 4811
rect 16439 4808 16451 4811
rect 16482 4808 16488 4820
rect 16439 4780 16488 4808
rect 16439 4777 16451 4780
rect 16393 4771 16451 4777
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 16942 4808 16948 4820
rect 16807 4780 16948 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17310 4808 17316 4820
rect 17271 4780 17316 4808
rect 17310 4768 17316 4780
rect 17368 4768 17374 4820
rect 17954 4768 17960 4820
rect 18012 4808 18018 4820
rect 18141 4811 18199 4817
rect 18141 4808 18153 4811
rect 18012 4780 18153 4808
rect 18012 4768 18018 4780
rect 18141 4777 18153 4780
rect 18187 4808 18199 4811
rect 18598 4808 18604 4820
rect 18187 4780 18604 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 1397 4743 1455 4749
rect 1397 4709 1409 4743
rect 1443 4740 1455 4743
rect 2038 4740 2044 4752
rect 1443 4712 2044 4740
rect 1443 4709 1455 4712
rect 1397 4703 1455 4709
rect 2038 4700 2044 4712
rect 2096 4700 2102 4752
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 3421 4743 3479 4749
rect 3421 4740 3433 4743
rect 3108 4712 3433 4740
rect 3108 4700 3114 4712
rect 3421 4709 3433 4712
rect 3467 4709 3479 4743
rect 3421 4703 3479 4709
rect 8110 4700 8116 4752
rect 8168 4740 8174 4752
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 8168 4712 8401 4740
rect 8168 4700 8174 4712
rect 8389 4709 8401 4712
rect 8435 4740 8447 4743
rect 8570 4740 8576 4752
rect 8435 4712 8576 4740
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 8662 4700 8668 4752
rect 8720 4740 8726 4752
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 8720 4712 9045 4740
rect 8720 4700 8726 4712
rect 9033 4709 9045 4712
rect 9079 4709 9091 4743
rect 9033 4703 9091 4709
rect 9582 4700 9588 4752
rect 9640 4740 9646 4752
rect 10042 4740 10048 4752
rect 9640 4712 10048 4740
rect 9640 4700 9646 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 2406 4632 2412 4684
rect 2464 4632 2470 4684
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 5626 4672 5632 4684
rect 2823 4644 3464 4672
rect 5587 4644 5632 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 2424 4604 2452 4632
rect 3436 4616 3464 4644
rect 5626 4632 5632 4644
rect 5684 4672 5690 4684
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 5684 4644 7849 4672
rect 5684 4632 5690 4644
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 7837 4635 7895 4641
rect 9493 4675 9551 4681
rect 9493 4641 9505 4675
rect 9539 4672 9551 4675
rect 10152 4672 10180 4768
rect 15105 4743 15163 4749
rect 15105 4709 15117 4743
rect 15151 4740 15163 4743
rect 15562 4740 15568 4752
rect 15151 4712 15568 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 15562 4700 15568 4712
rect 15620 4740 15626 4752
rect 15620 4712 15884 4740
rect 15620 4700 15626 4712
rect 9539 4644 10180 4672
rect 9539 4641 9551 4644
rect 9493 4635 9551 4641
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11885 4675 11943 4681
rect 11885 4672 11897 4675
rect 11112 4644 11897 4672
rect 11112 4632 11118 4644
rect 11885 4641 11897 4644
rect 11931 4672 11943 4675
rect 12158 4672 12164 4684
rect 11931 4644 12164 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 13446 4672 13452 4684
rect 13407 4644 13452 4672
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 14642 4632 14648 4684
rect 14700 4672 14706 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 14700 4644 15669 4672
rect 14700 4632 14706 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 3050 4604 3056 4616
rect 2004 4576 2912 4604
rect 3011 4576 3056 4604
rect 2004 4564 2010 4576
rect 2406 4536 2412 4548
rect 2367 4508 2412 4536
rect 2406 4496 2412 4508
rect 2464 4496 2470 4548
rect 2884 4536 2912 4576
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 3476 4576 4261 4604
rect 3476 4564 3482 4576
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 6178 4604 6184 4616
rect 5951 4576 6184 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 8478 4564 8484 4616
rect 8536 4604 8542 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8536 4576 8585 4604
rect 8536 4564 8542 4576
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 10226 4604 10232 4616
rect 10187 4576 10232 4604
rect 8573 4567 8631 4573
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 10962 4604 10968 4616
rect 10875 4576 10968 4604
rect 10962 4564 10968 4576
rect 11020 4604 11026 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11020 4576 11989 4604
rect 11020 4564 11026 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 12066 4564 12072 4616
rect 12124 4604 12130 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 12124 4576 12541 4604
rect 12124 4564 12130 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 13722 4604 13728 4616
rect 13683 4576 13728 4604
rect 12529 4567 12587 4573
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 15746 4604 15752 4616
rect 15707 4576 15752 4604
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 15856 4613 15884 4712
rect 16114 4672 16120 4684
rect 15948 4644 16120 4672
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 3786 4536 3792 4548
rect 2884 4508 3792 4536
rect 3786 4496 3792 4508
rect 3844 4536 3850 4548
rect 4338 4536 4344 4548
rect 3844 4508 4344 4536
rect 3844 4496 3850 4508
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 13078 4536 13084 4548
rect 13039 4508 13084 4536
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 13354 4496 13360 4548
rect 13412 4536 13418 4548
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 13412 4508 14473 4536
rect 13412 4496 13418 4508
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 15764 4536 15792 4564
rect 15948 4536 15976 4644
rect 16114 4632 16120 4644
rect 16172 4672 16178 4684
rect 17218 4672 17224 4684
rect 16172 4644 17224 4672
rect 16172 4632 16178 4644
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17954 4632 17960 4684
rect 18012 4672 18018 4684
rect 18417 4675 18475 4681
rect 18417 4672 18429 4675
rect 18012 4644 18429 4672
rect 18012 4632 18018 4644
rect 18417 4641 18429 4644
rect 18463 4672 18475 4675
rect 18598 4672 18604 4684
rect 18463 4644 18604 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 19334 4632 19340 4684
rect 19392 4672 19398 4684
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 19392 4644 19533 4672
rect 19392 4632 19398 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 19521 4635 19579 4641
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 21266 4632 21272 4684
rect 21324 4672 21330 4684
rect 21913 4675 21971 4681
rect 21913 4672 21925 4675
rect 21324 4644 21925 4672
rect 21324 4632 21330 4644
rect 21913 4641 21925 4644
rect 21959 4672 21971 4675
rect 22002 4672 22008 4684
rect 21959 4644 22008 4672
rect 21959 4641 21971 4644
rect 21913 4635 21971 4641
rect 22002 4632 22008 4644
rect 22060 4632 22066 4684
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4604 17555 4607
rect 17678 4604 17684 4616
rect 17543 4576 17684 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 16850 4536 16856 4548
rect 15764 4508 15976 4536
rect 16811 4508 16856 4536
rect 14461 4499 14519 4505
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 1762 4428 1768 4480
rect 1820 4468 1826 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1820 4440 1869 4468
rect 1820 4428 1826 4440
rect 1857 4437 1869 4440
rect 1903 4437 1915 4471
rect 4706 4468 4712 4480
rect 4667 4440 4712 4468
rect 1857 4431 1915 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 8018 4468 8024 4480
rect 7979 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 12894 4468 12900 4480
rect 12855 4440 12900 4468
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 14182 4468 14188 4480
rect 14143 4440 14188 4468
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 19518 4468 19524 4480
rect 18647 4440 19524 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 20806 4468 20812 4480
rect 19751 4440 20812 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 21082 4468 21088 4480
rect 21043 4440 21088 4468
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22152 4440 22197 4468
rect 22152 4428 22158 4440
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1762 4264 1768 4276
rect 1412 4236 1768 4264
rect 1412 4196 1440 4236
rect 1762 4224 1768 4236
rect 1820 4224 1826 4276
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3418 4264 3424 4276
rect 2832 4236 2877 4264
rect 3379 4236 3424 4264
rect 2832 4224 2838 4236
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 4338 4264 4344 4276
rect 4299 4236 4344 4264
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4893 4267 4951 4273
rect 4893 4233 4905 4267
rect 4939 4264 4951 4267
rect 6086 4264 6092 4276
rect 4939 4236 6092 4264
rect 4939 4233 4951 4236
rect 4893 4227 4951 4233
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8444 4236 8493 4264
rect 8444 4224 8450 4236
rect 8481 4233 8493 4236
rect 8527 4264 8539 4267
rect 8573 4267 8631 4273
rect 8573 4264 8585 4267
rect 8527 4236 8585 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 8573 4233 8585 4236
rect 8619 4233 8631 4267
rect 8573 4227 8631 4233
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 11974 4264 11980 4276
rect 11931 4236 11980 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 11974 4224 11980 4236
rect 12032 4264 12038 4276
rect 12710 4264 12716 4276
rect 12032 4236 12716 4264
rect 12032 4224 12038 4236
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13817 4267 13875 4273
rect 13817 4264 13829 4267
rect 13596 4236 13829 4264
rect 13596 4224 13602 4236
rect 13817 4233 13829 4236
rect 13863 4233 13875 4267
rect 15746 4264 15752 4276
rect 13817 4227 13875 4233
rect 15028 4236 15752 4264
rect 1320 4168 1440 4196
rect 290 4088 296 4140
rect 348 4128 354 4140
rect 1320 4128 1348 4168
rect 3050 4156 3056 4208
rect 3108 4196 3114 4208
rect 3697 4199 3755 4205
rect 3697 4196 3709 4199
rect 3108 4168 3709 4196
rect 3108 4156 3114 4168
rect 3697 4165 3709 4168
rect 3743 4196 3755 4199
rect 3970 4196 3976 4208
rect 3743 4168 3976 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 11241 4199 11299 4205
rect 6840 4168 8248 4196
rect 348 4100 1348 4128
rect 348 4088 354 4100
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 3660 4100 4813 4128
rect 3660 4088 3666 4100
rect 4801 4097 4813 4100
rect 4847 4128 4859 4131
rect 5166 4128 5172 4140
rect 4847 4100 5172 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 5166 4088 5172 4100
rect 5224 4128 5230 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5224 4100 5457 4128
rect 5224 4088 5230 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6840 4128 6868 4168
rect 7760 4137 7788 4168
rect 6687 4100 6868 4128
rect 7745 4131 7803 4137
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 8220 4128 8248 4168
rect 11241 4165 11253 4199
rect 11287 4196 11299 4199
rect 12066 4196 12072 4208
rect 11287 4168 12072 4196
rect 11287 4165 11299 4168
rect 11241 4159 11299 4165
rect 12066 4156 12072 4168
rect 12124 4196 12130 4208
rect 12986 4196 12992 4208
rect 12124 4168 12992 4196
rect 12124 4156 12130 4168
rect 12986 4156 12992 4168
rect 13044 4196 13050 4208
rect 13044 4168 13124 4196
rect 13044 4156 13050 4168
rect 12894 4128 12900 4140
rect 8220 4100 8892 4128
rect 12855 4100 12900 4128
rect 7745 4091 7803 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1486 4060 1492 4072
rect 1443 4032 1492 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1486 4020 1492 4032
rect 1544 4060 1550 4072
rect 2590 4060 2596 4072
rect 1544 4032 2596 4060
rect 1544 4020 1550 4032
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8202 4060 8208 4072
rect 7699 4032 8208 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8527 4032 8769 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8864 4060 8892 4100
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13096 4137 13124 4168
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 14148 4100 14473 4128
rect 14148 4088 14154 4100
rect 14461 4097 14473 4100
rect 14507 4128 14519 4131
rect 14642 4128 14648 4140
rect 14507 4100 14648 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 15028 4128 15056 4236
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 17037 4267 17095 4273
rect 17037 4233 17049 4267
rect 17083 4264 17095 4267
rect 17310 4264 17316 4276
rect 17083 4236 17316 4264
rect 17083 4233 17095 4236
rect 17037 4227 17095 4233
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 18598 4264 18604 4276
rect 18559 4236 18604 4264
rect 18598 4224 18604 4236
rect 18656 4224 18662 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 20073 4267 20131 4273
rect 20073 4264 20085 4267
rect 19392 4236 20085 4264
rect 19392 4224 19398 4236
rect 20073 4233 20085 4236
rect 20119 4233 20131 4267
rect 20073 4227 20131 4233
rect 21082 4224 21088 4276
rect 21140 4264 21146 4276
rect 21177 4267 21235 4273
rect 21177 4264 21189 4267
rect 21140 4236 21189 4264
rect 21140 4224 21146 4236
rect 21177 4233 21189 4236
rect 21223 4233 21235 4267
rect 22002 4264 22008 4276
rect 21963 4236 22008 4264
rect 21177 4227 21235 4233
rect 14844 4100 15056 4128
rect 9030 4069 9036 4072
rect 9013 4063 9036 4069
rect 9013 4060 9025 4063
rect 8864 4032 9025 4060
rect 8757 4023 8815 4029
rect 9013 4029 9025 4032
rect 9088 4060 9094 4072
rect 10226 4060 10232 4072
rect 9088 4032 10232 4060
rect 9013 4023 9036 4029
rect 9030 4020 9036 4023
rect 9088 4020 9094 4032
rect 10226 4020 10232 4032
rect 10284 4060 10290 4072
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10284 4032 10701 4060
rect 10284 4020 10290 4032
rect 10689 4029 10701 4032
rect 10735 4029 10747 4063
rect 11330 4060 11336 4072
rect 11243 4032 11336 4060
rect 10689 4023 10747 4029
rect 11330 4020 11336 4032
rect 11388 4060 11394 4072
rect 13354 4060 13360 4072
rect 11388 4032 13360 4060
rect 11388 4020 11394 4032
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13541 4063 13599 4069
rect 13541 4029 13553 4063
rect 13587 4060 13599 4063
rect 13814 4060 13820 4072
rect 13587 4032 13820 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 13998 4060 14004 4072
rect 13959 4032 14004 4060
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14844 4069 14872 4100
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 17276 4100 17325 4128
rect 17276 4088 17282 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14424 4032 14841 4060
rect 14424 4020 14430 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 15010 4060 15016 4072
rect 14971 4032 15016 4060
rect 14829 4023 14887 4029
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15280 4063 15338 4069
rect 15280 4029 15292 4063
rect 15326 4060 15338 4063
rect 15562 4060 15568 4072
rect 15326 4032 15568 4060
rect 15326 4029 15338 4032
rect 15280 4023 15338 4029
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18138 4060 18144 4072
rect 18095 4032 18144 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18138 4020 18144 4032
rect 18196 4060 18202 4072
rect 18969 4063 19027 4069
rect 18969 4060 18981 4063
rect 18196 4032 18981 4060
rect 18196 4020 18202 4032
rect 18969 4029 18981 4032
rect 19015 4029 19027 4063
rect 18969 4023 19027 4029
rect 19153 4063 19211 4069
rect 19153 4029 19165 4063
rect 19199 4060 19211 4063
rect 20257 4063 20315 4069
rect 19199 4032 19840 4060
rect 19199 4029 19211 4032
rect 19153 4023 19211 4029
rect 19812 4004 19840 4032
rect 20257 4029 20269 4063
rect 20303 4029 20315 4063
rect 21192 4060 21220 4227
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 21361 4063 21419 4069
rect 21361 4060 21373 4063
rect 21192 4032 21373 4060
rect 20257 4023 20315 4029
rect 21361 4029 21373 4032
rect 21407 4029 21419 4063
rect 22462 4060 22468 4072
rect 22423 4032 22468 4060
rect 21361 4023 21419 4029
rect 1664 3995 1722 4001
rect 1664 3961 1676 3995
rect 1710 3992 1722 3995
rect 2866 3992 2872 4004
rect 1710 3964 2872 3992
rect 1710 3961 1722 3964
rect 1664 3955 1722 3961
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 5261 3995 5319 4001
rect 5261 3961 5273 3995
rect 5307 3992 5319 3995
rect 5442 3992 5448 4004
rect 5307 3964 5448 3992
rect 5307 3961 5319 3964
rect 5261 3955 5319 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6178 3992 6184 4004
rect 6043 3964 6184 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6178 3952 6184 3964
rect 6236 3992 6242 4004
rect 6914 3992 6920 4004
rect 6236 3964 6920 3992
rect 6236 3952 6242 3964
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7561 3995 7619 4001
rect 7561 3992 7573 3995
rect 7024 3964 7573 3992
rect 7024 3936 7052 3964
rect 7561 3961 7573 3964
rect 7607 3961 7619 3995
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 7561 3955 7619 3961
rect 8496 3964 10180 3992
rect 8496 3936 8524 3964
rect 3878 3924 3884 3936
rect 3839 3896 3884 3924
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 5534 3924 5540 3936
rect 5399 3896 5540 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 8110 3924 8116 3936
rect 7239 3896 8116 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8294 3924 8300 3936
rect 8255 3896 8300 3924
rect 8294 3884 8300 3896
rect 8352 3924 8358 3936
rect 8478 3924 8484 3936
rect 8352 3896 8484 3924
rect 8352 3884 8358 3896
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 10152 3933 10180 3964
rect 12176 3964 12817 3992
rect 12176 3936 12204 3964
rect 12805 3961 12817 3964
rect 12851 3961 12863 3995
rect 14642 3992 14648 4004
rect 12805 3955 12863 3961
rect 14200 3964 14648 3992
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3893 10195 3927
rect 11514 3924 11520 3936
rect 11475 3896 11520 3924
rect 10137 3887 10195 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 12158 3924 12164 3936
rect 12119 3896 12164 3924
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 13446 3924 13452 3936
rect 12483 3896 13452 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 14200 3933 14228 3964
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 19794 3992 19800 4004
rect 19755 3964 19800 3992
rect 19794 3952 19800 3964
rect 19852 3952 19858 4004
rect 20272 3992 20300 4023
rect 22462 4020 22468 4032
rect 22520 4060 22526 4072
rect 22925 4063 22983 4069
rect 22925 4060 22937 4063
rect 22520 4032 22937 4060
rect 22520 4020 22526 4032
rect 22925 4029 22937 4032
rect 22971 4029 22983 4063
rect 22925 4023 22983 4029
rect 20901 3995 20959 4001
rect 20901 3992 20913 3995
rect 20272 3964 20913 3992
rect 20901 3961 20913 3964
rect 20947 3992 20959 3995
rect 22278 3992 22284 4004
rect 20947 3964 22284 3992
rect 20947 3961 20959 3964
rect 20901 3955 20959 3961
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 14185 3927 14243 3933
rect 14185 3893 14197 3927
rect 14231 3893 14243 3927
rect 16390 3924 16396 3936
rect 16351 3896 16396 3924
rect 14185 3887 14243 3893
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 17678 3924 17684 3936
rect 17639 3896 17684 3924
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 18012 3896 18245 3924
rect 18012 3884 18018 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 19337 3927 19395 3933
rect 19337 3893 19349 3927
rect 19383 3924 19395 3927
rect 20254 3924 20260 3936
rect 19383 3896 20260 3924
rect 19383 3893 19395 3896
rect 19337 3887 19395 3893
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20441 3927 20499 3933
rect 20441 3893 20453 3927
rect 20487 3924 20499 3927
rect 21358 3924 21364 3936
rect 20487 3896 21364 3924
rect 20487 3893 20499 3896
rect 20441 3887 20499 3893
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 21542 3924 21548 3936
rect 21503 3896 21548 3924
rect 21542 3884 21548 3896
rect 21600 3884 21606 3936
rect 22646 3924 22652 3936
rect 22607 3896 22652 3924
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2866 3720 2872 3732
rect 2827 3692 2872 3720
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 3476 3692 3525 3720
rect 3476 3680 3482 3692
rect 3513 3689 3525 3692
rect 3559 3720 3571 3723
rect 3602 3720 3608 3732
rect 3559 3692 3608 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 4246 3720 4252 3732
rect 4207 3692 4252 3720
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 4982 3720 4988 3732
rect 4943 3692 4988 3720
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5261 3723 5319 3729
rect 5261 3689 5273 3723
rect 5307 3720 5319 3723
rect 5442 3720 5448 3732
rect 5307 3692 5448 3720
rect 5307 3689 5319 3692
rect 5261 3683 5319 3689
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6641 3723 6699 3729
rect 6641 3720 6653 3723
rect 5592 3692 6653 3720
rect 5592 3680 5598 3692
rect 6641 3689 6653 3692
rect 6687 3689 6699 3723
rect 6641 3683 6699 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 9088 3692 9137 3720
rect 9088 3680 9094 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3720 10103 3723
rect 10778 3720 10784 3732
rect 10091 3692 10784 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11146 3720 11152 3732
rect 11107 3692 11152 3720
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 13909 3723 13967 3729
rect 13909 3720 13921 3723
rect 13504 3692 13921 3720
rect 13504 3680 13510 3692
rect 13909 3689 13921 3692
rect 13955 3689 13967 3723
rect 13909 3683 13967 3689
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15749 3723 15807 3729
rect 15749 3720 15761 3723
rect 15344 3692 15761 3720
rect 15344 3680 15350 3692
rect 15749 3689 15761 3692
rect 15795 3689 15807 3723
rect 18230 3720 18236 3732
rect 18191 3692 18236 3720
rect 15749 3683 15807 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 19242 3680 19248 3732
rect 19300 3720 19306 3732
rect 19889 3723 19947 3729
rect 19889 3720 19901 3723
rect 19300 3692 19901 3720
rect 19300 3680 19306 3692
rect 19889 3689 19901 3692
rect 19935 3720 19947 3723
rect 20162 3720 20168 3732
rect 19935 3692 20168 3720
rect 19935 3689 19947 3692
rect 19889 3683 19947 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20990 3680 20996 3732
rect 21048 3720 21054 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 21048 3692 21373 3720
rect 21048 3680 21054 3692
rect 21361 3689 21373 3692
rect 21407 3689 21419 3723
rect 21361 3683 21419 3689
rect 1756 3655 1814 3661
rect 1756 3621 1768 3655
rect 1802 3652 1814 3655
rect 1946 3652 1952 3664
rect 1802 3624 1952 3652
rect 1802 3621 1814 3624
rect 1756 3615 1814 3621
rect 1946 3612 1952 3624
rect 2004 3612 2010 3664
rect 5718 3652 5724 3664
rect 5679 3624 5724 3652
rect 5718 3612 5724 3624
rect 5776 3652 5782 3664
rect 6178 3652 6184 3664
rect 5776 3624 6184 3652
rect 5776 3612 5782 3624
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 7006 3612 7012 3664
rect 7064 3661 7070 3664
rect 7064 3655 7128 3661
rect 7064 3621 7082 3655
rect 7116 3621 7128 3655
rect 7064 3615 7128 3621
rect 7064 3612 7070 3615
rect 9674 3612 9680 3664
rect 9732 3652 9738 3664
rect 10505 3655 10563 3661
rect 10505 3652 10517 3655
rect 9732 3624 10517 3652
rect 9732 3612 9738 3624
rect 10505 3621 10517 3624
rect 10551 3621 10563 3655
rect 11514 3652 11520 3664
rect 11427 3624 11520 3652
rect 10505 3615 10563 3621
rect 11514 3612 11520 3624
rect 11572 3652 11578 3664
rect 11876 3655 11934 3661
rect 11876 3652 11888 3655
rect 11572 3624 11888 3652
rect 11572 3612 11578 3624
rect 11876 3621 11888 3624
rect 11922 3652 11934 3655
rect 11974 3652 11980 3664
rect 11922 3624 11980 3652
rect 11922 3621 11934 3624
rect 11876 3615 11934 3621
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 13004 3652 13032 3680
rect 13541 3655 13599 3661
rect 13541 3652 13553 3655
rect 13004 3624 13553 3652
rect 13541 3621 13553 3624
rect 13587 3621 13599 3655
rect 13541 3615 13599 3621
rect 14737 3655 14795 3661
rect 14737 3621 14749 3655
rect 14783 3652 14795 3655
rect 15562 3652 15568 3664
rect 14783 3624 15568 3652
rect 14783 3621 14795 3624
rect 14737 3615 14795 3621
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 20898 3652 20904 3664
rect 20859 3624 20904 3652
rect 20898 3612 20904 3624
rect 20956 3612 20962 3664
rect 1486 3584 1492 3596
rect 1447 3556 1492 3584
rect 1486 3544 1492 3556
rect 1544 3544 1550 3596
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 6086 3584 6092 3596
rect 5675 3556 6092 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6788 3556 6837 3584
rect 6788 3544 6794 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 10410 3584 10416 3596
rect 10371 3556 10416 3584
rect 6825 3547 6883 3553
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 11606 3584 11612 3596
rect 11567 3556 11612 3584
rect 11606 3544 11612 3556
rect 11664 3584 11670 3596
rect 14093 3587 14151 3593
rect 11664 3556 12747 3584
rect 11664 3544 11670 3556
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 5951 3488 6408 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6380 3392 6408 3488
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9640 3488 9965 3516
rect 9640 3476 9646 3488
rect 9953 3485 9965 3488
rect 9999 3516 10011 3519
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 9999 3488 10701 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10689 3485 10701 3488
rect 10735 3516 10747 3519
rect 11514 3516 11520 3528
rect 10735 3488 11520 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 12719 3516 12747 3556
rect 14093 3553 14105 3587
rect 14139 3584 14151 3587
rect 14182 3584 14188 3596
rect 14139 3556 14188 3584
rect 14139 3553 14151 3556
rect 14093 3547 14151 3553
rect 14182 3544 14188 3556
rect 14240 3584 14246 3596
rect 15470 3584 15476 3596
rect 14240 3556 15476 3584
rect 14240 3544 14246 3556
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 15654 3584 15660 3596
rect 15615 3556 15660 3584
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 16758 3544 16764 3596
rect 16816 3584 16822 3596
rect 17109 3587 17167 3593
rect 17109 3584 17121 3587
rect 16816 3556 17121 3584
rect 16816 3544 16822 3556
rect 17109 3553 17121 3556
rect 17155 3553 17167 3587
rect 17109 3547 17167 3553
rect 19337 3587 19395 3593
rect 19337 3553 19349 3587
rect 19383 3584 19395 3587
rect 20622 3584 20628 3596
rect 19383 3556 20628 3584
rect 19383 3553 19395 3556
rect 19337 3547 19395 3553
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 23290 3584 23296 3596
rect 23251 3556 23296 3584
rect 23290 3544 23296 3556
rect 23348 3544 23354 3596
rect 15010 3516 15016 3528
rect 12719 3488 15016 3516
rect 15010 3476 15016 3488
rect 15068 3516 15074 3528
rect 15378 3516 15384 3528
rect 15068 3488 15384 3516
rect 15068 3476 15074 3488
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15838 3516 15844 3528
rect 15799 3488 15844 3516
rect 15838 3476 15844 3488
rect 15896 3516 15902 3528
rect 16301 3519 16359 3525
rect 16301 3516 16313 3519
rect 15896 3488 16313 3516
rect 15896 3476 15902 3488
rect 16301 3485 16313 3488
rect 16347 3516 16359 3519
rect 16390 3516 16396 3528
rect 16347 3488 16396 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 8205 3451 8263 3457
rect 8205 3417 8217 3451
rect 8251 3448 8263 3451
rect 8849 3451 8907 3457
rect 8849 3448 8861 3451
rect 8251 3420 8861 3448
rect 8251 3417 8263 3420
rect 8205 3411 8263 3417
rect 8849 3417 8861 3420
rect 8895 3448 8907 3451
rect 8938 3448 8944 3460
rect 8895 3420 8944 3448
rect 8895 3417 8907 3420
rect 8849 3411 8907 3417
rect 8938 3408 8944 3420
rect 8996 3408 9002 3460
rect 15396 3448 15424 3476
rect 16868 3448 16896 3479
rect 15396 3420 16896 3448
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3752 3352 3801 3380
rect 3752 3340 3758 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 6362 3380 6368 3392
rect 6323 3352 6368 3380
rect 3789 3343 3847 3349
rect 6362 3340 6368 3352
rect 6420 3340 6426 3392
rect 14274 3380 14280 3392
rect 14235 3352 14280 3380
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 15286 3380 15292 3392
rect 15247 3352 15292 3380
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 16758 3380 16764 3392
rect 16719 3352 16764 3380
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 16868 3380 16896 3420
rect 17218 3380 17224 3392
rect 16868 3352 17224 3380
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 18564 3352 18797 3380
rect 18564 3340 18570 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 19058 3340 19064 3392
rect 19116 3380 19122 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 19116 3352 19533 3380
rect 19116 3340 19122 3352
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 23474 3380 23480 3392
rect 23435 3352 23480 3380
rect 19521 3343 19579 3349
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1544 3148 1593 3176
rect 1544 3136 1550 3148
rect 1581 3145 1593 3148
rect 1627 3176 1639 3179
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1627 3148 1961 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 1949 3145 1961 3148
rect 1995 3176 2007 3179
rect 2317 3179 2375 3185
rect 2317 3176 2329 3179
rect 1995 3148 2329 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2317 3145 2329 3148
rect 2363 3145 2375 3179
rect 2317 3139 2375 3145
rect 2332 3040 2360 3139
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 3844 3148 3893 3176
rect 3844 3136 3850 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 4890 3176 4896 3188
rect 4851 3148 4896 3176
rect 3881 3139 3939 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5534 3176 5540 3188
rect 5031 3148 5540 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6089 3179 6147 3185
rect 6089 3145 6101 3179
rect 6135 3176 6147 3179
rect 6178 3176 6184 3188
rect 6135 3148 6184 3176
rect 6135 3145 6147 3148
rect 6089 3139 6147 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9677 3179 9735 3185
rect 9677 3176 9689 3179
rect 9088 3148 9689 3176
rect 9088 3136 9094 3148
rect 9677 3145 9689 3148
rect 9723 3145 9735 3179
rect 9677 3139 9735 3145
rect 10781 3179 10839 3185
rect 10781 3145 10793 3179
rect 10827 3176 10839 3179
rect 10962 3176 10968 3188
rect 10827 3148 10968 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 11664 3148 12173 3176
rect 11664 3136 11670 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 15013 3179 15071 3185
rect 15013 3145 15025 3179
rect 15059 3176 15071 3179
rect 15654 3176 15660 3188
rect 15059 3148 15660 3176
rect 15059 3145 15071 3148
rect 15013 3139 15071 3145
rect 2406 3040 2412 3052
rect 2319 3012 2412 3040
rect 2406 3000 2412 3012
rect 2464 3040 2470 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2464 3012 2513 3040
rect 2464 3000 2470 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 4908 3040 4936 3136
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 7009 3111 7067 3117
rect 7009 3108 7021 3111
rect 6788 3080 7021 3108
rect 6788 3068 6794 3080
rect 7009 3077 7021 3080
rect 7055 3108 7067 3111
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 7055 3080 8217 3108
rect 7055 3077 7067 3080
rect 7009 3071 7067 3077
rect 8205 3077 8217 3080
rect 8251 3108 8263 3111
rect 8251 3080 8340 3108
rect 8251 3077 8263 3080
rect 8205 3071 8263 3077
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 4908 3012 5457 3040
rect 2501 3003 2559 3009
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 6362 3040 6368 3052
rect 5675 3012 6368 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 8110 3040 8116 3052
rect 7331 3012 8116 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8312 3049 8340 3080
rect 10410 3068 10416 3120
rect 10468 3108 10474 3120
rect 11793 3111 11851 3117
rect 11793 3108 11805 3111
rect 10468 3080 11805 3108
rect 10468 3068 10474 3080
rect 11793 3077 11805 3080
rect 11839 3077 11851 3111
rect 11793 3071 11851 3077
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 9732 3012 10241 3040
rect 9732 3000 9738 3012
rect 10229 3009 10241 3012
rect 10275 3040 10287 3043
rect 10778 3040 10784 3052
rect 10275 3012 10784 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11241 3043 11299 3049
rect 11241 3040 11253 3043
rect 11204 3012 11253 3040
rect 11204 3000 11210 3012
rect 11241 3009 11253 3012
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 11425 3043 11483 3049
rect 11425 3009 11437 3043
rect 11471 3040 11483 3043
rect 11514 3040 11520 3052
rect 11471 3012 11520 3040
rect 11471 3009 11483 3012
rect 11425 3003 11483 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 12066 3000 12072 3052
rect 12124 3040 12130 3052
rect 12176 3040 12204 3139
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16816 3148 16865 3176
rect 16816 3136 16822 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17276 3148 17417 3176
rect 17276 3136 17282 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19484 3148 19625 3176
rect 19484 3136 19490 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 20622 3176 20628 3188
rect 20583 3148 20628 3176
rect 19613 3139 19671 3145
rect 20622 3136 20628 3148
rect 20680 3176 20686 3188
rect 22646 3176 22652 3188
rect 20680 3148 22652 3176
rect 20680 3136 20686 3148
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 15378 3108 15384 3120
rect 15339 3080 15384 3108
rect 15378 3068 15384 3080
rect 15436 3108 15442 3120
rect 15436 3080 15516 3108
rect 15436 3068 15442 3080
rect 15488 3049 15516 3080
rect 20714 3068 20720 3120
rect 20772 3108 20778 3120
rect 21361 3111 21419 3117
rect 21361 3108 21373 3111
rect 20772 3080 21373 3108
rect 20772 3068 20778 3080
rect 21361 3077 21373 3080
rect 21407 3077 21419 3111
rect 23290 3108 23296 3120
rect 23251 3080 23296 3108
rect 21361 3071 21419 3077
rect 23290 3068 23296 3080
rect 23348 3068 23354 3120
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12124 3012 12449 3040
rect 12124 3000 12130 3012
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 18288 3012 18613 3040
rect 18288 3000 18294 3012
rect 18601 3009 18613 3012
rect 18647 3040 18659 3043
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 18647 3012 19073 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 19061 3009 19073 3012
rect 19107 3009 19119 3043
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 19061 3003 19119 3009
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 2768 2975 2826 2981
rect 2768 2941 2780 2975
rect 2814 2972 2826 2975
rect 3694 2972 3700 2984
rect 2814 2944 3700 2972
rect 2814 2941 2826 2944
rect 2768 2935 2826 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4525 2975 4583 2981
rect 4525 2972 4537 2975
rect 4028 2944 4537 2972
rect 4028 2932 4034 2944
rect 4525 2941 4537 2944
rect 4571 2972 4583 2975
rect 6086 2972 6092 2984
rect 4571 2944 6092 2972
rect 4571 2941 4583 2944
rect 4525 2935 4583 2941
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 7006 2972 7012 2984
rect 6687 2944 7012 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 8202 2972 8208 2984
rect 7064 2944 8208 2972
rect 7064 2932 7070 2944
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8564 2975 8622 2981
rect 8564 2941 8576 2975
rect 8610 2972 8622 2975
rect 8938 2972 8944 2984
rect 8610 2944 8944 2972
rect 8610 2941 8622 2944
rect 8564 2935 8622 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 12704 2975 12762 2981
rect 12704 2941 12716 2975
rect 12750 2972 12762 2975
rect 12986 2972 12992 2984
rect 12750 2944 12992 2972
rect 12750 2941 12762 2944
rect 12704 2935 12762 2941
rect 12986 2932 12992 2944
rect 13044 2932 13050 2984
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 20070 2972 20076 2984
rect 19392 2944 20076 2972
rect 19392 2932 19398 2944
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 21082 2932 21088 2984
rect 21140 2972 21146 2984
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 21140 2944 21189 2972
rect 21140 2932 21146 2944
rect 21177 2941 21189 2944
rect 21223 2972 21235 2975
rect 21637 2975 21695 2981
rect 21637 2972 21649 2975
rect 21223 2944 21649 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 21637 2941 21649 2944
rect 21683 2941 21695 2975
rect 22186 2972 22192 2984
rect 22147 2944 22192 2972
rect 21637 2935 21695 2941
rect 22186 2932 22192 2944
rect 22244 2972 22250 2984
rect 22649 2975 22707 2981
rect 22649 2972 22661 2975
rect 22244 2944 22661 2972
rect 22244 2932 22250 2944
rect 22649 2941 22661 2944
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 24397 2975 24455 2981
rect 24397 2972 24409 2975
rect 23532 2944 24409 2972
rect 23532 2932 23538 2944
rect 24397 2941 24409 2944
rect 24443 2972 24455 2975
rect 24949 2975 25007 2981
rect 24949 2972 24961 2975
rect 24443 2944 24961 2972
rect 24443 2941 24455 2944
rect 24397 2935 24455 2941
rect 24949 2941 24961 2944
rect 24995 2941 25007 2975
rect 24949 2935 25007 2941
rect 4982 2864 4988 2916
rect 5040 2904 5046 2916
rect 5353 2907 5411 2913
rect 5353 2904 5365 2907
rect 5040 2876 5365 2904
rect 5040 2864 5046 2876
rect 5353 2873 5365 2876
rect 5399 2873 5411 2907
rect 5353 2867 5411 2873
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 15718 2907 15776 2913
rect 15718 2904 15730 2907
rect 14691 2876 15730 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15718 2873 15730 2876
rect 15764 2904 15776 2907
rect 15838 2904 15844 2916
rect 15764 2876 15844 2904
rect 15764 2873 15776 2876
rect 15718 2867 15776 2873
rect 15838 2864 15844 2876
rect 15896 2864 15902 2916
rect 17865 2907 17923 2913
rect 17865 2873 17877 2907
rect 17911 2904 17923 2907
rect 18414 2904 18420 2916
rect 17911 2876 18420 2904
rect 17911 2873 17923 2876
rect 17865 2867 17923 2873
rect 18414 2864 18420 2876
rect 18472 2864 18478 2916
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 19521 2907 19579 2913
rect 19521 2904 19533 2907
rect 19484 2876 19533 2904
rect 19484 2864 19490 2876
rect 19521 2873 19533 2876
rect 19567 2904 19579 2907
rect 19981 2907 20039 2913
rect 19981 2904 19993 2907
rect 19567 2876 19993 2904
rect 19567 2873 19579 2876
rect 19521 2867 19579 2873
rect 19981 2873 19993 2876
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 7742 2836 7748 2848
rect 7703 2808 7748 2836
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 10689 2839 10747 2845
rect 10689 2836 10701 2839
rect 9824 2808 10701 2836
rect 9824 2796 9830 2808
rect 10689 2805 10701 2808
rect 10735 2836 10747 2839
rect 11146 2836 11152 2848
rect 10735 2808 11152 2836
rect 10735 2805 10747 2808
rect 10689 2799 10747 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 13814 2836 13820 2848
rect 13775 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 18049 2839 18107 2845
rect 18049 2805 18061 2839
rect 18095 2836 18107 2839
rect 18230 2836 18236 2848
rect 18095 2808 18236 2836
rect 18095 2805 18107 2808
rect 18049 2799 18107 2805
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 18506 2836 18512 2848
rect 18467 2808 18512 2836
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 22370 2836 22376 2848
rect 22331 2808 22376 2836
rect 22370 2796 22376 2808
rect 22428 2796 22434 2848
rect 24578 2836 24584 2848
rect 24539 2808 24584 2836
rect 24578 2796 24584 2808
rect 24636 2796 24642 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 1854 2632 1860 2644
rect 1443 2604 1860 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2777 2635 2835 2641
rect 2777 2632 2789 2635
rect 1995 2604 2789 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2777 2601 2789 2604
rect 2823 2632 2835 2635
rect 3878 2632 3884 2644
rect 2823 2604 3884 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5224 2604 5733 2632
rect 5224 2592 5230 2604
rect 5721 2601 5733 2604
rect 5767 2601 5779 2635
rect 6730 2632 6736 2644
rect 6691 2604 6736 2632
rect 5721 2595 5779 2601
rect 2406 2524 2412 2576
rect 2464 2564 2470 2576
rect 3697 2567 3755 2573
rect 3697 2564 3709 2567
rect 2464 2536 3709 2564
rect 2464 2524 2470 2536
rect 3697 2533 3709 2536
rect 3743 2564 3755 2567
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 3743 2536 3801 2564
rect 3743 2533 3755 2536
rect 3697 2527 3755 2533
rect 3789 2533 3801 2536
rect 3835 2533 3847 2567
rect 5736 2564 5764 2595
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10928 2604 10977 2632
rect 10928 2592 10934 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 12066 2632 12072 2644
rect 12027 2604 12072 2632
rect 10965 2595 11023 2601
rect 12066 2592 12072 2604
rect 12124 2632 12130 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 12124 2604 12357 2632
rect 12124 2592 12130 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 12345 2595 12403 2601
rect 7184 2567 7242 2573
rect 7184 2564 7196 2567
rect 5736 2536 7196 2564
rect 3789 2527 3847 2533
rect 7184 2533 7196 2536
rect 7230 2564 7242 2567
rect 7742 2564 7748 2576
rect 7230 2536 7748 2564
rect 7230 2533 7242 2536
rect 7184 2527 7242 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 3513 2499 3571 2505
rect 3513 2465 3525 2499
rect 3559 2496 3571 2499
rect 4608 2499 4666 2505
rect 4608 2496 4620 2499
rect 3559 2468 4620 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 4608 2465 4620 2468
rect 4654 2496 4666 2499
rect 6362 2496 6368 2508
rect 4654 2468 6368 2496
rect 4654 2465 4666 2468
rect 4608 2459 4666 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6788 2468 6929 2496
rect 6788 2456 6794 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9858 2496 9864 2508
rect 9263 2468 9864 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 10410 2456 10416 2508
rect 10468 2496 10474 2508
rect 11330 2496 11336 2508
rect 10468 2468 11336 2496
rect 10468 2456 10474 2468
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 12360 2496 12388 2595
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 16206 2632 16212 2644
rect 16167 2604 16212 2632
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 16390 2632 16396 2644
rect 16351 2604 16396 2632
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2632 18110 2644
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18104 2604 18797 2632
rect 18104 2592 18110 2604
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 18785 2595 18843 2601
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 20070 2632 20076 2644
rect 19751 2604 20076 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 20441 2635 20499 2641
rect 20441 2632 20453 2635
rect 20220 2604 20453 2632
rect 20220 2592 20226 2604
rect 20441 2601 20453 2604
rect 20487 2601 20499 2635
rect 24762 2632 24768 2644
rect 24723 2604 24768 2632
rect 20441 2595 20499 2601
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 13814 2524 13820 2576
rect 13872 2524 13878 2576
rect 16224 2564 16252 2592
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 16224 2536 16865 2564
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 21174 2564 21180 2576
rect 21135 2536 21180 2564
rect 16853 2527 16911 2533
rect 21174 2524 21180 2536
rect 21232 2524 21238 2576
rect 23385 2567 23443 2573
rect 23385 2564 23397 2567
rect 22940 2536 23397 2564
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12360 2468 12909 2496
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13164 2499 13222 2505
rect 13164 2465 13176 2499
rect 13210 2496 13222 2499
rect 13832 2496 13860 2524
rect 22940 2508 22968 2536
rect 23385 2533 23397 2536
rect 23431 2533 23443 2567
rect 23385 2527 23443 2533
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 13210 2468 14841 2496
rect 13210 2465 13222 2468
rect 13164 2459 13222 2465
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 15838 2456 15844 2508
rect 15896 2496 15902 2508
rect 16761 2499 16819 2505
rect 16761 2496 16773 2499
rect 15896 2468 16773 2496
rect 15896 2456 15902 2468
rect 16761 2465 16773 2468
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2465 18751 2499
rect 19886 2496 19892 2508
rect 19847 2468 19892 2496
rect 18693 2459 18751 2465
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2240 2400 2881 2428
rect 2240 2304 2268 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3418 2428 3424 2440
rect 3099 2400 3424 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 3697 2431 3755 2437
rect 3697 2397 3709 2431
rect 3743 2428 3755 2431
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 3743 2400 4353 2428
rect 3743 2397 3755 2400
rect 3697 2391 3755 2397
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2397 11483 2431
rect 11606 2428 11612 2440
rect 11567 2400 11612 2428
rect 11425 2391 11483 2397
rect 2409 2363 2467 2369
rect 2409 2329 2421 2363
rect 2455 2360 2467 2363
rect 2682 2360 2688 2372
rect 2455 2332 2688 2360
rect 2455 2329 2467 2332
rect 2409 2323 2467 2329
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 11440 2360 11468 2391
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 16850 2428 16856 2440
rect 15335 2400 16856 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 16850 2388 16856 2400
rect 16908 2428 16914 2440
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 16908 2400 16957 2428
rect 16908 2388 16914 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 12342 2360 12348 2372
rect 11440 2332 12348 2360
rect 2222 2292 2228 2304
rect 2183 2264 2228 2292
rect 2222 2252 2228 2264
rect 2280 2252 2286 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10410 2292 10416 2304
rect 10371 2264 10416 2292
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 10778 2292 10784 2304
rect 10739 2264 10784 2292
rect 10778 2252 10784 2264
rect 10836 2292 10842 2304
rect 11440 2292 11468 2332
rect 12342 2320 12348 2332
rect 12400 2320 12406 2372
rect 17678 2360 17684 2372
rect 17639 2332 17684 2360
rect 17678 2320 17684 2332
rect 17736 2360 17742 2372
rect 18708 2360 18736 2459
rect 19886 2456 19892 2468
rect 19944 2496 19950 2508
rect 20809 2499 20867 2505
rect 20809 2496 20821 2499
rect 19944 2468 20821 2496
rect 19944 2456 19950 2468
rect 20809 2465 20821 2468
rect 20855 2465 20867 2499
rect 22922 2496 22928 2508
rect 22883 2468 22928 2496
rect 20809 2459 20867 2465
rect 22922 2456 22928 2468
rect 22980 2456 22986 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23124 2468 24593 2496
rect 18969 2431 19027 2437
rect 18969 2397 18981 2431
rect 19015 2428 19027 2431
rect 19242 2428 19248 2440
rect 19015 2400 19248 2428
rect 19015 2397 19027 2400
rect 18969 2391 19027 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 23124 2369 23152 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 17736 2332 18736 2360
rect 23109 2363 23167 2369
rect 17736 2320 17742 2332
rect 23109 2329 23121 2363
rect 23155 2329 23167 2363
rect 23109 2323 23167 2329
rect 10836 2264 11468 2292
rect 10836 2252 10842 2264
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 15654 2292 15660 2304
rect 13688 2264 15660 2292
rect 13688 2252 13694 2264
rect 15654 2252 15660 2264
rect 15712 2252 15718 2304
rect 15838 2292 15844 2304
rect 15799 2264 15844 2292
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 18322 2292 18328 2304
rect 18283 2264 18328 2292
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 18506 2252 18512 2304
rect 18564 2292 18570 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 18564 2264 20085 2292
rect 18564 2252 18570 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 7190 620 7196 672
rect 7248 660 7254 672
rect 7248 632 8248 660
rect 7248 620 7254 632
rect 8220 604 8248 632
rect 8202 552 8208 604
rect 8260 552 8266 604
rect 21542 552 21548 604
rect 21600 592 21606 604
rect 21910 592 21916 604
rect 21600 564 21916 592
rect 21600 552 21606 564
rect 21910 552 21916 564
rect 21968 552 21974 604
<< via1 >>
rect 3332 27072 3384 27124
rect 6276 27072 6328 27124
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 2504 24216 2556 24268
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1492 23808 1544 23860
rect 2688 23851 2740 23860
rect 2688 23817 2697 23851
rect 2697 23817 2731 23851
rect 2731 23817 2740 23851
rect 2688 23808 2740 23817
rect 3148 23579 3200 23588
rect 3148 23545 3157 23579
rect 3157 23545 3191 23579
rect 3191 23545 3200 23579
rect 3148 23536 3200 23545
rect 2044 23511 2096 23520
rect 2044 23477 2053 23511
rect 2053 23477 2087 23511
rect 2087 23477 2096 23511
rect 2044 23468 2096 23477
rect 2504 23468 2556 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1400 23264 1452 23316
rect 2412 23128 2464 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1676 22720 1728 22772
rect 2044 22627 2096 22636
rect 2044 22593 2053 22627
rect 2053 22593 2087 22627
rect 2087 22593 2096 22627
rect 2044 22584 2096 22593
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1860 22040 1912 22092
rect 1584 21947 1636 21956
rect 1584 21913 1593 21947
rect 1593 21913 1627 21947
rect 1627 21913 1636 21947
rect 1584 21904 1636 21913
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1860 21292 1912 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1492 21088 1544 21140
rect 1676 20952 1728 21004
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1676 20383 1728 20392
rect 1676 20349 1685 20383
rect 1685 20349 1719 20383
rect 1719 20349 1728 20383
rect 1676 20340 1728 20349
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 1676 19864 1728 19916
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 11612 19252 11664 19304
rect 12072 19252 12124 19304
rect 12716 19252 12768 19304
rect 13268 19252 13320 19304
rect 9956 19116 10008 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 7748 18411 7800 18420
rect 7748 18377 7757 18411
rect 7757 18377 7791 18411
rect 7791 18377 7800 18411
rect 7748 18368 7800 18377
rect 2872 18028 2924 18080
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 8208 18028 8260 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1400 17824 1452 17876
rect 1584 17688 1636 17740
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17212 1636 17264
rect 14280 17212 14332 17264
rect 14740 17212 14792 17264
rect 3056 17119 3108 17128
rect 3056 17085 3065 17119
rect 3065 17085 3099 17119
rect 3099 17085 3108 17119
rect 3056 17076 3108 17085
rect 1492 16940 1544 16992
rect 2044 16983 2096 16992
rect 2044 16949 2053 16983
rect 2053 16949 2087 16983
rect 2087 16949 2096 16983
rect 2044 16940 2096 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 5724 16779 5776 16788
rect 5724 16745 5733 16779
rect 5733 16745 5767 16779
rect 5767 16745 5776 16779
rect 5724 16736 5776 16745
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 6552 16600 6604 16652
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 5448 16235 5500 16244
rect 5448 16201 5457 16235
rect 5457 16201 5491 16235
rect 5491 16201 5500 16235
rect 5448 16192 5500 16201
rect 6092 16192 6144 16244
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 5908 15963 5960 15972
rect 5908 15929 5917 15963
rect 5917 15929 5951 15963
rect 5951 15929 5960 15963
rect 5908 15920 5960 15929
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 6552 15648 6604 15700
rect 6276 15580 6328 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 4620 15308 4672 15360
rect 6920 15308 6972 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 6552 15104 6604 15156
rect 8116 15104 8168 15156
rect 1400 15036 1452 15088
rect 6276 15036 6328 15088
rect 6644 15036 6696 15088
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 4252 14832 4304 14884
rect 6552 14832 6604 14884
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 6460 14764 6512 14816
rect 7196 14764 7248 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1492 14560 1544 14612
rect 4252 14603 4304 14612
rect 4252 14569 4261 14603
rect 4261 14569 4295 14603
rect 4295 14569 4304 14603
rect 4252 14560 4304 14569
rect 6552 14560 6604 14612
rect 4712 14492 4764 14544
rect 5540 14492 5592 14544
rect 2044 14424 2096 14476
rect 6736 14424 6788 14476
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 4620 14016 4672 14068
rect 5540 13948 5592 14000
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 2688 13812 2740 13864
rect 6736 13948 6788 14000
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 5448 13744 5500 13796
rect 6552 13719 6604 13728
rect 6552 13685 6561 13719
rect 6561 13685 6595 13719
rect 6595 13685 6604 13719
rect 6552 13676 6604 13685
rect 6920 13676 6972 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1400 13472 1452 13524
rect 2688 13515 2740 13524
rect 2688 13481 2697 13515
rect 2697 13481 2731 13515
rect 2731 13481 2740 13515
rect 2688 13472 2740 13481
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 7380 13472 7432 13524
rect 5540 13404 5592 13456
rect 6644 13404 6696 13456
rect 6920 13447 6972 13456
rect 6920 13413 6929 13447
rect 6929 13413 6963 13447
rect 6963 13413 6972 13447
rect 6920 13404 6972 13413
rect 1676 13336 1728 13388
rect 2228 13336 2280 13388
rect 3332 13336 3384 13388
rect 5448 13336 5500 13388
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 2688 13132 2740 13184
rect 3884 13175 3936 13184
rect 3884 13141 3893 13175
rect 3893 13141 3927 13175
rect 3927 13141 3936 13175
rect 3884 13132 3936 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 3332 12971 3384 12980
rect 3332 12937 3341 12971
rect 3341 12937 3375 12971
rect 3375 12937 3384 12971
rect 3332 12928 3384 12937
rect 4068 12928 4120 12980
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 2320 12724 2372 12776
rect 3332 12792 3384 12844
rect 3884 12792 3936 12844
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 2780 12656 2832 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 2320 12427 2372 12436
rect 2320 12393 2329 12427
rect 2329 12393 2363 12427
rect 2363 12393 2372 12427
rect 2320 12384 2372 12393
rect 2780 12384 2832 12436
rect 4252 12384 4304 12436
rect 5172 12384 5224 12436
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 5448 12384 5500 12393
rect 2228 12316 2280 12368
rect 4344 12359 4396 12368
rect 4344 12325 4378 12359
rect 4378 12325 4396 12359
rect 4344 12316 4396 12325
rect 1584 12248 1636 12300
rect 3700 12248 3752 12300
rect 3976 12248 4028 12300
rect 12256 12291 12308 12300
rect 12256 12257 12290 12291
rect 12290 12257 12308 12291
rect 12256 12248 12308 12257
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 4068 12044 4120 12096
rect 12716 12044 12768 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 3700 11883 3752 11892
rect 3700 11849 3709 11883
rect 3709 11849 3743 11883
rect 3743 11849 3752 11883
rect 3700 11840 3752 11849
rect 12256 11840 12308 11892
rect 2872 11636 2924 11688
rect 8852 11636 8904 11688
rect 4068 11611 4120 11620
rect 4068 11577 4102 11611
rect 4102 11577 4120 11611
rect 4068 11568 4120 11577
rect 2688 11500 2740 11552
rect 4344 11500 4396 11552
rect 11980 11500 12032 11552
rect 13176 11500 13228 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3700 11296 3752 11348
rect 4344 11339 4396 11348
rect 4344 11305 4353 11339
rect 4353 11305 4387 11339
rect 4387 11305 4396 11339
rect 4344 11296 4396 11305
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 4988 11160 5040 11212
rect 3608 11092 3660 11144
rect 5448 11024 5500 11076
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3608 10795 3660 10804
rect 3608 10761 3617 10795
rect 3617 10761 3651 10795
rect 3651 10761 3660 10795
rect 3608 10752 3660 10761
rect 4436 10752 4488 10804
rect 2780 10684 2832 10736
rect 4068 10616 4120 10668
rect 5448 10616 5500 10668
rect 3608 10548 3660 10600
rect 1584 10412 1636 10464
rect 2504 10412 2556 10464
rect 4712 10412 4764 10464
rect 4988 10412 5040 10464
rect 5448 10412 5500 10464
rect 9680 10412 9732 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 4068 10208 4120 10260
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 6368 10140 6420 10192
rect 2504 10072 2556 10124
rect 6644 10072 6696 10124
rect 11060 10072 11112 10124
rect 17224 10115 17276 10124
rect 17224 10081 17258 10115
rect 17258 10081 17276 10115
rect 17224 10072 17276 10081
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 2780 9936 2832 9988
rect 6828 9936 6880 9988
rect 9864 10004 9916 10056
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 8392 9936 8444 9988
rect 18328 9979 18380 9988
rect 18328 9945 18337 9979
rect 18337 9945 18371 9979
rect 18371 9945 18380 9979
rect 18328 9936 18380 9945
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 1768 9868 1820 9920
rect 4160 9868 4212 9920
rect 5356 9868 5408 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 8208 9868 8260 9920
rect 11612 9868 11664 9920
rect 11888 9868 11940 9920
rect 12440 9868 12492 9920
rect 13544 9868 13596 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2872 9664 2924 9716
rect 4712 9664 4764 9716
rect 6736 9664 6788 9716
rect 7196 9664 7248 9716
rect 7748 9664 7800 9716
rect 11060 9707 11112 9716
rect 11060 9673 11069 9707
rect 11069 9673 11103 9707
rect 11103 9673 11112 9707
rect 11060 9664 11112 9673
rect 17224 9664 17276 9716
rect 18236 9596 18288 9648
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 5540 9528 5592 9580
rect 6184 9528 6236 9580
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 9588 9503 9640 9512
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 10968 9460 11020 9512
rect 3148 9392 3200 9444
rect 6920 9392 6972 9444
rect 7196 9392 7248 9444
rect 10048 9392 10100 9444
rect 1952 9324 2004 9376
rect 2136 9324 2188 9376
rect 2688 9324 2740 9376
rect 3332 9324 3384 9376
rect 6368 9324 6420 9376
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 7380 9324 7432 9376
rect 10968 9324 11020 9376
rect 12164 9324 12216 9376
rect 13084 9324 13136 9376
rect 14372 9460 14424 9512
rect 13544 9435 13596 9444
rect 13544 9401 13578 9435
rect 13578 9401 13596 9435
rect 13544 9392 13596 9401
rect 14280 9324 14332 9376
rect 16948 9324 17000 9376
rect 17500 9324 17552 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2044 9120 2096 9172
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 6092 9163 6144 9172
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 8300 9120 8352 9172
rect 7380 9095 7432 9104
rect 7380 9061 7414 9095
rect 7414 9061 7432 9095
rect 7380 9052 7432 9061
rect 2320 8984 2372 9036
rect 4620 8984 4672 9036
rect 7196 8984 7248 9036
rect 9680 9120 9732 9172
rect 10140 9120 10192 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 14280 9163 14332 9172
rect 14280 9129 14289 9163
rect 14289 9129 14323 9163
rect 14323 9129 14332 9163
rect 14280 9120 14332 9129
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 9772 9052 9824 9104
rect 10968 9052 11020 9104
rect 12440 9095 12492 9104
rect 12440 9061 12474 9095
rect 12474 9061 12492 9095
rect 12440 9052 12492 9061
rect 16120 8984 16172 9036
rect 22192 9027 22244 9036
rect 22192 8993 22201 9027
rect 22201 8993 22235 9027
rect 22235 8993 22244 9027
rect 22192 8984 22244 8993
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 2872 8916 2924 8968
rect 3608 8916 3660 8968
rect 3976 8916 4028 8968
rect 10048 8916 10100 8968
rect 12164 8959 12216 8968
rect 12164 8925 12173 8959
rect 12173 8925 12207 8959
rect 12207 8925 12216 8959
rect 12164 8916 12216 8925
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 8392 8848 8444 8900
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 2228 8780 2280 8832
rect 4252 8780 4304 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 6920 8780 6972 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 16488 8780 16540 8832
rect 23480 8780 23532 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 7380 8576 7432 8628
rect 8116 8576 8168 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 12440 8576 12492 8628
rect 1400 8551 1452 8560
rect 1400 8517 1409 8551
rect 1409 8517 1443 8551
rect 1443 8517 1452 8551
rect 1400 8508 1452 8517
rect 9496 8508 9548 8560
rect 10048 8508 10100 8560
rect 1676 8440 1728 8492
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 11060 8440 11112 8492
rect 12164 8440 12216 8492
rect 12900 8483 12952 8492
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 2044 8372 2096 8424
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 4068 8372 4120 8424
rect 4252 8415 4304 8424
rect 4252 8381 4286 8415
rect 4286 8381 4304 8415
rect 4252 8372 4304 8381
rect 2320 8304 2372 8356
rect 4436 8304 4488 8356
rect 5172 8304 5224 8356
rect 6920 8304 6972 8356
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 5356 8236 5408 8245
rect 7196 8236 7248 8288
rect 12348 8372 12400 8424
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 15660 8576 15712 8628
rect 22192 8576 22244 8628
rect 17868 8508 17920 8560
rect 22100 8508 22152 8560
rect 8392 8304 8444 8356
rect 10968 8304 11020 8356
rect 12072 8304 12124 8356
rect 8300 8236 8352 8288
rect 12532 8236 12584 8288
rect 14280 8372 14332 8424
rect 16856 8415 16908 8424
rect 16856 8381 16865 8415
rect 16865 8381 16899 8415
rect 16899 8381 16908 8415
rect 16856 8372 16908 8381
rect 21640 8415 21692 8424
rect 21640 8381 21649 8415
rect 21649 8381 21683 8415
rect 21683 8381 21692 8415
rect 21640 8372 21692 8381
rect 16120 8347 16172 8356
rect 16120 8313 16129 8347
rect 16129 8313 16163 8347
rect 16163 8313 16172 8347
rect 16120 8304 16172 8313
rect 14372 8236 14424 8288
rect 15568 8279 15620 8288
rect 15568 8245 15577 8279
rect 15577 8245 15611 8279
rect 15611 8245 15620 8279
rect 15568 8236 15620 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1768 8032 1820 8084
rect 4068 8032 4120 8084
rect 6460 8075 6512 8084
rect 6460 8041 6469 8075
rect 6469 8041 6503 8075
rect 6503 8041 6512 8075
rect 6460 8032 6512 8041
rect 6920 8032 6972 8084
rect 7656 8032 7708 8084
rect 8392 8032 8444 8084
rect 9496 8075 9548 8084
rect 9496 8041 9505 8075
rect 9505 8041 9539 8075
rect 9539 8041 9548 8075
rect 9496 8032 9548 8041
rect 12072 8032 12124 8084
rect 12440 8032 12492 8084
rect 12900 8032 12952 8084
rect 13820 8032 13872 8084
rect 15660 8075 15712 8084
rect 15660 8041 15669 8075
rect 15669 8041 15703 8075
rect 15703 8041 15712 8075
rect 15660 8032 15712 8041
rect 17224 8075 17276 8084
rect 17224 8041 17233 8075
rect 17233 8041 17267 8075
rect 17267 8041 17276 8075
rect 17224 8032 17276 8041
rect 8300 7964 8352 8016
rect 9588 7964 9640 8016
rect 10140 7964 10192 8016
rect 15844 7964 15896 8016
rect 1768 7939 1820 7948
rect 1768 7905 1777 7939
rect 1777 7905 1811 7939
rect 1811 7905 1820 7939
rect 1768 7896 1820 7905
rect 5172 7896 5224 7948
rect 5356 7939 5408 7948
rect 5356 7905 5390 7939
rect 5390 7905 5408 7939
rect 5356 7896 5408 7905
rect 6920 7896 6972 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 21088 7939 21140 7948
rect 21088 7905 21097 7939
rect 21097 7905 21131 7939
rect 21131 7905 21140 7939
rect 21088 7896 21140 7905
rect 22100 7896 22152 7948
rect 22744 7939 22796 7948
rect 22744 7905 22753 7939
rect 22753 7905 22787 7939
rect 22787 7905 22796 7939
rect 22744 7896 22796 7905
rect 23848 7939 23900 7948
rect 23848 7905 23857 7939
rect 23857 7905 23891 7939
rect 23891 7905 23900 7939
rect 23848 7896 23900 7905
rect 1584 7828 1636 7880
rect 2872 7828 2924 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 12532 7828 12584 7880
rect 14280 7871 14332 7880
rect 7564 7803 7616 7812
rect 7564 7769 7573 7803
rect 7573 7769 7607 7803
rect 7607 7769 7616 7803
rect 7564 7760 7616 7769
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 18420 7871 18472 7880
rect 17408 7828 17460 7837
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 17960 7760 18012 7812
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 4620 7735 4672 7744
rect 2780 7692 2832 7701
rect 4620 7701 4629 7735
rect 4629 7701 4663 7735
rect 4663 7701 4672 7735
rect 4620 7692 4672 7701
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 4896 7692 4948 7701
rect 8392 7692 8444 7744
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 15292 7735 15344 7744
rect 15292 7701 15301 7735
rect 15301 7701 15335 7735
rect 15335 7701 15344 7735
rect 15292 7692 15344 7701
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 18880 7735 18932 7744
rect 18880 7701 18889 7735
rect 18889 7701 18923 7735
rect 18923 7701 18932 7735
rect 18880 7692 18932 7701
rect 22100 7692 22152 7744
rect 22928 7735 22980 7744
rect 22928 7701 22937 7735
rect 22937 7701 22971 7735
rect 22971 7701 22980 7735
rect 22928 7692 22980 7701
rect 24032 7735 24084 7744
rect 24032 7701 24041 7735
rect 24041 7701 24075 7735
rect 24075 7701 24084 7735
rect 24032 7692 24084 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1676 7488 1728 7540
rect 4896 7488 4948 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 9312 7531 9364 7540
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2780 7352 2832 7404
rect 2964 7352 3016 7404
rect 3976 7352 4028 7404
rect 6920 7420 6972 7472
rect 8392 7395 8444 7404
rect 3516 7284 3568 7336
rect 5356 7284 5408 7336
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 11704 7488 11756 7540
rect 12256 7488 12308 7540
rect 12532 7531 12584 7540
rect 12532 7497 12541 7531
rect 12541 7497 12575 7531
rect 12575 7497 12584 7531
rect 12532 7488 12584 7497
rect 13820 7488 13872 7540
rect 14372 7488 14424 7540
rect 15476 7488 15528 7540
rect 15844 7488 15896 7540
rect 15936 7488 15988 7540
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 21088 7488 21140 7540
rect 22744 7531 22796 7540
rect 22744 7497 22753 7531
rect 22753 7497 22787 7531
rect 22787 7497 22796 7531
rect 22744 7488 22796 7497
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 10968 7352 11020 7404
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 13544 7420 13596 7472
rect 15660 7420 15712 7472
rect 17224 7420 17276 7472
rect 23848 7420 23900 7472
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 17500 7284 17552 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 20536 7327 20588 7336
rect 20536 7293 20545 7327
rect 20545 7293 20579 7327
rect 20579 7293 20588 7327
rect 20536 7284 20588 7293
rect 23480 7284 23532 7336
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 2136 7191 2188 7200
rect 2136 7157 2145 7191
rect 2145 7157 2179 7191
rect 2179 7157 2188 7191
rect 2136 7148 2188 7157
rect 2412 7148 2464 7200
rect 3148 7148 3200 7200
rect 3976 7191 4028 7200
rect 3976 7157 3985 7191
rect 3985 7157 4019 7191
rect 4019 7157 4028 7191
rect 3976 7148 4028 7157
rect 5172 7148 5224 7200
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 12808 7216 12860 7268
rect 14832 7216 14884 7268
rect 18880 7216 18932 7268
rect 9772 7148 9824 7200
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 19432 7191 19484 7200
rect 19432 7157 19441 7191
rect 19441 7157 19475 7191
rect 19475 7157 19484 7191
rect 19432 7148 19484 7157
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 23848 7191 23900 7200
rect 23848 7157 23857 7191
rect 23857 7157 23891 7191
rect 23891 7157 23900 7191
rect 23848 7148 23900 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2136 6944 2188 6996
rect 3516 6987 3568 6996
rect 1676 6740 1728 6792
rect 1860 6604 1912 6656
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 4068 6944 4120 6996
rect 5448 6944 5500 6996
rect 7196 6944 7248 6996
rect 8116 6944 8168 6996
rect 8392 6944 8444 6996
rect 12808 6944 12860 6996
rect 8208 6919 8260 6928
rect 8208 6885 8217 6919
rect 8217 6885 8251 6919
rect 8251 6885 8260 6919
rect 8208 6876 8260 6885
rect 9772 6876 9824 6928
rect 3884 6808 3936 6860
rect 5448 6808 5500 6860
rect 2504 6740 2556 6792
rect 3148 6740 3200 6792
rect 5172 6740 5224 6792
rect 3240 6604 3292 6656
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 6276 6604 6328 6656
rect 6460 6604 6512 6656
rect 6920 6740 6972 6792
rect 8392 6740 8444 6792
rect 9680 6808 9732 6860
rect 8576 6740 8628 6792
rect 9312 6740 9364 6792
rect 10876 6808 10928 6860
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 9496 6715 9548 6724
rect 9496 6681 9505 6715
rect 9505 6681 9539 6715
rect 9539 6681 9548 6715
rect 10968 6740 11020 6792
rect 11152 6740 11204 6792
rect 9496 6672 9548 6681
rect 10784 6672 10836 6724
rect 12440 6740 12492 6792
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 15752 6944 15804 6996
rect 16212 6987 16264 6996
rect 16212 6953 16221 6987
rect 16221 6953 16255 6987
rect 16255 6953 16264 6987
rect 16212 6944 16264 6953
rect 16948 6987 17000 6996
rect 16948 6953 16957 6987
rect 16957 6953 16991 6987
rect 16991 6953 17000 6987
rect 16948 6944 17000 6953
rect 17408 6944 17460 6996
rect 18880 6944 18932 6996
rect 15476 6919 15528 6928
rect 15476 6885 15485 6919
rect 15485 6885 15519 6919
rect 15519 6885 15528 6919
rect 15476 6876 15528 6885
rect 15936 6740 15988 6792
rect 18052 6808 18104 6860
rect 22100 6808 22152 6860
rect 22560 6808 22612 6860
rect 24032 6808 24084 6860
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 8300 6604 8352 6656
rect 11244 6604 11296 6656
rect 11612 6647 11664 6656
rect 11612 6613 11621 6647
rect 11621 6613 11655 6647
rect 11655 6613 11664 6647
rect 11612 6604 11664 6613
rect 14832 6604 14884 6656
rect 15844 6647 15896 6656
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 22376 6647 22428 6656
rect 22376 6613 22385 6647
rect 22385 6613 22419 6647
rect 22419 6613 22428 6647
rect 22376 6604 22428 6613
rect 24124 6647 24176 6656
rect 24124 6613 24133 6647
rect 24133 6613 24167 6647
rect 24167 6613 24176 6647
rect 24124 6604 24176 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 3056 6400 3108 6452
rect 1676 6264 1728 6316
rect 3240 6264 3292 6316
rect 5172 6400 5224 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 11520 6400 11572 6452
rect 13820 6400 13872 6452
rect 15752 6400 15804 6452
rect 18880 6400 18932 6452
rect 22560 6443 22612 6452
rect 22560 6409 22569 6443
rect 22569 6409 22603 6443
rect 22603 6409 22612 6443
rect 22560 6400 22612 6409
rect 24032 6443 24084 6452
rect 24032 6409 24041 6443
rect 24041 6409 24075 6443
rect 24075 6409 24084 6443
rect 24032 6400 24084 6409
rect 6276 6307 6328 6316
rect 6276 6273 6285 6307
rect 6285 6273 6319 6307
rect 6319 6273 6328 6307
rect 6276 6264 6328 6273
rect 7196 6264 7248 6316
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 848 6196 900 6248
rect 2872 6128 2924 6180
rect 4344 6196 4396 6248
rect 6368 6196 6420 6248
rect 6920 6196 6972 6248
rect 10968 6196 11020 6248
rect 11888 6196 11940 6248
rect 13084 6196 13136 6248
rect 15752 6239 15804 6248
rect 15752 6205 15786 6239
rect 15786 6205 15804 6239
rect 15752 6196 15804 6205
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 20720 6196 20772 6248
rect 7748 6128 7800 6180
rect 10784 6128 10836 6180
rect 18328 6128 18380 6180
rect 2504 6060 2556 6112
rect 3884 6060 3936 6112
rect 5356 6060 5408 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 11336 6060 11388 6112
rect 11980 6060 12032 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 15936 6060 15988 6112
rect 16948 6060 17000 6112
rect 17500 6103 17552 6112
rect 17500 6069 17509 6103
rect 17509 6069 17543 6103
rect 17543 6069 17552 6103
rect 17500 6060 17552 6069
rect 19248 6060 19300 6112
rect 20168 6103 20220 6112
rect 20168 6069 20177 6103
rect 20177 6069 20211 6103
rect 20211 6069 20220 6103
rect 20168 6060 20220 6069
rect 21916 6060 21968 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 4160 5856 4212 5908
rect 4896 5856 4948 5908
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 8576 5856 8628 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 11152 5899 11204 5908
rect 11152 5865 11161 5899
rect 11161 5865 11195 5899
rect 11195 5865 11204 5899
rect 11152 5856 11204 5865
rect 13084 5856 13136 5908
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 16212 5856 16264 5908
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 1676 5788 1728 5840
rect 1952 5788 2004 5840
rect 2780 5788 2832 5840
rect 10232 5788 10284 5840
rect 10784 5831 10836 5840
rect 10784 5797 10793 5831
rect 10793 5797 10827 5831
rect 10827 5797 10836 5831
rect 10784 5788 10836 5797
rect 11520 5831 11572 5840
rect 11520 5797 11554 5831
rect 11554 5797 11572 5831
rect 11520 5788 11572 5797
rect 12164 5788 12216 5840
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 16948 5831 17000 5840
rect 16948 5797 16982 5831
rect 16982 5797 17000 5831
rect 16948 5788 17000 5797
rect 17960 5788 18012 5840
rect 18512 5788 18564 5840
rect 4712 5720 4764 5772
rect 6276 5720 6328 5772
rect 6460 5720 6512 5772
rect 7012 5720 7064 5772
rect 7196 5720 7248 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10968 5720 11020 5772
rect 14188 5763 14240 5772
rect 14188 5729 14197 5763
rect 14197 5729 14231 5763
rect 14231 5729 14240 5763
rect 14188 5720 14240 5729
rect 4344 5584 4396 5636
rect 8668 5652 8720 5704
rect 9588 5584 9640 5636
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15476 5720 15528 5772
rect 17500 5720 17552 5772
rect 19156 5763 19208 5772
rect 19156 5729 19165 5763
rect 19165 5729 19199 5763
rect 19199 5729 19208 5763
rect 19156 5720 19208 5729
rect 20168 5720 20220 5772
rect 20904 5720 20956 5772
rect 15016 5652 15068 5661
rect 11060 5584 11112 5636
rect 2872 5516 2924 5568
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 4160 5516 4212 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 5448 5516 5500 5568
rect 6092 5559 6144 5568
rect 6092 5525 6101 5559
rect 6101 5525 6135 5559
rect 6135 5525 6144 5559
rect 6092 5516 6144 5525
rect 8208 5516 8260 5568
rect 8392 5559 8444 5568
rect 8392 5525 8401 5559
rect 8401 5525 8435 5559
rect 8435 5525 8444 5559
rect 8392 5516 8444 5525
rect 12440 5516 12492 5568
rect 15844 5516 15896 5568
rect 19340 5559 19392 5568
rect 19340 5525 19349 5559
rect 19349 5525 19383 5559
rect 19383 5525 19392 5559
rect 19340 5516 19392 5525
rect 21180 5559 21232 5568
rect 21180 5525 21189 5559
rect 21189 5525 21223 5559
rect 21223 5525 21232 5559
rect 21180 5516 21232 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2228 5312 2280 5364
rect 2412 5244 2464 5296
rect 2596 5176 2648 5228
rect 3240 5312 3292 5364
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 6276 5312 6328 5364
rect 6828 5355 6880 5364
rect 6828 5321 6837 5355
rect 6837 5321 6871 5355
rect 6871 5321 6880 5355
rect 6828 5312 6880 5321
rect 7748 5312 7800 5364
rect 10784 5312 10836 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11612 5312 11664 5364
rect 11888 5355 11940 5364
rect 11888 5321 11897 5355
rect 11897 5321 11931 5355
rect 11931 5321 11940 5355
rect 11888 5312 11940 5321
rect 4896 5287 4948 5296
rect 4896 5253 4905 5287
rect 4905 5253 4939 5287
rect 4939 5253 4948 5287
rect 4896 5244 4948 5253
rect 10048 5244 10100 5296
rect 17500 5312 17552 5364
rect 19156 5355 19208 5364
rect 19156 5321 19165 5355
rect 19165 5321 19199 5355
rect 19199 5321 19208 5355
rect 19156 5312 19208 5321
rect 20904 5355 20956 5364
rect 20904 5321 20913 5355
rect 20913 5321 20947 5355
rect 20947 5321 20956 5355
rect 20904 5312 20956 5321
rect 16212 5287 16264 5296
rect 16212 5253 16221 5287
rect 16221 5253 16255 5287
rect 16255 5253 16264 5287
rect 16212 5244 16264 5253
rect 16948 5176 17000 5228
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 1400 5108 1452 5160
rect 3056 5108 3108 5160
rect 7840 5108 7892 5160
rect 8668 5151 8720 5160
rect 8668 5117 8702 5151
rect 8702 5117 8720 5151
rect 6276 5040 6328 5092
rect 6736 5040 6788 5092
rect 8668 5108 8720 5117
rect 16856 5108 16908 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 21088 5151 21140 5160
rect 21088 5117 21097 5151
rect 21097 5117 21131 5151
rect 21131 5117 21140 5151
rect 21088 5108 21140 5117
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22100 5108 22152 5117
rect 10232 5040 10284 5092
rect 13728 5040 13780 5092
rect 16488 5040 16540 5092
rect 1768 4972 1820 5024
rect 6828 4972 6880 5024
rect 8392 4972 8444 5024
rect 10048 4972 10100 5024
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 12164 5015 12216 5024
rect 12164 4981 12173 5015
rect 12173 4981 12207 5015
rect 12207 4981 12216 5015
rect 12164 4972 12216 4981
rect 14832 4972 14884 5024
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 22284 5015 22336 5024
rect 22284 4981 22293 5015
rect 22293 4981 22327 5015
rect 22327 4981 22336 5015
rect 22284 4972 22336 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2596 4768 2648 4820
rect 4068 4768 4120 4820
rect 5356 4768 5408 4820
rect 6092 4768 6144 4820
rect 6460 4811 6512 4820
rect 6460 4777 6469 4811
rect 6469 4777 6503 4811
rect 6503 4777 6512 4811
rect 6460 4768 6512 4777
rect 6828 4811 6880 4820
rect 6828 4777 6837 4811
rect 6837 4777 6871 4811
rect 6871 4777 6880 4811
rect 6828 4768 6880 4777
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7840 4768 7892 4820
rect 8944 4768 8996 4820
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 11428 4768 11480 4820
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 15292 4811 15344 4820
rect 15292 4777 15301 4811
rect 15301 4777 15335 4811
rect 15335 4777 15344 4811
rect 15292 4768 15344 4777
rect 16488 4768 16540 4820
rect 16948 4768 17000 4820
rect 17316 4811 17368 4820
rect 17316 4777 17325 4811
rect 17325 4777 17359 4811
rect 17359 4777 17368 4811
rect 17316 4768 17368 4777
rect 17960 4768 18012 4820
rect 18604 4768 18656 4820
rect 2044 4700 2096 4752
rect 3056 4700 3108 4752
rect 8116 4700 8168 4752
rect 8576 4700 8628 4752
rect 8668 4700 8720 4752
rect 9588 4700 9640 4752
rect 10048 4743 10100 4752
rect 10048 4709 10057 4743
rect 10057 4709 10091 4743
rect 10091 4709 10100 4743
rect 10048 4700 10100 4709
rect 2412 4632 2464 4684
rect 5632 4675 5684 4684
rect 1952 4564 2004 4616
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 15568 4700 15620 4752
rect 11060 4632 11112 4684
rect 12164 4632 12216 4684
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 14648 4632 14700 4684
rect 3056 4607 3108 4616
rect 2412 4539 2464 4548
rect 2412 4505 2421 4539
rect 2421 4505 2455 4539
rect 2455 4505 2464 4539
rect 2412 4496 2464 4505
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 3424 4564 3476 4616
rect 6184 4564 6236 4616
rect 8484 4564 8536 4616
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 15752 4607 15804 4616
rect 15752 4573 15761 4607
rect 15761 4573 15795 4607
rect 15795 4573 15804 4607
rect 15752 4564 15804 4573
rect 3792 4539 3844 4548
rect 3792 4505 3801 4539
rect 3801 4505 3835 4539
rect 3835 4505 3844 4539
rect 3792 4496 3844 4505
rect 4344 4496 4396 4548
rect 13084 4539 13136 4548
rect 13084 4505 13093 4539
rect 13093 4505 13127 4539
rect 13127 4505 13136 4539
rect 13084 4496 13136 4505
rect 13360 4496 13412 4548
rect 16120 4632 16172 4684
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 17960 4632 18012 4684
rect 18604 4632 18656 4684
rect 19340 4632 19392 4684
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 21272 4632 21324 4684
rect 22008 4632 22060 4684
rect 17684 4564 17736 4616
rect 16856 4539 16908 4548
rect 16856 4505 16865 4539
rect 16865 4505 16899 4539
rect 16899 4505 16908 4539
rect 16856 4496 16908 4505
rect 1768 4428 1820 4480
rect 4712 4471 4764 4480
rect 4712 4437 4721 4471
rect 4721 4437 4755 4471
rect 4755 4437 4764 4471
rect 4712 4428 4764 4437
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 12900 4471 12952 4480
rect 12900 4437 12909 4471
rect 12909 4437 12943 4471
rect 12943 4437 12952 4471
rect 12900 4428 12952 4437
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 19524 4428 19576 4480
rect 20812 4428 20864 4480
rect 21088 4471 21140 4480
rect 21088 4437 21097 4471
rect 21097 4437 21131 4471
rect 21131 4437 21140 4471
rect 21088 4428 21140 4437
rect 22100 4471 22152 4480
rect 22100 4437 22109 4471
rect 22109 4437 22143 4471
rect 22143 4437 22152 4471
rect 22100 4428 22152 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1768 4224 1820 4276
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 3424 4267 3476 4276
rect 2780 4224 2832 4233
rect 3424 4233 3433 4267
rect 3433 4233 3467 4267
rect 3467 4233 3476 4267
rect 3424 4224 3476 4233
rect 4344 4267 4396 4276
rect 4344 4233 4353 4267
rect 4353 4233 4387 4267
rect 4387 4233 4396 4267
rect 4344 4224 4396 4233
rect 6092 4224 6144 4276
rect 8392 4224 8444 4276
rect 11980 4224 12032 4276
rect 12716 4224 12768 4276
rect 13544 4224 13596 4276
rect 296 4088 348 4140
rect 3056 4156 3108 4208
rect 3976 4156 4028 4208
rect 3608 4088 3660 4140
rect 5172 4088 5224 4140
rect 12072 4156 12124 4208
rect 12992 4156 13044 4208
rect 12900 4131 12952 4140
rect 1492 4020 1544 4072
rect 2596 4020 2648 4072
rect 8208 4020 8260 4072
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 14096 4088 14148 4140
rect 14648 4088 14700 4140
rect 15752 4224 15804 4276
rect 17316 4224 17368 4276
rect 18604 4267 18656 4276
rect 18604 4233 18613 4267
rect 18613 4233 18647 4267
rect 18647 4233 18656 4267
rect 18604 4224 18656 4233
rect 19340 4224 19392 4276
rect 21088 4224 21140 4276
rect 22008 4267 22060 4276
rect 9036 4063 9088 4072
rect 9036 4029 9059 4063
rect 9059 4029 9088 4063
rect 9036 4020 9088 4029
rect 10232 4020 10284 4072
rect 11336 4063 11388 4072
rect 11336 4029 11345 4063
rect 11345 4029 11379 4063
rect 11379 4029 11388 4063
rect 11336 4020 11388 4029
rect 13360 4020 13412 4072
rect 13820 4020 13872 4072
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14372 4020 14424 4072
rect 17224 4088 17276 4140
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 15568 4020 15620 4072
rect 18144 4020 18196 4072
rect 22008 4233 22017 4267
rect 22017 4233 22051 4267
rect 22051 4233 22060 4267
rect 22008 4224 22060 4233
rect 22468 4063 22520 4072
rect 2872 3952 2924 4004
rect 5448 3952 5500 4004
rect 6184 3952 6236 4004
rect 6920 3952 6972 4004
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 5540 3884 5592 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 8116 3884 8168 3936
rect 8300 3927 8352 3936
rect 8300 3893 8309 3927
rect 8309 3893 8343 3927
rect 8343 3893 8352 3927
rect 8300 3884 8352 3893
rect 8484 3884 8536 3936
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12164 3884 12216 3893
rect 13452 3884 13504 3936
rect 14648 3952 14700 4004
rect 19800 3995 19852 4004
rect 19800 3961 19809 3995
rect 19809 3961 19843 3995
rect 19843 3961 19852 3995
rect 19800 3952 19852 3961
rect 22468 4029 22477 4063
rect 22477 4029 22511 4063
rect 22511 4029 22520 4063
rect 22468 4020 22520 4029
rect 22284 3952 22336 4004
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 17684 3927 17736 3936
rect 17684 3893 17693 3927
rect 17693 3893 17727 3927
rect 17727 3893 17736 3927
rect 17684 3884 17736 3893
rect 17960 3884 18012 3936
rect 20260 3884 20312 3936
rect 21364 3884 21416 3936
rect 21548 3927 21600 3936
rect 21548 3893 21557 3927
rect 21557 3893 21591 3927
rect 21591 3893 21600 3927
rect 21548 3884 21600 3893
rect 22652 3927 22704 3936
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 3424 3680 3476 3732
rect 3608 3680 3660 3732
rect 4252 3723 4304 3732
rect 4252 3689 4261 3723
rect 4261 3689 4295 3723
rect 4295 3689 4304 3723
rect 4252 3680 4304 3689
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 5448 3680 5500 3732
rect 5540 3680 5592 3732
rect 9036 3680 9088 3732
rect 10784 3680 10836 3732
rect 11152 3723 11204 3732
rect 11152 3689 11161 3723
rect 11161 3689 11195 3723
rect 11195 3689 11204 3723
rect 11152 3680 11204 3689
rect 12992 3723 13044 3732
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 13452 3680 13504 3732
rect 15292 3680 15344 3732
rect 18236 3723 18288 3732
rect 18236 3689 18245 3723
rect 18245 3689 18279 3723
rect 18279 3689 18288 3723
rect 18236 3680 18288 3689
rect 19248 3680 19300 3732
rect 20168 3680 20220 3732
rect 20996 3680 21048 3732
rect 1952 3612 2004 3664
rect 5724 3655 5776 3664
rect 5724 3621 5733 3655
rect 5733 3621 5767 3655
rect 5767 3621 5776 3655
rect 5724 3612 5776 3621
rect 6184 3612 6236 3664
rect 7012 3612 7064 3664
rect 9680 3612 9732 3664
rect 11520 3655 11572 3664
rect 11520 3621 11529 3655
rect 11529 3621 11563 3655
rect 11563 3621 11572 3655
rect 11520 3612 11572 3621
rect 11980 3612 12032 3664
rect 15568 3612 15620 3664
rect 20904 3655 20956 3664
rect 20904 3621 20913 3655
rect 20913 3621 20947 3655
rect 20947 3621 20956 3655
rect 20904 3612 20956 3621
rect 1492 3587 1544 3596
rect 1492 3553 1501 3587
rect 1501 3553 1535 3587
rect 1535 3553 1544 3587
rect 1492 3544 1544 3553
rect 6092 3544 6144 3596
rect 6736 3544 6788 3596
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 9588 3476 9640 3528
rect 11520 3476 11572 3528
rect 14188 3544 14240 3596
rect 15476 3544 15528 3596
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 16764 3544 16816 3596
rect 20628 3544 20680 3596
rect 23296 3587 23348 3596
rect 23296 3553 23305 3587
rect 23305 3553 23339 3587
rect 23339 3553 23348 3587
rect 23296 3544 23348 3553
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 15384 3476 15436 3528
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 16396 3476 16448 3528
rect 8944 3408 8996 3460
rect 3700 3340 3752 3392
rect 6368 3383 6420 3392
rect 6368 3349 6377 3383
rect 6377 3349 6411 3383
rect 6411 3349 6420 3383
rect 6368 3340 6420 3349
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 15292 3383 15344 3392
rect 15292 3349 15301 3383
rect 15301 3349 15335 3383
rect 15335 3349 15344 3383
rect 15292 3340 15344 3349
rect 16764 3383 16816 3392
rect 16764 3349 16773 3383
rect 16773 3349 16807 3383
rect 16807 3349 16816 3383
rect 16764 3340 16816 3349
rect 17224 3340 17276 3392
rect 18512 3340 18564 3392
rect 19064 3340 19116 3392
rect 23480 3383 23532 3392
rect 23480 3349 23489 3383
rect 23489 3349 23523 3383
rect 23523 3349 23532 3383
rect 23480 3340 23532 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1492 3136 1544 3188
rect 3792 3136 3844 3188
rect 4896 3179 4948 3188
rect 4896 3145 4905 3179
rect 4905 3145 4939 3179
rect 4939 3145 4948 3179
rect 4896 3136 4948 3145
rect 5540 3136 5592 3188
rect 6184 3136 6236 3188
rect 9036 3136 9088 3188
rect 10968 3136 11020 3188
rect 11612 3136 11664 3188
rect 2412 3000 2464 3052
rect 6736 3068 6788 3120
rect 6368 3000 6420 3052
rect 8116 3000 8168 3052
rect 10416 3068 10468 3120
rect 9680 3000 9732 3052
rect 10784 3000 10836 3052
rect 11152 3000 11204 3052
rect 11520 3000 11572 3052
rect 12072 3000 12124 3052
rect 15660 3136 15712 3188
rect 16764 3136 16816 3188
rect 17224 3136 17276 3188
rect 19432 3136 19484 3188
rect 20628 3179 20680 3188
rect 20628 3145 20637 3179
rect 20637 3145 20671 3179
rect 20671 3145 20680 3179
rect 20628 3136 20680 3145
rect 22652 3136 22704 3188
rect 15384 3111 15436 3120
rect 15384 3077 15393 3111
rect 15393 3077 15427 3111
rect 15427 3077 15436 3111
rect 15384 3068 15436 3077
rect 20720 3068 20772 3120
rect 23296 3111 23348 3120
rect 23296 3077 23305 3111
rect 23305 3077 23339 3111
rect 23339 3077 23348 3111
rect 23296 3068 23348 3077
rect 18236 3000 18288 3052
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 3700 2932 3752 2984
rect 3976 2932 4028 2984
rect 6092 2932 6144 2984
rect 7012 2932 7064 2984
rect 8208 2932 8260 2984
rect 8944 2932 8996 2984
rect 12992 2932 13044 2984
rect 19340 2932 19392 2984
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 21088 2932 21140 2984
rect 22192 2975 22244 2984
rect 22192 2941 22201 2975
rect 22201 2941 22235 2975
rect 22235 2941 22244 2975
rect 22192 2932 22244 2941
rect 23480 2932 23532 2984
rect 4988 2864 5040 2916
rect 15844 2864 15896 2916
rect 18420 2907 18472 2916
rect 18420 2873 18429 2907
rect 18429 2873 18463 2907
rect 18463 2873 18472 2907
rect 18420 2864 18472 2873
rect 19432 2864 19484 2916
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 9772 2796 9824 2848
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 18236 2796 18288 2848
rect 18512 2839 18564 2848
rect 18512 2805 18521 2839
rect 18521 2805 18555 2839
rect 18555 2805 18564 2839
rect 18512 2796 18564 2805
rect 22376 2839 22428 2848
rect 22376 2805 22385 2839
rect 22385 2805 22419 2839
rect 22419 2805 22428 2839
rect 22376 2796 22428 2805
rect 24584 2839 24636 2848
rect 24584 2805 24593 2839
rect 24593 2805 24627 2839
rect 24627 2805 24636 2839
rect 24584 2796 24636 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1860 2592 1912 2644
rect 3884 2592 3936 2644
rect 5172 2592 5224 2644
rect 6736 2635 6788 2644
rect 2412 2524 2464 2576
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 10876 2592 10928 2644
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 14280 2635 14332 2644
rect 7748 2524 7800 2576
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 6736 2456 6788 2508
rect 9864 2499 9916 2508
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 10416 2456 10468 2508
rect 11336 2499 11388 2508
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 16212 2635 16264 2644
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 16396 2635 16448 2644
rect 16396 2601 16405 2635
rect 16405 2601 16439 2635
rect 16439 2601 16448 2635
rect 16396 2592 16448 2601
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 20076 2592 20128 2644
rect 20168 2592 20220 2644
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 13820 2524 13872 2576
rect 21180 2567 21232 2576
rect 21180 2533 21189 2567
rect 21189 2533 21223 2567
rect 21223 2533 21232 2567
rect 21180 2524 21232 2533
rect 15844 2456 15896 2508
rect 19892 2499 19944 2508
rect 3424 2388 3476 2440
rect 11612 2431 11664 2440
rect 2688 2320 2740 2372
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 16856 2388 16908 2440
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 10416 2295 10468 2304
rect 10416 2261 10425 2295
rect 10425 2261 10459 2295
rect 10459 2261 10468 2295
rect 10416 2252 10468 2261
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 12348 2320 12400 2372
rect 17684 2363 17736 2372
rect 17684 2329 17693 2363
rect 17693 2329 17727 2363
rect 17727 2329 17736 2363
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 22928 2499 22980 2508
rect 22928 2465 22937 2499
rect 22937 2465 22971 2499
rect 22971 2465 22980 2499
rect 22928 2456 22980 2465
rect 19248 2388 19300 2440
rect 17684 2320 17736 2329
rect 10784 2252 10836 2261
rect 13636 2252 13688 2304
rect 15660 2252 15712 2304
rect 15844 2295 15896 2304
rect 15844 2261 15853 2295
rect 15853 2261 15887 2295
rect 15887 2261 15896 2295
rect 15844 2252 15896 2261
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 18512 2252 18564 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 7196 620 7248 672
rect 8208 552 8260 604
rect 21548 552 21600 604
rect 21916 552 21968 604
<< metal2 >>
rect 3330 27568 3386 27577
rect 3330 27503 3386 27512
rect 3344 27130 3372 27503
rect 3332 27124 3384 27130
rect 3332 27066 3384 27072
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 2686 26888 2742 26897
rect 2686 26823 2742 26832
rect 1582 26208 1638 26217
rect 1582 26143 1638 26152
rect 1490 25528 1546 25537
rect 1490 25463 1546 25472
rect 1398 24848 1454 24857
rect 1398 24783 1454 24792
rect 1412 23322 1440 24783
rect 1504 23866 1532 25463
rect 1596 24410 1624 26143
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 1674 24168 1730 24177
rect 1674 24103 1730 24112
rect 1492 23860 1544 23866
rect 1492 23802 1544 23808
rect 1582 23488 1638 23497
rect 1582 23423 1638 23432
rect 1400 23316 1452 23322
rect 1400 23258 1452 23264
rect 1490 22808 1546 22817
rect 1490 22743 1546 22752
rect 1398 22128 1454 22137
rect 1398 22063 1454 22072
rect 1412 17882 1440 22063
rect 1504 21146 1532 22743
rect 1596 21962 1624 23423
rect 1688 22778 1716 24103
rect 2516 23526 2544 24210
rect 2700 23866 2728 26823
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 3146 23624 3202 23633
rect 3146 23559 3148 23568
rect 3200 23559 3202 23568
rect 3148 23530 3200 23536
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2504 23520 2556 23526
rect 2504 23462 2556 23468
rect 2056 23089 2084 23462
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2042 23080 2098 23089
rect 2042 23015 2098 23024
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 2042 22672 2098 22681
rect 2042 22607 2044 22616
rect 2096 22607 2098 22616
rect 2044 22578 2096 22584
rect 2424 22438 2452 23122
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1584 21956 1636 21962
rect 1584 21898 1636 21904
rect 1582 21448 1638 21457
rect 1582 21383 1638 21392
rect 1492 21140 1544 21146
rect 1492 21082 1544 21088
rect 1596 20058 1624 21383
rect 1872 21350 1900 22034
rect 2424 21457 2452 22374
rect 2410 21448 2466 21457
rect 2410 21383 2466 21392
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 1688 20398 1716 20946
rect 1676 20392 1728 20398
rect 1674 20360 1676 20369
rect 1728 20360 1730 20369
rect 1674 20295 1730 20304
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1490 18728 1546 18737
rect 1490 18663 1546 18672
rect 1400 17876 1452 17882
rect 1400 17818 1452 17824
rect 1504 16998 1532 18663
rect 1596 18426 1624 19343
rect 1688 19174 1716 19858
rect 1676 19168 1728 19174
rect 1674 19136 1676 19145
rect 1728 19136 1730 19145
rect 1674 19071 1730 19080
rect 1872 18986 1900 21286
rect 1688 18958 1900 18986
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1596 17270 1624 17682
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1596 16794 1624 17206
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1490 16008 1546 16017
rect 1490 15943 1546 15952
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 15094 1440 15506
rect 1400 15088 1452 15094
rect 1400 15030 1452 15036
rect 1398 14648 1454 14657
rect 1504 14618 1532 15943
rect 1596 15706 1624 16623
rect 1688 16153 1716 18958
rect 2516 18873 2544 23462
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 4066 20768 4122 20777
rect 4066 20703 4122 20712
rect 3330 20088 3386 20097
rect 3330 20023 3386 20032
rect 3344 19009 3372 20023
rect 4080 19281 4108 20703
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 4066 19272 4122 19281
rect 4066 19207 4122 19216
rect 3330 19000 3386 19009
rect 3330 18935 3386 18944
rect 2502 18864 2558 18873
rect 2502 18799 2558 18808
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 16833 2084 16934
rect 2042 16824 2098 16833
rect 2042 16759 2098 16768
rect 1674 16144 1730 16153
rect 1674 16079 1730 16088
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 1398 14583 1454 14592
rect 1492 14612 1544 14618
rect 1412 13530 1440 14583
rect 1492 14554 1544 14560
rect 1596 14074 1624 15263
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1582 13968 1638 13977
rect 2056 13938 2084 14418
rect 1582 13903 1638 13912
rect 2044 13932 2096 13938
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 1596 12442 1624 13903
rect 2044 13874 2096 13880
rect 2056 13841 2084 13874
rect 2688 13864 2740 13870
rect 2042 13832 2098 13841
rect 2688 13806 2740 13812
rect 2042 13767 2098 13776
rect 2700 13530 2728 13806
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 1688 12646 1716 13330
rect 2240 12646 2268 13330
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12850 2728 13126
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1596 11898 1624 12242
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1688 10985 1716 12582
rect 2240 12374 2268 12582
rect 2332 12442 2360 12718
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12442 2820 12650
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 2884 11694 2912 18022
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5446 17368 5502 17377
rect 5622 17360 5918 17380
rect 5446 17303 5502 17312
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 3068 16969 3096 17070
rect 3054 16960 3110 16969
rect 3054 16895 3110 16904
rect 5460 16250 5488 17303
rect 5722 16960 5778 16969
rect 5722 16895 5778 16904
rect 5736 16794 5764 16895
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6104 16250 6132 16594
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 5906 16008 5962 16017
rect 5906 15943 5908 15952
rect 5960 15943 5962 15952
rect 5908 15914 5960 15920
rect 5172 15904 5224 15910
rect 5170 15872 5172 15881
rect 5224 15872 5226 15881
rect 5170 15807 5226 15816
rect 6288 15638 6316 27066
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 14278 23624 14334 23633
rect 14278 23559 14334 23568
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 13910 23080 13966 23089
rect 13910 23015 13966 23024
rect 9678 22672 9734 22681
rect 9678 22607 9734 22616
rect 8298 19272 8354 19281
rect 8298 19207 8354 19216
rect 8312 19174 8340 19207
rect 8300 19168 8352 19174
rect 6734 19136 6790 19145
rect 8300 19110 8352 19116
rect 6734 19071 6790 19080
rect 6748 16697 6776 19071
rect 7746 19000 7802 19009
rect 7746 18935 7802 18944
rect 7760 18426 7788 18935
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 7470 17912 7526 17921
rect 7470 17847 7526 17856
rect 7010 16824 7066 16833
rect 7484 16794 7512 17847
rect 7010 16759 7066 16768
rect 7472 16788 7524 16794
rect 6734 16688 6790 16697
rect 6552 16652 6604 16658
rect 6734 16623 6790 16632
rect 6552 16594 6604 16600
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6380 16017 6408 16526
rect 6564 16250 6592 16594
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6366 16008 6422 16017
rect 6366 15943 6422 15952
rect 6564 15706 6592 16186
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 4264 14618 4292 14826
rect 4632 14822 4660 15302
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6288 15094 6316 15574
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4632 14074 4660 14758
rect 4724 14550 4752 14962
rect 6472 14822 6500 15438
rect 6564 15162 6592 15438
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6564 14890 6592 15098
rect 6644 15088 6696 15094
rect 6932 15042 6960 15302
rect 6644 15030 6696 15036
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6564 14618 6592 14826
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 5552 14006 5580 14486
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4172 13682 4200 13874
rect 5354 13832 5410 13841
rect 5354 13767 5410 13776
rect 5448 13796 5500 13802
rect 4080 13654 4200 13682
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3146 13288 3202 13297
rect 3146 13223 3202 13232
rect 2872 11688 2924 11694
rect 3160 11665 3188 13223
rect 3344 12986 3372 13330
rect 4080 13326 4108 13654
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3344 12850 3372 12922
rect 3896 12850 3924 13126
rect 4080 12986 4108 13262
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4080 12866 4108 12922
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3988 12838 4108 12866
rect 4158 12880 4214 12889
rect 3422 12608 3478 12617
rect 3422 12543 3478 12552
rect 3436 11801 3464 12543
rect 3988 12306 4016 12838
rect 4158 12815 4214 12824
rect 4344 12844 4396 12850
rect 4172 12782 4200 12815
rect 4344 12786 4396 12792
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3712 11898 3740 12242
rect 4068 12096 4120 12102
rect 4172 12084 4200 12718
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 12442 4292 12582
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4356 12374 4384 12786
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4120 12056 4200 12084
rect 4068 12038 4120 12044
rect 3974 11928 4030 11937
rect 3700 11892 3752 11898
rect 3974 11863 4030 11872
rect 3700 11834 3752 11840
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 2872 11630 2924 11636
rect 3146 11656 3202 11665
rect 3146 11591 3202 11600
rect 2688 11552 2740 11558
rect 2740 11500 2820 11506
rect 2688 11494 2820 11500
rect 2700 11478 2820 11494
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 2792 10742 2820 11478
rect 3712 11354 3740 11834
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3620 10810 3648 11086
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 2780 10736 2832 10742
rect 2410 10704 2466 10713
rect 2780 10678 2832 10684
rect 2410 10639 2466 10648
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 9178 1624 10406
rect 2424 10266 2452 10639
rect 3620 10606 3648 10746
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2516 10130 2544 10406
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1214 9072 1270 9081
rect 1214 9007 1270 9016
rect 1228 8537 1256 9007
rect 1400 8560 1452 8566
rect 1214 8528 1270 8537
rect 1214 8463 1270 8472
rect 1398 8528 1400 8537
rect 1452 8528 1454 8537
rect 1688 8498 1716 9862
rect 1398 8463 1454 8472
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7206 1624 7822
rect 1688 7546 1716 8434
rect 1780 8430 1808 9862
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 1964 8498 1992 9318
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8090 1808 8366
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 848 6248 900 6254
rect 848 6190 900 6196
rect 296 4140 348 4146
rect 296 4082 348 4088
rect 308 480 336 4082
rect 860 480 888 6190
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4321 1440 5102
rect 1398 4312 1454 4321
rect 1398 4247 1454 4256
rect 1412 480 1440 4247
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3602 1532 4014
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1504 3194 1532 3538
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1596 3097 1624 7142
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1780 6746 1808 7890
rect 1688 6322 1716 6734
rect 1780 6718 1900 6746
rect 1872 6662 1900 6718
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1688 5846 1716 6258
rect 1676 5840 1728 5846
rect 1676 5782 1728 5788
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4486 1808 4966
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 4282 1808 4422
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1780 4185 1808 4218
rect 1766 4176 1822 4185
rect 1766 4111 1822 4120
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 1872 2650 1900 6598
rect 1964 5846 1992 8434
rect 2056 8430 2084 9114
rect 2148 8974 2176 9318
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 2056 4758 2084 8366
rect 2240 7410 2268 8774
rect 2332 8362 2360 8978
rect 2700 8786 2728 9318
rect 2792 9058 2820 9930
rect 2884 9722 2912 9998
rect 3514 9888 3570 9897
rect 3514 9823 3570 9832
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 9178 3188 9386
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 2792 9030 3096 9058
rect 2792 8786 2820 9030
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2700 8758 2820 8786
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2148 7002 2176 7142
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2240 5370 2268 7346
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2044 4752 2096 4758
rect 2044 4694 2096 4700
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 3670 1992 4558
rect 2332 3777 2360 8298
rect 2884 7886 2912 8910
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7410 2820 7686
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 5302 2452 7142
rect 2502 6896 2558 6905
rect 2502 6831 2558 6840
rect 2516 6798 2544 6831
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2516 6118 2544 6734
rect 2884 6186 2912 7822
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2424 4690 2452 5238
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2410 4584 2466 4593
rect 2410 4519 2412 4528
rect 2464 4519 2466 4528
rect 2412 4490 2464 4496
rect 2318 3768 2374 3777
rect 2318 3703 2374 3712
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 2424 2582 2452 2994
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 1950 2000 2006 2009
rect 1950 1935 2006 1944
rect 1964 480 1992 1935
rect 2240 1737 2268 2246
rect 2226 1728 2282 1737
rect 2226 1663 2282 1672
rect 2516 480 2544 6054
rect 2884 5914 2912 6122
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2608 4826 2636 5170
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2608 4078 2636 4762
rect 2686 4720 2742 4729
rect 2686 4655 2742 4664
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2700 2378 2728 4655
rect 2792 4282 2820 5782
rect 2872 5568 2924 5574
rect 2976 5556 3004 7346
rect 3068 6458 3096 9030
rect 3160 7290 3188 9114
rect 3160 7262 3280 7290
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 6798 3188 7142
rect 3148 6792 3200 6798
rect 3252 6769 3280 7262
rect 3148 6734 3200 6740
rect 3238 6760 3294 6769
rect 3238 6695 3294 6704
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2924 5528 3004 5556
rect 2872 5510 2924 5516
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2884 4010 2912 5510
rect 3068 5166 3096 6394
rect 3252 6322 3280 6598
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3252 5370 3280 6258
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4758 3096 5102
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3068 4214 3096 4558
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2884 3738 2912 3946
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 3344 3641 3372 9318
rect 3528 7342 3556 9823
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3620 8974 3648 9522
rect 3698 9480 3754 9489
rect 3698 9415 3754 9424
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3712 7857 3740 9415
rect 3988 9217 4016 11863
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4080 10674 4108 11562
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4080 10266 4108 10610
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4172 9926 4200 12056
rect 4356 11558 4384 12310
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11354 4384 11494
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 4448 10810 4476 11154
rect 4802 10976 4858 10985
rect 4802 10911 4858 10920
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3790 9208 3846 9217
rect 3790 9143 3846 9152
rect 3974 9208 4030 9217
rect 3974 9143 4030 9152
rect 3804 8129 3832 9143
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 8430 4016 8910
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4264 8430 4292 8774
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 3882 8256 3938 8265
rect 3882 8191 3938 8200
rect 3790 8120 3846 8129
rect 3790 8055 3846 8064
rect 3698 7848 3754 7857
rect 3698 7783 3754 7792
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3528 7002 3556 7278
rect 3896 7177 3924 8191
rect 4080 8090 4108 8366
rect 4448 8362 4476 10746
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 9722 4752 10406
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4068 8084 4120 8090
rect 3988 8044 4068 8072
rect 3988 7410 4016 8044
rect 4068 8026 4120 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3976 7200 4028 7206
rect 3882 7168 3938 7177
rect 3976 7142 4028 7148
rect 3882 7103 3938 7112
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3896 6118 3924 6802
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3436 4282 3464 4558
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 3738 3648 4082
rect 3698 3768 3754 3777
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3608 3732 3660 3738
rect 3698 3703 3754 3712
rect 3608 3674 3660 3680
rect 3330 3632 3386 3641
rect 3330 3567 3386 3576
rect 3436 2446 3464 3674
rect 3712 3398 3740 3703
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3712 2990 3740 3334
rect 3804 3194 3832 4490
rect 3896 4026 3924 6054
rect 3988 5930 4016 7142
rect 4080 7002 4108 7822
rect 4632 7750 4660 8978
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7449 4660 7686
rect 4618 7440 4674 7449
rect 4618 7375 4674 7384
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6254 4384 6598
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 3988 5914 4200 5930
rect 3988 5908 4212 5914
rect 3988 5902 4160 5908
rect 4160 5850 4212 5856
rect 3988 5630 4200 5658
rect 4356 5642 4384 6190
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 3988 4214 4016 5630
rect 4172 5574 4200 5630
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4080 4826 4108 5510
rect 4356 5370 4384 5578
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4356 4282 4384 4490
rect 4724 4486 4752 5714
rect 4712 4480 4764 4486
rect 4710 4448 4712 4457
rect 4764 4448 4766 4457
rect 4710 4383 4766 4392
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4342 4040 4398 4049
rect 3896 3998 4016 4026
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3896 2650 3924 3878
rect 3988 2990 4016 3998
rect 4342 3975 4398 3984
rect 4250 3904 4306 3913
rect 4250 3839 4306 3848
rect 4264 3738 4292 3839
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4250 3632 4306 3641
rect 4356 3618 4384 3975
rect 4306 3590 4384 3618
rect 4250 3567 4306 3576
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4066 2952 4122 2961
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3988 2530 4016 2926
rect 4066 2887 4122 2896
rect 3712 2502 4016 2530
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 3146 1864 3202 1873
rect 3146 1799 3202 1808
rect 3160 480 3188 1799
rect 3712 480 3740 2502
rect 4080 1057 4108 2887
rect 4066 1048 4122 1057
rect 4066 983 4122 992
rect 4264 480 4292 3567
rect 4816 480 4844 10911
rect 5000 10470 5028 11154
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5184 9704 5212 12378
rect 5368 10033 5396 13767
rect 5448 13738 5500 13744
rect 5460 13530 5488 13738
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5552 13462 5580 13942
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5460 12442 5488 13330
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6564 12458 6592 13670
rect 6656 13462 6684 15030
rect 6840 15026 6960 15042
rect 6828 15020 6960 15026
rect 6880 15014 6960 15020
rect 6828 14962 6880 14968
rect 6840 14906 6868 14962
rect 6748 14878 6868 14906
rect 6748 14482 6776 14878
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6748 14006 6776 14418
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13462 6960 13670
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6656 12889 6684 13398
rect 6642 12880 6698 12889
rect 6642 12815 6698 12824
rect 5448 12436 5500 12442
rect 6564 12430 6684 12458
rect 5448 12378 5500 12384
rect 6656 12356 6684 12430
rect 6564 12328 6684 12356
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 10674 5488 11018
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 6090 10568 6146 10577
rect 6090 10503 6146 10512
rect 5448 10464 5500 10470
rect 5500 10424 5580 10452
rect 5448 10406 5500 10412
rect 5354 10024 5410 10033
rect 5354 9959 5410 9968
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5184 9676 5304 9704
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5078 7984 5134 7993
rect 5184 7954 5212 8298
rect 5078 7919 5134 7928
rect 5172 7948 5224 7954
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7546 4936 7686
rect 5092 7546 5120 7919
rect 5172 7890 5224 7896
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7206 5212 7890
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 6798 5212 7142
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 6458 5212 6734
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4908 5302 4936 5850
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4908 4185 4936 5238
rect 5276 5148 5304 9676
rect 5368 9518 5396 9862
rect 5446 9616 5502 9625
rect 5552 9586 5580 10424
rect 6104 10266 6132 10503
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 5998 10024 6054 10033
rect 5998 9959 6054 9968
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5446 9551 5448 9560
rect 5500 9551 5502 9560
rect 5540 9580 5592 9586
rect 5448 9522 5500 9528
rect 5540 9522 5592 9528
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7954 5396 8230
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5368 7342 5396 7890
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5538 7304 5594 7313
rect 5538 7239 5594 7248
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 7002 5488 7142
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5552 6905 5580 7239
rect 5538 6896 5594 6905
rect 5448 6860 5500 6866
rect 5538 6831 5594 6840
rect 5448 6802 5500 6808
rect 5460 6746 5488 6802
rect 5368 6718 5488 6746
rect 5368 6118 5396 6718
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 5574 5396 6054
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5184 5120 5304 5148
rect 4986 4992 5042 5001
rect 4986 4927 5042 4936
rect 5000 4321 5028 4927
rect 5184 4706 5212 5120
rect 5354 4856 5410 4865
rect 5354 4791 5356 4800
rect 5408 4791 5410 4800
rect 5356 4762 5408 4768
rect 5184 4678 5396 4706
rect 4986 4312 5042 4321
rect 4986 4247 5042 4256
rect 4894 4176 4950 4185
rect 4894 4111 4950 4120
rect 4908 3194 4936 4111
rect 5000 3738 5028 4247
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5000 2922 5028 3674
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 5184 2650 5212 4082
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5368 480 5396 4678
rect 5460 4010 5488 5510
rect 5552 4162 5580 6831
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5630 4720 5686 4729
rect 5630 4655 5632 4664
rect 5684 4655 5686 4664
rect 5632 4626 5684 4632
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5552 4134 5764 4162
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5460 3738 5488 3946
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3738 5580 3878
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5552 3194 5580 3674
rect 5736 3670 5764 4134
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 480 6040 9959
rect 6104 9178 6132 10202
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6182 10024 6238 10033
rect 6182 9959 6238 9968
rect 6196 9586 6224 9959
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6380 9382 6408 10134
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6322 6316 6598
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 5778 6316 6258
rect 6380 6254 6408 9318
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6472 8090 6500 8774
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6472 5778 6500 6598
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6104 4826 6132 5510
rect 6288 5370 6316 5714
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6288 5098 6316 5306
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6472 4826 6500 5714
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6104 4282 6132 4762
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6196 4010 6224 4558
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6104 3233 6132 3538
rect 6090 3224 6146 3233
rect 6196 3194 6224 3606
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6090 3159 6146 3168
rect 6184 3188 6236 3194
rect 6104 2990 6132 3159
rect 6184 3130 6236 3136
rect 6380 3058 6408 3334
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6380 2553 6408 2994
rect 6366 2544 6422 2553
rect 6366 2479 6368 2488
rect 6420 2479 6422 2488
rect 6368 2450 6420 2456
rect 6564 480 6592 12328
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9382 6684 10066
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 5001 6684 9318
rect 6748 6905 6776 9658
rect 6840 7970 6868 9930
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9450 6960 9862
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6932 8838 6960 9386
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8090 6960 8298
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6840 7954 6960 7970
rect 6840 7948 6972 7954
rect 6840 7942 6920 7948
rect 6920 7890 6972 7896
rect 6920 7472 6972 7478
rect 6918 7440 6920 7449
rect 6972 7440 6974 7449
rect 6918 7375 6974 7384
rect 6734 6896 6790 6905
rect 6734 6831 6790 6840
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6932 6254 6960 6734
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7024 5778 7052 16759
rect 7472 16730 7524 16736
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7300 15910 7328 16594
rect 8114 16008 8170 16017
rect 8114 15943 8170 15952
rect 7288 15904 7340 15910
rect 7102 15872 7158 15881
rect 7288 15846 7340 15852
rect 7102 15807 7158 15816
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7010 5672 7066 5681
rect 7010 5607 7066 5616
rect 6826 5400 6882 5409
rect 6826 5335 6828 5344
rect 6880 5335 6882 5344
rect 6828 5306 6880 5312
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6642 4992 6698 5001
rect 6642 4927 6698 4936
rect 6748 3602 6776 5034
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4826 6868 4966
rect 7024 4826 7052 5607
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6932 3754 6960 3946
rect 7012 3936 7064 3942
rect 7010 3904 7012 3913
rect 7064 3904 7066 3913
rect 7010 3839 7066 3848
rect 6932 3726 7052 3754
rect 7024 3670 7052 3726
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3126 6776 3538
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6748 2650 6776 3062
rect 7024 2990 7052 3606
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6748 2514 6776 2586
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7116 480 7144 15807
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 9722 7236 14758
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9042 7236 9386
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7208 8294 7236 8978
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7002 7236 8230
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7208 6322 7236 6938
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 678 7236 5714
rect 7300 4842 7328 15846
rect 8128 15162 8156 15943
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7392 13530 7420 13874
rect 8220 13705 8248 18022
rect 9692 17785 9720 22607
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 12714 21448 12770 21457
rect 12714 21383 12770 21392
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 12070 20360 12126 20369
rect 12070 20295 12126 20304
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 12084 19310 12112 20295
rect 12728 19310 12756 21383
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9678 17776 9734 17785
rect 9678 17711 9734 17720
rect 8206 13696 8262 13705
rect 8206 13631 8262 13640
rect 9402 13696 9458 13705
rect 9402 13631 9458 13640
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 7746 11248 7802 11257
rect 7746 11183 7802 11192
rect 7760 10266 7788 11183
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7760 9722 7788 10202
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 9110 7420 9318
rect 8220 9194 8248 9862
rect 8220 9178 8340 9194
rect 8220 9172 8352 9178
rect 8220 9166 8300 9172
rect 8300 9114 8352 9120
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7392 8634 7420 9046
rect 8404 8906 8432 9930
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7562 7848 7618 7857
rect 7562 7783 7564 7792
rect 7616 7783 7618 7792
rect 7564 7754 7616 7760
rect 7668 7546 7696 8026
rect 8128 7886 8156 8570
rect 8404 8362 8432 8842
rect 8482 8664 8538 8673
rect 8482 8599 8538 8608
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8312 8022 8340 8230
rect 8404 8090 8432 8298
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7930 7712 7986 7721
rect 7930 7647 7986 7656
rect 7944 7546 7972 7647
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8128 7002 8156 7822
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7410 8432 7686
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 7002 8432 7346
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7760 5914 7788 6122
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7760 5370 7788 5850
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7852 5166 7880 6598
rect 8220 5574 8248 6870
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 6656 8352 6662
rect 8404 6633 8432 6734
rect 8300 6598 8352 6604
rect 8390 6624 8446 6633
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7300 4814 7696 4842
rect 7852 4826 7880 5102
rect 7196 672 7248 678
rect 7196 614 7248 620
rect 7668 480 7696 4814
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 4185 8064 4422
rect 8022 4176 8078 4185
rect 8022 4111 8078 4120
rect 8128 3942 8156 4694
rect 8208 4072 8260 4078
rect 8312 4026 8340 6598
rect 8390 6559 8446 6568
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8404 5137 8432 5510
rect 8496 5409 8524 8599
rect 8574 7440 8630 7449
rect 8574 7375 8576 7384
rect 8628 7375 8630 7384
rect 8576 7346 8628 7352
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8588 5914 8616 6734
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8680 5710 8708 6054
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8482 5400 8538 5409
rect 8482 5335 8538 5344
rect 8680 5166 8708 5646
rect 8668 5160 8720 5166
rect 8390 5128 8446 5137
rect 8390 5063 8446 5072
rect 8574 5128 8630 5137
rect 8668 5102 8720 5108
rect 8574 5063 8630 5072
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8404 4282 8432 4966
rect 8588 4758 8616 5063
rect 8680 4758 8708 5102
rect 8758 4856 8814 4865
rect 8758 4791 8814 4800
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8260 4020 8432 4026
rect 8208 4014 8432 4020
rect 8220 3998 8432 4014
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3777 8340 3878
rect 8298 3768 8354 3777
rect 8298 3703 8354 3712
rect 8114 3632 8170 3641
rect 8114 3567 8170 3576
rect 8128 3058 8156 3567
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8208 2984 8260 2990
rect 8260 2944 8340 2972
rect 8208 2926 8260 2932
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7760 2582 7788 2790
rect 8312 2650 8340 2944
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 8404 1737 8432 3998
rect 8496 3942 8524 4558
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8772 3097 8800 4791
rect 8758 3088 8814 3097
rect 8758 3023 8814 3032
rect 8390 1728 8446 1737
rect 8390 1663 8446 1672
rect 8208 604 8260 610
rect 8208 546 8260 552
rect 8220 480 8248 546
rect 8864 480 8892 11630
rect 9310 8120 9366 8129
rect 9310 8055 9366 8064
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 4826 8984 7686
rect 9324 7546 9352 8055
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9324 6798 9352 6829
rect 9312 6792 9364 6798
rect 9310 6760 9312 6769
rect 9364 6760 9366 6769
rect 9310 6695 9366 6704
rect 9324 6458 9352 6695
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9048 3738 9076 4014
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8942 3496 8998 3505
rect 8942 3431 8944 3440
rect 8996 3431 8998 3440
rect 8944 3402 8996 3408
rect 8956 2990 8984 3402
rect 9048 3194 9076 3674
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9416 480 9444 13631
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9600 8514 9628 9454
rect 9692 9178 9720 10406
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9770 9208 9826 9217
rect 9680 9172 9732 9178
rect 9770 9143 9826 9152
rect 9680 9114 9732 9120
rect 9784 9110 9812 9143
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9678 8936 9734 8945
rect 9678 8871 9680 8880
rect 9732 8871 9734 8880
rect 9680 8842 9732 8848
rect 9508 8090 9536 8502
rect 9600 8486 9720 8514
rect 9692 8344 9720 8486
rect 9600 8316 9720 8344
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9600 8022 9628 8316
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9692 7954 9720 8316
rect 9680 7948 9732 7954
rect 9732 7908 9812 7936
rect 9680 7890 9732 7896
rect 9784 7206 9812 7908
rect 9876 7342 9904 9998
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6934 9812 7142
rect 9772 6928 9824 6934
rect 9824 6888 9904 6916
rect 9772 6870 9824 6876
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9508 5914 9536 6666
rect 9692 6118 9720 6802
rect 9770 6624 9826 6633
rect 9770 6559 9826 6568
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9600 4758 9628 5578
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9692 4049 9720 6054
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 9692 3670 9720 3975
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 2650 9628 3470
rect 9692 3058 9720 3606
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9784 2854 9812 6559
rect 9876 6322 9904 6888
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9876 1601 9904 2450
rect 9862 1592 9918 1601
rect 9862 1527 9918 1536
rect 9968 480 9996 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10690 16688 10746 16697
rect 10690 16623 10746 16632
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10060 8974 10088 9386
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8566 10088 8910
rect 10152 8634 10180 9114
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10152 7410 10180 7958
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10232 5840 10284 5846
rect 10046 5808 10102 5817
rect 10232 5782 10284 5788
rect 10046 5743 10048 5752
rect 10100 5743 10102 5752
rect 10048 5714 10100 5720
rect 10060 5302 10088 5714
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 10138 5264 10194 5273
rect 10138 5199 10194 5208
rect 10048 5024 10100 5030
rect 10046 4992 10048 5001
rect 10100 4992 10102 5001
rect 10046 4927 10102 4936
rect 10152 4826 10180 5199
rect 10244 5098 10272 5782
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10048 4752 10100 4758
rect 10046 4720 10048 4729
rect 10100 4720 10102 4729
rect 10046 4655 10102 4664
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4078 10272 4558
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10428 3126 10456 3538
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10428 2961 10456 3062
rect 10414 2952 10470 2961
rect 10414 2887 10470 2896
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2632 10732 16623
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9518 11008 9998
rect 11072 9722 11100 10066
rect 11624 9926 11652 19246
rect 12622 17776 12678 17785
rect 12622 17711 12678 17720
rect 11702 16144 11758 16153
rect 11702 16079 11758 16088
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 9382 11008 9454
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11072 9178 11100 9658
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10980 8362 11008 9046
rect 11072 8498 11100 9114
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 11334 8120 11390 8129
rect 11334 8055 11390 8064
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7449 11100 7686
rect 11058 7440 11114 7449
rect 10968 7404 11020 7410
rect 11348 7410 11376 8055
rect 11716 7546 11744 16079
rect 12254 13832 12310 13841
rect 12254 13767 12310 13776
rect 12268 12306 12296 13767
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11558 12020 12174
rect 12268 11898 12296 12242
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 11891 9602 11919 9862
rect 11808 9574 11919 9602
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11058 7375 11114 7384
rect 11336 7404 11388 7410
rect 10968 7346 11020 7352
rect 11336 7346 11388 7352
rect 10980 7206 11008 7346
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 7041 11008 7142
rect 10966 7032 11022 7041
rect 10966 6967 11022 6976
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6186 10824 6666
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10796 5846 10824 6122
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10796 5370 10824 5782
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10888 4808 10916 6802
rect 10980 6798 11008 6967
rect 11058 6896 11114 6905
rect 11058 6831 11114 6840
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 5778 11008 6190
rect 11072 5794 11100 6831
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11164 5914 11192 6734
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 10968 5772 11020 5778
rect 11072 5766 11192 5794
rect 10968 5714 11020 5720
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11072 5370 11100 5578
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10796 4780 10916 4808
rect 10796 4049 10824 4780
rect 10888 4690 11100 4706
rect 10888 4684 11112 4690
rect 10888 4678 11060 4684
rect 10782 4040 10838 4049
rect 10782 3975 10838 3984
rect 10782 3904 10838 3913
rect 10782 3839 10838 3848
rect 10796 3738 10824 3839
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10796 2689 10824 2994
rect 10520 2604 10732 2632
rect 10782 2680 10838 2689
rect 10888 2650 10916 4678
rect 11060 4626 11112 4632
rect 10968 4616 11020 4622
rect 11164 4570 11192 5766
rect 11256 5137 11284 6598
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11348 5681 11376 6054
rect 11532 5846 11560 6394
rect 11624 6361 11652 6598
rect 11808 6440 11836 9574
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 8974 12204 9318
rect 12452 9110 12480 9862
rect 12530 9344 12586 9353
rect 12530 9279 12586 9288
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8498 12204 8910
rect 12452 8634 12480 9046
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12084 8090 12112 8298
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12164 7336 12216 7342
rect 12162 7304 12164 7313
rect 12216 7304 12218 7313
rect 12162 7239 12218 7248
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11716 6412 11836 6440
rect 11610 6352 11666 6361
rect 11610 6287 11666 6296
rect 11520 5840 11572 5846
rect 11440 5788 11520 5794
rect 11440 5782 11572 5788
rect 11440 5766 11560 5782
rect 11334 5672 11390 5681
rect 11334 5607 11390 5616
rect 11242 5128 11298 5137
rect 11242 5063 11298 5072
rect 11336 5024 11388 5030
rect 11334 4992 11336 5001
rect 11388 4992 11390 5001
rect 11334 4927 11390 4936
rect 11440 4826 11468 5766
rect 11518 5672 11574 5681
rect 11518 5607 11574 5616
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 10968 4558 11020 4564
rect 10980 3194 11008 4558
rect 11072 4542 11192 4570
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10782 2615 10838 2624
rect 10876 2644 10928 2650
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10428 2310 10456 2450
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10060 1465 10088 2246
rect 10428 1873 10456 2246
rect 10414 1864 10470 1873
rect 10414 1799 10470 1808
rect 10046 1456 10102 1465
rect 10046 1391 10102 1400
rect 10520 480 10548 2604
rect 10876 2586 10928 2592
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 2009 10824 2246
rect 10782 2000 10838 2009
rect 10782 1935 10838 1944
rect 11072 480 11100 4542
rect 11334 4176 11390 4185
rect 11334 4111 11390 4120
rect 11348 4078 11376 4111
rect 11336 4072 11388 4078
rect 11150 4040 11206 4049
rect 11336 4014 11388 4020
rect 11150 3975 11206 3984
rect 11164 3777 11192 3975
rect 11532 3942 11560 5607
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11150 3768 11206 3777
rect 11150 3703 11152 3712
rect 11204 3703 11206 3712
rect 11152 3674 11204 3680
rect 11164 3058 11192 3674
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3534 11560 3606
rect 11624 3602 11652 5306
rect 11716 5080 11744 6412
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11900 5370 11928 6190
rect 11992 6118 12020 6802
rect 12162 6216 12218 6225
rect 12162 6151 12218 6160
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 12176 5846 12204 6151
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11716 5052 11836 5080
rect 11808 4842 11836 5052
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11716 4814 11836 4842
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11532 3058 11560 3470
rect 11624 3194 11652 3538
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11532 2938 11560 2994
rect 11532 2910 11652 2938
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 1873 11192 2790
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11348 2281 11376 2450
rect 11624 2446 11652 2910
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11334 2272 11390 2281
rect 11334 2207 11390 2216
rect 11150 1864 11206 1873
rect 11150 1799 11206 1808
rect 11716 480 11744 4814
rect 12176 4690 12204 4966
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11992 3670 12020 4218
rect 12084 4214 12112 4558
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11980 3664 12032 3670
rect 12176 3641 12204 3878
rect 11980 3606 12032 3612
rect 12162 3632 12218 3641
rect 12162 3567 12218 3576
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 12084 2650 12112 2994
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12268 480 12296 7482
rect 12360 6780 12388 8366
rect 12452 8090 12480 8570
rect 12544 8294 12572 9279
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12544 7546 12572 7822
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12440 6792 12492 6798
rect 12360 6752 12440 6780
rect 12360 5522 12388 6752
rect 12440 6734 12492 6740
rect 12440 5568 12492 5574
rect 12360 5516 12440 5522
rect 12360 5510 12492 5516
rect 12360 5494 12480 5510
rect 12360 2378 12388 5494
rect 12636 2802 12664 17711
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 4282 12756 12038
rect 12806 11792 12862 11801
rect 12806 11727 12862 11736
rect 12820 7274 12848 11727
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 9636 13216 11494
rect 13096 9608 13216 9636
rect 13096 9382 13124 9608
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12912 8090 12940 8434
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12990 7440 13046 7449
rect 12990 7375 12992 7384
rect 13044 7375 13046 7384
rect 12992 7346 13044 7352
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12820 7002 12848 7210
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 13082 6896 13138 6905
rect 13082 6831 13084 6840
rect 13136 6831 13138 6840
rect 13084 6802 13136 6808
rect 13096 6254 13124 6802
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13096 5914 13124 6190
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13082 4584 13138 4593
rect 13082 4519 13084 4528
rect 13136 4519 13138 4528
rect 13084 4490 13136 4496
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12912 4146 12940 4422
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12912 3913 12940 4082
rect 12898 3904 12954 3913
rect 12898 3839 12954 3848
rect 13004 3738 13032 4150
rect 13280 3924 13308 19246
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13450 9616 13506 9625
rect 13450 9551 13506 9560
rect 13464 4978 13492 9551
rect 13556 9450 13584 9862
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13556 8838 13584 9386
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 7478 13584 8774
rect 13832 8090 13860 9998
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13726 7712 13782 7721
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13648 7313 13676 7686
rect 13726 7647 13782 7656
rect 13634 7304 13690 7313
rect 13634 7239 13690 7248
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13556 5846 13584 6802
rect 13636 6792 13688 6798
rect 13740 6769 13768 7647
rect 13832 7546 13860 8026
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13820 6792 13872 6798
rect 13636 6734 13688 6740
rect 13726 6760 13782 6769
rect 13648 5953 13676 6734
rect 13820 6734 13872 6740
rect 13726 6695 13782 6704
rect 13832 6458 13860 6734
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13818 6216 13874 6225
rect 13818 6151 13874 6160
rect 13832 6118 13860 6151
rect 13820 6112 13872 6118
rect 13740 6072 13820 6100
rect 13634 5944 13690 5953
rect 13634 5879 13690 5888
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13740 5098 13768 6072
rect 13820 6054 13872 6060
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13464 4950 13676 4978
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13372 4078 13400 4490
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13464 3942 13492 4626
rect 13556 4282 13584 4762
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13452 3936 13504 3942
rect 13280 3896 13400 3924
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13004 2990 13032 3674
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12636 2774 12756 2802
rect 12728 2666 12756 2774
rect 12728 2638 12848 2666
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12820 480 12848 2638
rect 13372 480 13400 3896
rect 13452 3878 13504 3884
rect 13464 3738 13492 3878
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13648 2310 13676 4950
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 4026 13768 4558
rect 13820 4072 13872 4078
rect 13740 4020 13820 4026
rect 13740 4014 13872 4020
rect 13740 3998 13860 4014
rect 13832 2854 13860 3998
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 2582 13860 2790
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13924 480 13952 23015
rect 14292 17270 14320 23559
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 24122 23352 24178 23361
rect 24122 23287 24178 23296
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 14554 18864 14610 18873
rect 14554 18799 14610 18808
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14094 11656 14150 11665
rect 14094 11591 14150 11600
rect 14002 10704 14058 10713
rect 14002 10639 14058 10648
rect 14016 5914 14044 10639
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14016 4078 14044 5850
rect 14108 4146 14136 11591
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 9178 14320 9318
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14186 8528 14242 8537
rect 14186 8463 14242 8472
rect 14200 5778 14228 8463
rect 14292 8430 14320 9114
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14292 7886 14320 8366
rect 14384 8294 14412 9454
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14384 7546 14412 8230
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14384 5817 14412 5850
rect 14370 5808 14426 5817
rect 14188 5772 14240 5778
rect 14370 5743 14426 5752
rect 14188 5714 14240 5720
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14200 3602 14228 4422
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 2961 14320 3334
rect 14278 2952 14334 2961
rect 14278 2887 14334 2896
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14292 2553 14320 2586
rect 14278 2544 14334 2553
rect 14278 2479 14334 2488
rect 14384 2281 14412 4014
rect 14462 3904 14518 3913
rect 14462 3839 14518 3848
rect 14476 3505 14504 3839
rect 14462 3496 14518 3505
rect 14462 3431 14518 3440
rect 14462 3224 14518 3233
rect 14462 3159 14518 3168
rect 14476 2825 14504 3159
rect 14462 2816 14518 2825
rect 14462 2751 14518 2760
rect 14370 2272 14426 2281
rect 14370 2207 14426 2216
rect 14568 480 14596 18799
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14660 4146 14688 4626
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14660 2009 14688 3946
rect 14646 2000 14702 2009
rect 14646 1935 14702 1944
rect 14752 1306 14780 17206
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 24136 16017 24164 23287
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24122 16008 24178 16017
rect 24122 15943 24178 15952
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15658 9480 15714 9489
rect 15658 9415 15714 9424
rect 15672 9178 15700 9415
rect 16960 9382 16988 9998
rect 17236 9722 17264 10066
rect 18326 10024 18382 10033
rect 18326 9959 18328 9968
rect 18380 9959 18382 9968
rect 18328 9930 18380 9936
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15672 8634 15700 9114
rect 16210 9072 16266 9081
rect 16120 9036 16172 9042
rect 16210 9007 16266 9016
rect 16120 8978 16172 8984
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14844 6662 14872 7210
rect 15304 7177 15332 7686
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15290 7168 15346 7177
rect 15290 7103 15346 7112
rect 15488 6934 15516 7482
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 5030 14872 6598
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15488 6322 15516 6870
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15488 5778 15516 6258
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15016 5704 15068 5710
rect 15014 5672 15016 5681
rect 15068 5672 15070 5681
rect 15014 5607 15070 5616
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 14844 4865 14872 4966
rect 14830 4856 14886 4865
rect 15304 4826 15332 4966
rect 14830 4791 14886 4800
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15028 3534 15056 4014
rect 15304 3738 15332 4762
rect 15580 4758 15608 8230
rect 15658 8120 15714 8129
rect 15658 8055 15660 8064
rect 15712 8055 15714 8064
rect 15660 8026 15712 8032
rect 15672 7478 15700 8026
rect 15856 8022 15884 8910
rect 16132 8362 16160 8978
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15764 7002 15792 7822
rect 15856 7546 15884 7958
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15948 7546 15976 7822
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15856 6746 15884 7482
rect 15948 6905 15976 7482
rect 15934 6896 15990 6905
rect 15934 6831 15990 6840
rect 15764 6718 15884 6746
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15764 6458 15792 6718
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15764 6254 15792 6394
rect 15856 6361 15884 6598
rect 15842 6352 15898 6361
rect 15842 6287 15898 6296
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15948 6118 15976 6734
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15580 4078 15608 4694
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15764 4282 15792 4558
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15750 4176 15806 4185
rect 15750 4111 15806 4120
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15580 3670 15608 4014
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15658 3632 15714 3641
rect 15476 3596 15528 3602
rect 15658 3567 15660 3576
rect 15476 3538 15528 3544
rect 15712 3567 15714 3576
rect 15660 3538 15712 3544
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15304 3097 15332 3334
rect 15396 3126 15424 3470
rect 15488 3369 15516 3538
rect 15474 3360 15530 3369
rect 15474 3295 15530 3304
rect 15672 3194 15700 3538
rect 15764 3233 15792 4111
rect 15856 4049 15884 5510
rect 15842 4040 15898 4049
rect 15842 3975 15898 3984
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15750 3224 15806 3233
rect 15660 3188 15712 3194
rect 15750 3159 15806 3168
rect 15660 3130 15712 3136
rect 15384 3120 15436 3126
rect 15290 3088 15346 3097
rect 15384 3062 15436 3068
rect 15290 3023 15346 3032
rect 15856 2922 15884 3470
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15948 2825 15976 6054
rect 16132 4690 16160 8298
rect 16224 7002 16252 9007
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16224 5914 16252 6938
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16212 5296 16264 5302
rect 16210 5264 16212 5273
rect 16264 5264 16266 5273
rect 16210 5199 16266 5208
rect 16500 5098 16528 8774
rect 16854 8528 16910 8537
rect 16854 8463 16910 8472
rect 16868 8430 16896 8463
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 17222 8256 17278 8265
rect 17222 8191 17278 8200
rect 17236 8090 17264 8191
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17236 7478 17264 8026
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17328 7546 17356 7822
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17224 7472 17276 7478
rect 17328 7449 17356 7482
rect 17224 7414 17276 7420
rect 17314 7440 17370 7449
rect 17314 7375 17370 7384
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 5166 16896 7142
rect 17420 7002 17448 7822
rect 17512 7342 17540 9318
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 16960 6225 16988 6938
rect 17408 6792 17460 6798
rect 17512 6780 17540 7278
rect 17460 6752 17540 6780
rect 17408 6734 17460 6740
rect 16946 6216 17002 6225
rect 16946 6151 17002 6160
rect 17512 6118 17540 6752
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 16960 5846 16988 6054
rect 17314 5944 17370 5953
rect 17314 5879 17370 5888
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16960 5234 16988 5782
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16500 4826 16528 5034
rect 16960 4826 16988 5170
rect 17328 4826 17356 5879
rect 17512 5778 17540 6054
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 5370 17540 5714
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17776 5024 17828 5030
rect 17774 4992 17776 5001
rect 17828 4992 17830 5001
rect 17774 4927 17830 4936
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 16854 4720 16910 4729
rect 16120 4684 16172 4690
rect 16854 4655 16910 4664
rect 17224 4684 17276 4690
rect 16120 4626 16172 4632
rect 16868 4554 16896 4655
rect 17224 4626 17276 4632
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 17236 4146 17264 4626
rect 17328 4282 17356 4762
rect 17880 4672 17908 8502
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17972 5846 18000 7754
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 7342 18092 7686
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18064 5914 18092 6802
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18142 5808 18198 5817
rect 18142 5743 18198 5752
rect 18050 5128 18106 5137
rect 18050 5063 18106 5072
rect 18064 5030 18092 5063
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17958 4856 18014 4865
rect 17958 4791 17960 4800
rect 18012 4791 18014 4800
rect 17960 4762 18012 4768
rect 17960 4684 18012 4690
rect 17880 4644 17960 4672
rect 17960 4626 18012 4632
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17406 4040 17462 4049
rect 17406 3975 17462 3984
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16408 3534 16436 3878
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16776 3398 16804 3538
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 16776 3194 16804 3334
rect 17236 3194 17264 3334
rect 16764 3188 16816 3194
rect 17224 3188 17276 3194
rect 16816 3148 16896 3176
rect 16764 3130 16816 3136
rect 16762 2952 16818 2961
rect 16762 2887 16818 2896
rect 15934 2816 15990 2825
rect 15934 2751 15990 2760
rect 16210 2816 16266 2825
rect 16210 2751 16266 2760
rect 16394 2816 16450 2825
rect 16394 2751 16450 2760
rect 16224 2650 16252 2751
rect 16408 2650 16436 2751
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15856 2310 15884 2450
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14752 1278 15148 1306
rect 15120 480 15148 1278
rect 15672 480 15700 2246
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3146 0 3202 480
rect 3698 0 3754 480
rect 4250 0 4306 480
rect 4802 0 4858 480
rect 5354 0 5410 480
rect 5998 0 6054 480
rect 6550 0 6606 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8206 0 8262 480
rect 8850 0 8906 480
rect 9402 0 9458 480
rect 9954 0 10010 480
rect 10506 0 10562 480
rect 11058 0 11114 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 15856 105 15884 2246
rect 16210 1456 16266 1465
rect 16210 1391 16266 1400
rect 16224 480 16252 1391
rect 16776 480 16804 2887
rect 16868 2446 16896 3148
rect 17224 3130 17276 3136
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17420 480 17448 3975
rect 17696 3942 17724 4558
rect 18156 4078 18184 5743
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 17684 3936 17736 3942
rect 17682 3904 17684 3913
rect 17960 3936 18012 3942
rect 17736 3904 17738 3913
rect 17960 3878 18012 3884
rect 17682 3839 17738 3848
rect 17682 2408 17738 2417
rect 17682 2343 17684 2352
rect 17736 2343 17738 2352
rect 17684 2314 17736 2320
rect 17972 480 18000 3878
rect 18248 3738 18276 9590
rect 22190 9480 22246 9489
rect 22190 9415 22246 9424
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 22204 9042 22232 9415
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 21638 8936 21694 8945
rect 21638 8871 21694 8880
rect 21652 8430 21680 8871
rect 22204 8634 22232 8978
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20534 7984 20590 7993
rect 22112 7954 22140 8502
rect 20534 7919 20590 7928
rect 21088 7948 21140 7954
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18432 6254 18460 7822
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 7274 18920 7686
rect 20548 7342 20576 7919
rect 21088 7890 21140 7896
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 21100 7857 21128 7890
rect 21086 7848 21142 7857
rect 21086 7783 21142 7792
rect 21100 7546 21128 7783
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18892 7002 18920 7210
rect 19432 7200 19484 7206
rect 19154 7168 19210 7177
rect 19432 7142 19484 7148
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 19154 7103 19210 7112
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18892 6458 18920 6938
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18510 6352 18566 6361
rect 18510 6287 18512 6296
rect 18564 6287 18566 6296
rect 18512 6258 18564 6264
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18340 5817 18368 6122
rect 18512 5840 18564 5846
rect 18326 5808 18382 5817
rect 18512 5782 18564 5788
rect 18326 5743 18382 5752
rect 18524 5166 18552 5782
rect 19168 5778 19196 7103
rect 19444 7041 19472 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19430 7032 19486 7041
rect 19622 7024 19918 7044
rect 19430 6967 19486 6976
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19996 6254 20024 6695
rect 20732 6254 20760 7142
rect 22112 6866 22140 7686
rect 22756 7546 22784 7890
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 21270 6488 21326 6497
rect 21270 6423 21326 6432
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19168 5370 19196 5714
rect 19260 5681 19288 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20180 5778 20208 6054
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 19246 5672 19302 5681
rect 19246 5607 19302 5616
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18616 4826 18644 5170
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 19352 4690 19380 5510
rect 19430 5400 19486 5409
rect 20916 5370 20944 5714
rect 21086 5672 21142 5681
rect 21086 5607 21142 5616
rect 19430 5335 19486 5344
rect 20904 5364 20956 5370
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 18616 4282 18644 4626
rect 19352 4282 19380 4626
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19246 3904 19302 3913
rect 19246 3839 19302 3848
rect 19260 3738 19288 3839
rect 19338 3768 19394 3777
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 19248 3732 19300 3738
rect 19338 3703 19394 3712
rect 19248 3674 19300 3680
rect 18248 3058 18276 3674
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18420 2916 18472 2922
rect 18420 2858 18472 2864
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18050 2680 18106 2689
rect 18050 2615 18052 2624
rect 18104 2615 18106 2624
rect 18052 2586 18104 2592
rect 18248 2417 18276 2790
rect 18432 2553 18460 2858
rect 18524 2854 18552 3334
rect 18512 2848 18564 2854
rect 18510 2816 18512 2825
rect 18564 2816 18566 2825
rect 18510 2751 18566 2760
rect 18418 2544 18474 2553
rect 18418 2479 18474 2488
rect 18234 2408 18290 2417
rect 18234 2343 18290 2352
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18340 1737 18368 2246
rect 18326 1728 18382 1737
rect 18326 1663 18382 1672
rect 18524 480 18552 2246
rect 19076 480 19104 3334
rect 19260 2446 19288 3674
rect 19352 2990 19380 3703
rect 19444 3194 19472 5335
rect 20904 5306 20956 5312
rect 20902 5264 20958 5273
rect 20902 5199 20958 5208
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19444 1873 19472 2858
rect 19430 1864 19486 1873
rect 19430 1799 19486 1808
rect 19536 1442 19564 4422
rect 20180 4185 20208 4966
rect 20916 4690 20944 5199
rect 21100 5166 21128 5607
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 20904 4684 20956 4690
rect 20956 4644 21036 4672
rect 20904 4626 20956 4632
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20166 4176 20222 4185
rect 20166 4111 20222 4120
rect 19798 4040 19854 4049
rect 19798 3975 19800 3984
rect 19852 3975 19854 3984
rect 19800 3946 19852 3952
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20180 3058 20208 3674
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20076 2984 20128 2990
rect 20074 2952 20076 2961
rect 20128 2952 20130 2961
rect 20074 2887 20130 2896
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20088 2650 20116 2887
rect 20180 2650 20208 2994
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19904 2009 19932 2450
rect 19890 2000 19946 2009
rect 19890 1935 19946 1944
rect 19536 1414 19656 1442
rect 19628 480 19656 1414
rect 20272 480 20300 3878
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20640 3194 20668 3538
rect 20718 3360 20774 3369
rect 20718 3295 20774 3304
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20732 3126 20760 3295
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20824 480 20852 4422
rect 21008 3738 21036 4644
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 21100 4282 21128 4422
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 20904 3664 20956 3670
rect 20902 3632 20904 3641
rect 20956 3632 20958 3641
rect 20902 3567 20958 3576
rect 21086 3496 21142 3505
rect 21086 3431 21142 3440
rect 21100 2990 21128 3431
rect 21192 3369 21220 5510
rect 21284 4690 21312 6423
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21270 3496 21326 3505
rect 21270 3431 21326 3440
rect 21178 3360 21234 3369
rect 21178 3295 21234 3304
rect 21284 3233 21312 3431
rect 21270 3224 21326 3233
rect 21270 3159 21326 3168
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 21180 2576 21232 2582
rect 21178 2544 21180 2553
rect 21232 2544 21234 2553
rect 21178 2479 21234 2488
rect 21376 480 21404 3878
rect 21560 610 21588 3878
rect 21928 3233 21956 6054
rect 22100 5160 22152 5166
rect 22098 5128 22100 5137
rect 22152 5128 22154 5137
rect 22098 5063 22154 5072
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 22020 4282 22048 4626
rect 22190 4584 22246 4593
rect 22190 4519 22246 4528
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22112 4049 22140 4422
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 21914 3224 21970 3233
rect 21914 3159 21970 3168
rect 22204 2990 22232 4519
rect 22296 4010 22324 4966
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22388 3777 22416 6598
rect 22572 6458 22600 6802
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22558 4176 22614 4185
rect 22558 4111 22614 4120
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22374 3768 22430 3777
rect 22374 3703 22430 3712
rect 22480 3505 22508 4014
rect 22466 3496 22522 3505
rect 22466 3431 22522 3440
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22388 1601 22416 2790
rect 22572 2530 22600 4111
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22664 3194 22692 3878
rect 22940 3641 22968 7686
rect 23492 7342 23520 8774
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 23860 7478 23888 7890
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23480 7336 23532 7342
rect 23860 7313 23888 7414
rect 23480 7278 23532 7284
rect 23846 7304 23902 7313
rect 23846 7239 23902 7248
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 23860 3913 23888 7142
rect 24044 6866 24072 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24044 6458 24072 6802
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24136 4049 24164 6598
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24674 5808 24730 5817
rect 24674 5743 24730 5752
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 4729 24716 5743
rect 24674 4720 24730 4729
rect 24674 4655 24730 4664
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24122 4040 24178 4049
rect 24122 3975 24178 3984
rect 25962 4040 26018 4049
rect 25962 3975 26018 3984
rect 23846 3904 23902 3913
rect 23846 3839 23902 3848
rect 25318 3904 25374 3913
rect 25318 3839 25374 3848
rect 24214 3768 24270 3777
rect 24214 3703 24270 3712
rect 22926 3632 22982 3641
rect 22926 3567 22982 3576
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23110 3360 23166 3369
rect 23110 3295 23166 3304
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22480 2502 22600 2530
rect 22928 2508 22980 2514
rect 22374 1592 22430 1601
rect 22374 1527 22430 1536
rect 21548 604 21600 610
rect 21548 546 21600 552
rect 21916 604 21968 610
rect 21916 546 21968 552
rect 21928 480 21956 546
rect 22480 480 22508 2502
rect 22928 2450 22980 2456
rect 22940 2417 22968 2450
rect 22926 2408 22982 2417
rect 22926 2343 22982 2352
rect 23124 480 23152 3295
rect 23308 3126 23336 3538
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23296 3120 23348 3126
rect 23294 3088 23296 3097
rect 23348 3088 23350 3097
rect 23294 3023 23350 3032
rect 23492 2990 23520 3334
rect 23662 3224 23718 3233
rect 23662 3159 23718 3168
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23676 480 23704 3159
rect 24228 480 24256 3703
rect 24674 3632 24730 3641
rect 24674 3567 24730 3576
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24582 2952 24638 2961
rect 24582 2887 24638 2896
rect 24596 2854 24624 2887
rect 24584 2848 24636 2854
rect 24584 2790 24636 2796
rect 24688 2530 24716 3567
rect 24766 2816 24822 2825
rect 24766 2751 24822 2760
rect 24780 2650 24808 2751
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24688 2502 24808 2530
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24780 480 24808 2502
rect 25332 480 25360 3839
rect 25976 480 26004 3975
rect 27618 3088 27674 3097
rect 27618 3023 27674 3032
rect 26514 2952 26570 2961
rect 26514 2887 26570 2896
rect 26528 480 26556 2887
rect 27066 2816 27122 2825
rect 27066 2751 27122 2760
rect 27080 480 27108 2751
rect 27632 480 27660 3023
rect 15842 96 15898 105
rect 15842 31 15898 40
rect 16210 0 16266 480
rect 16762 0 16818 480
rect 17406 0 17462 480
rect 17958 0 18014 480
rect 18510 0 18566 480
rect 19062 0 19118 480
rect 19614 0 19670 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
rect 23110 0 23166 480
rect 23662 0 23718 480
rect 24214 0 24270 480
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3330 27512 3386 27568
rect 2686 26832 2742 26888
rect 1582 26152 1638 26208
rect 1490 25472 1546 25528
rect 1398 24792 1454 24848
rect 1674 24112 1730 24168
rect 1582 23432 1638 23488
rect 1490 22752 1546 22808
rect 1398 22072 1454 22128
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 3146 23588 3202 23624
rect 3146 23568 3148 23588
rect 3148 23568 3200 23588
rect 3200 23568 3202 23588
rect 2042 23024 2098 23080
rect 2042 22636 2098 22672
rect 2042 22616 2044 22636
rect 2044 22616 2096 22636
rect 2096 22616 2098 22636
rect 1582 21392 1638 21448
rect 2410 21392 2466 21448
rect 1674 20340 1676 20360
rect 1676 20340 1728 20360
rect 1728 20340 1730 20360
rect 1674 20304 1730 20340
rect 1582 19352 1638 19408
rect 1490 18672 1546 18728
rect 1674 19116 1676 19136
rect 1676 19116 1728 19136
rect 1728 19116 1730 19136
rect 1674 19080 1730 19116
rect 1582 16632 1638 16688
rect 1490 15952 1546 16008
rect 1398 14592 1454 14648
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 4066 20712 4122 20768
rect 3330 20032 3386 20088
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4066 19216 4122 19272
rect 3330 18944 3386 19000
rect 2502 18808 2558 18864
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 2042 16768 2098 16824
rect 1674 16088 1730 16144
rect 1582 15272 1638 15328
rect 1582 13912 1638 13968
rect 2042 13776 2098 13832
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5446 17312 5502 17368
rect 3054 16904 3110 16960
rect 5722 16904 5778 16960
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5906 15972 5962 16008
rect 5906 15952 5908 15972
rect 5908 15952 5960 15972
rect 5960 15952 5962 15972
rect 5170 15852 5172 15872
rect 5172 15852 5224 15872
rect 5224 15852 5226 15872
rect 5170 15816 5226 15852
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 14278 23568 14334 23624
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 13910 23024 13966 23080
rect 9678 22616 9734 22672
rect 8298 19216 8354 19272
rect 6734 19080 6790 19136
rect 7746 18944 7802 19000
rect 7470 17856 7526 17912
rect 7010 16768 7066 16824
rect 6734 16632 6790 16688
rect 6366 15952 6422 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5354 13776 5410 13832
rect 3146 13232 3202 13288
rect 3422 12552 3478 12608
rect 4158 12824 4214 12880
rect 3974 11872 4030 11928
rect 3422 11736 3478 11792
rect 3146 11600 3202 11656
rect 1674 10920 1730 10976
rect 2410 10648 2466 10704
rect 1214 9016 1270 9072
rect 1214 8472 1270 8528
rect 1398 8508 1400 8528
rect 1400 8508 1452 8528
rect 1452 8508 1454 8528
rect 1398 8472 1454 8508
rect 1398 4256 1454 4312
rect 1766 4120 1822 4176
rect 1582 3032 1638 3088
rect 3514 9832 3570 9888
rect 2502 6840 2558 6896
rect 2410 4548 2466 4584
rect 2410 4528 2412 4548
rect 2412 4528 2464 4548
rect 2464 4528 2466 4548
rect 2318 3712 2374 3768
rect 1950 1944 2006 2000
rect 2226 1672 2282 1728
rect 2686 4664 2742 4720
rect 3238 6704 3294 6760
rect 3698 9424 3754 9480
rect 4802 10920 4858 10976
rect 3790 9152 3846 9208
rect 3974 9152 4030 9208
rect 3882 8200 3938 8256
rect 3790 8064 3846 8120
rect 3698 7792 3754 7848
rect 3882 7112 3938 7168
rect 3698 3712 3754 3768
rect 3330 3576 3386 3632
rect 4618 7384 4674 7440
rect 4710 4428 4712 4448
rect 4712 4428 4764 4448
rect 4764 4428 4766 4448
rect 4710 4392 4766 4428
rect 4342 3984 4398 4040
rect 4250 3848 4306 3904
rect 4250 3576 4306 3632
rect 4066 2896 4122 2952
rect 3146 1808 3202 1864
rect 4066 992 4122 1048
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6642 12824 6698 12880
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6090 10512 6146 10568
rect 5354 9968 5410 10024
rect 5078 7928 5134 7984
rect 5446 9580 5502 9616
rect 5998 9968 6054 10024
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5446 9560 5448 9580
rect 5448 9560 5500 9580
rect 5500 9560 5502 9580
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5538 7248 5594 7304
rect 5538 6840 5594 6896
rect 4986 4936 5042 4992
rect 5354 4820 5410 4856
rect 5354 4800 5356 4820
rect 5356 4800 5408 4820
rect 5408 4800 5410 4820
rect 4986 4256 5042 4312
rect 4894 4120 4950 4176
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5630 4684 5686 4720
rect 5630 4664 5632 4684
rect 5632 4664 5684 4684
rect 5684 4664 5686 4684
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6182 9968 6238 10024
rect 6090 3168 6146 3224
rect 6366 2508 6422 2544
rect 6366 2488 6368 2508
rect 6368 2488 6420 2508
rect 6420 2488 6422 2508
rect 6918 7420 6920 7440
rect 6920 7420 6972 7440
rect 6972 7420 6974 7440
rect 6918 7384 6974 7420
rect 6734 6840 6790 6896
rect 8114 15952 8170 16008
rect 7102 15816 7158 15872
rect 7010 5616 7066 5672
rect 6826 5364 6882 5400
rect 6826 5344 6828 5364
rect 6828 5344 6880 5364
rect 6880 5344 6882 5364
rect 6642 4936 6698 4992
rect 7010 3884 7012 3904
rect 7012 3884 7064 3904
rect 7064 3884 7066 3904
rect 7010 3848 7066 3884
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 12714 21392 12770 21448
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 12070 20304 12126 20360
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9678 17720 9734 17776
rect 8206 13640 8262 13696
rect 9402 13640 9458 13696
rect 7746 11192 7802 11248
rect 7562 7812 7618 7848
rect 7562 7792 7564 7812
rect 7564 7792 7616 7812
rect 7616 7792 7618 7812
rect 8482 8608 8538 8664
rect 7930 7656 7986 7712
rect 8022 4120 8078 4176
rect 8390 6568 8446 6624
rect 8574 7404 8630 7440
rect 8574 7384 8576 7404
rect 8576 7384 8628 7404
rect 8628 7384 8630 7404
rect 8482 5344 8538 5400
rect 8390 5072 8446 5128
rect 8574 5072 8630 5128
rect 8758 4800 8814 4856
rect 8298 3712 8354 3768
rect 8114 3576 8170 3632
rect 8758 3032 8814 3088
rect 8390 1672 8446 1728
rect 9310 8064 9366 8120
rect 9310 6740 9312 6760
rect 9312 6740 9364 6760
rect 9364 6740 9366 6760
rect 9310 6704 9366 6740
rect 8942 3460 8998 3496
rect 8942 3440 8944 3460
rect 8944 3440 8996 3460
rect 8996 3440 8998 3460
rect 9770 9152 9826 9208
rect 9678 8900 9734 8936
rect 9678 8880 9680 8900
rect 9680 8880 9732 8900
rect 9732 8880 9734 8900
rect 9770 6568 9826 6624
rect 9678 3984 9734 4040
rect 9862 1536 9918 1592
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 16632 10746 16688
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10046 5772 10102 5808
rect 10046 5752 10048 5772
rect 10048 5752 10100 5772
rect 10100 5752 10102 5772
rect 10138 5208 10194 5264
rect 10046 4972 10048 4992
rect 10048 4972 10100 4992
rect 10100 4972 10102 4992
rect 10046 4936 10102 4972
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10046 4700 10048 4720
rect 10048 4700 10100 4720
rect 10100 4700 10102 4720
rect 10046 4664 10102 4700
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10414 2896 10470 2952
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12622 17720 12678 17776
rect 11702 16088 11758 16144
rect 11334 8064 11390 8120
rect 11058 7384 11114 7440
rect 12254 13776 12310 13832
rect 10966 6976 11022 7032
rect 11058 6840 11114 6896
rect 10782 3984 10838 4040
rect 10782 3848 10838 3904
rect 10782 2624 10838 2680
rect 12530 9288 12586 9344
rect 12162 7284 12164 7304
rect 12164 7284 12216 7304
rect 12216 7284 12218 7304
rect 12162 7248 12218 7284
rect 11610 6296 11666 6352
rect 11334 5616 11390 5672
rect 11242 5072 11298 5128
rect 11334 4972 11336 4992
rect 11336 4972 11388 4992
rect 11388 4972 11390 4992
rect 11334 4936 11390 4972
rect 11518 5616 11574 5672
rect 10414 1808 10470 1864
rect 10046 1400 10102 1456
rect 10782 1944 10838 2000
rect 11334 4120 11390 4176
rect 11150 3984 11206 4040
rect 11150 3732 11206 3768
rect 11150 3712 11152 3732
rect 11152 3712 11204 3732
rect 11204 3712 11206 3732
rect 12162 6160 12218 6216
rect 11334 2216 11390 2272
rect 11150 1808 11206 1864
rect 12162 3576 12218 3632
rect 12806 11736 12862 11792
rect 12990 7404 13046 7440
rect 12990 7384 12992 7404
rect 12992 7384 13044 7404
rect 13044 7384 13046 7404
rect 13082 6860 13138 6896
rect 13082 6840 13084 6860
rect 13084 6840 13136 6860
rect 13136 6840 13138 6860
rect 13082 4548 13138 4584
rect 13082 4528 13084 4548
rect 13084 4528 13136 4548
rect 13136 4528 13138 4548
rect 12898 3848 12954 3904
rect 13450 9560 13506 9616
rect 13726 7656 13782 7712
rect 13634 7248 13690 7304
rect 13726 6704 13782 6760
rect 13818 6160 13874 6216
rect 13634 5888 13690 5944
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 24122 23296 24178 23352
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 14554 18808 14610 18864
rect 14094 11600 14150 11656
rect 14002 10648 14058 10704
rect 14186 8472 14242 8528
rect 14370 5752 14426 5808
rect 14278 2896 14334 2952
rect 14278 2488 14334 2544
rect 14462 3848 14518 3904
rect 14462 3440 14518 3496
rect 14462 3168 14518 3224
rect 14462 2760 14518 2816
rect 14370 2216 14426 2272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14646 1944 14702 2000
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24122 15952 24178 16008
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15658 9424 15714 9480
rect 18326 9988 18382 10024
rect 18326 9968 18328 9988
rect 18328 9968 18380 9988
rect 18380 9968 18382 9988
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 16210 9016 16266 9072
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15290 7112 15346 7168
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15014 5652 15016 5672
rect 15016 5652 15068 5672
rect 15068 5652 15070 5672
rect 15014 5616 15070 5652
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14830 4800 14886 4856
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15658 8084 15714 8120
rect 15658 8064 15660 8084
rect 15660 8064 15712 8084
rect 15712 8064 15714 8084
rect 15934 6840 15990 6896
rect 15842 6296 15898 6352
rect 15750 4120 15806 4176
rect 15658 3596 15714 3632
rect 15658 3576 15660 3596
rect 15660 3576 15712 3596
rect 15712 3576 15714 3596
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15474 3304 15530 3360
rect 15842 3984 15898 4040
rect 15750 3168 15806 3224
rect 15290 3032 15346 3088
rect 16210 5244 16212 5264
rect 16212 5244 16264 5264
rect 16264 5244 16266 5264
rect 16210 5208 16266 5244
rect 16854 8472 16910 8528
rect 17222 8200 17278 8256
rect 17314 7384 17370 7440
rect 16946 6160 17002 6216
rect 17314 5888 17370 5944
rect 17774 4972 17776 4992
rect 17776 4972 17828 4992
rect 17828 4972 17830 4992
rect 17774 4936 17830 4972
rect 16854 4664 16910 4720
rect 18142 5752 18198 5808
rect 18050 5072 18106 5128
rect 17958 4820 18014 4856
rect 17958 4800 17960 4820
rect 17960 4800 18012 4820
rect 18012 4800 18014 4820
rect 17406 3984 17462 4040
rect 16762 2896 16818 2952
rect 15934 2760 15990 2816
rect 16210 2760 16266 2816
rect 16394 2760 16450 2816
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16210 1400 16266 1456
rect 17682 3884 17684 3904
rect 17684 3884 17736 3904
rect 17736 3884 17738 3904
rect 17682 3848 17738 3884
rect 17682 2372 17738 2408
rect 17682 2352 17684 2372
rect 17684 2352 17736 2372
rect 17736 2352 17738 2372
rect 22190 9424 22246 9480
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 21638 8880 21694 8936
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 20534 7928 20590 7984
rect 21086 7792 21142 7848
rect 19154 7112 19210 7168
rect 18510 6316 18566 6352
rect 18510 6296 18512 6316
rect 18512 6296 18564 6316
rect 18564 6296 18566 6316
rect 18326 5752 18382 5808
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19430 6976 19486 7032
rect 19982 6704 20038 6760
rect 21270 6432 21326 6488
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19246 5616 19302 5672
rect 19430 5344 19486 5400
rect 21086 5616 21142 5672
rect 19246 3848 19302 3904
rect 19338 3712 19394 3768
rect 18050 2644 18106 2680
rect 18050 2624 18052 2644
rect 18052 2624 18104 2644
rect 18104 2624 18106 2644
rect 18510 2796 18512 2816
rect 18512 2796 18564 2816
rect 18564 2796 18566 2816
rect 18510 2760 18566 2796
rect 18418 2488 18474 2544
rect 18234 2352 18290 2408
rect 18326 1672 18382 1728
rect 20902 5208 20958 5264
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19430 1808 19486 1864
rect 20166 4120 20222 4176
rect 19798 4004 19854 4040
rect 19798 3984 19800 4004
rect 19800 3984 19852 4004
rect 19852 3984 19854 4004
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20074 2932 20076 2952
rect 20076 2932 20128 2952
rect 20128 2932 20130 2952
rect 20074 2896 20130 2932
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19890 1944 19946 2000
rect 20718 3304 20774 3360
rect 20902 3612 20904 3632
rect 20904 3612 20956 3632
rect 20956 3612 20958 3632
rect 20902 3576 20958 3612
rect 21086 3440 21142 3496
rect 21270 3440 21326 3496
rect 21178 3304 21234 3360
rect 21270 3168 21326 3224
rect 21178 2524 21180 2544
rect 21180 2524 21232 2544
rect 21232 2524 21234 2544
rect 21178 2488 21234 2524
rect 22098 5108 22100 5128
rect 22100 5108 22152 5128
rect 22152 5108 22154 5128
rect 22098 5072 22154 5108
rect 22190 4528 22246 4584
rect 22098 3984 22154 4040
rect 21914 3168 21970 3224
rect 22558 4120 22614 4176
rect 22374 3712 22430 3768
rect 22466 3440 22522 3496
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 23846 7248 23902 7304
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24674 5752 24730 5808
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24674 4664 24730 4720
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24122 3984 24178 4040
rect 25962 3984 26018 4040
rect 23846 3848 23902 3904
rect 25318 3848 25374 3904
rect 24214 3712 24270 3768
rect 22926 3576 22982 3632
rect 23110 3304 23166 3360
rect 22374 1536 22430 1592
rect 22926 2352 22982 2408
rect 23294 3068 23296 3088
rect 23296 3068 23348 3088
rect 23348 3068 23350 3088
rect 23294 3032 23350 3068
rect 23662 3168 23718 3224
rect 24674 3576 24730 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24582 2896 24638 2952
rect 24766 2760 24822 2816
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27618 3032 27674 3088
rect 26514 2896 26570 2952
rect 27066 2760 27122 2816
rect 15842 40 15898 96
<< metal3 >>
rect 0 27570 480 27600
rect 3325 27570 3391 27573
rect 0 27568 3391 27570
rect 0 27512 3330 27568
rect 3386 27512 3391 27568
rect 0 27510 3391 27512
rect 0 27480 480 27510
rect 3325 27507 3391 27510
rect 0 26890 480 26920
rect 2681 26890 2747 26893
rect 0 26888 2747 26890
rect 0 26832 2686 26888
rect 2742 26832 2747 26888
rect 0 26830 2747 26832
rect 0 26800 480 26830
rect 2681 26827 2747 26830
rect 0 26210 480 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 0 26120 480 26150
rect 1577 26147 1643 26150
rect 10277 25600 10597 25601
rect 0 25530 480 25560
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1485 25530 1551 25533
rect 0 25528 1551 25530
rect 0 25472 1490 25528
rect 1546 25472 1551 25528
rect 0 25470 1551 25472
rect 0 25440 480 25470
rect 1485 25467 1551 25470
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 1393 24850 1459 24853
rect 0 24848 1459 24850
rect 0 24792 1398 24848
rect 1454 24792 1459 24848
rect 0 24790 1459 24792
rect 0 24760 480 24790
rect 1393 24787 1459 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24170 480 24200
rect 1669 24170 1735 24173
rect 0 24168 1735 24170
rect 0 24112 1674 24168
rect 1730 24112 1735 24168
rect 0 24110 1735 24112
rect 0 24080 480 24110
rect 1669 24107 1735 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 3141 23626 3207 23629
rect 14273 23626 14339 23629
rect 3141 23624 14339 23626
rect 3141 23568 3146 23624
rect 3202 23568 14278 23624
rect 14334 23568 14339 23624
rect 3141 23566 14339 23568
rect 3141 23563 3207 23566
rect 14273 23563 14339 23566
rect 0 23490 480 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 480 23430
rect 1577 23427 1643 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 24117 23354 24183 23357
rect 27520 23354 28000 23384
rect 24117 23352 28000 23354
rect 24117 23296 24122 23352
rect 24178 23296 28000 23352
rect 24117 23294 28000 23296
rect 24117 23291 24183 23294
rect 27520 23264 28000 23294
rect 2037 23082 2103 23085
rect 13905 23082 13971 23085
rect 2037 23080 13971 23082
rect 2037 23024 2042 23080
rect 2098 23024 13910 23080
rect 13966 23024 13971 23080
rect 2037 23022 13971 23024
rect 2037 23019 2103 23022
rect 13905 23019 13971 23022
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1485 22810 1551 22813
rect 0 22808 1551 22810
rect 0 22752 1490 22808
rect 1546 22752 1551 22808
rect 0 22750 1551 22752
rect 0 22720 480 22750
rect 1485 22747 1551 22750
rect 2037 22674 2103 22677
rect 9673 22674 9739 22677
rect 2037 22672 9739 22674
rect 2037 22616 2042 22672
rect 2098 22616 9678 22672
rect 9734 22616 9739 22672
rect 2037 22614 9739 22616
rect 2037 22611 2103 22614
rect 9673 22611 9739 22614
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 0 22130 480 22160
rect 1393 22130 1459 22133
rect 0 22128 1459 22130
rect 0 22072 1398 22128
rect 1454 22072 1459 22128
rect 0 22070 1459 22072
rect 0 22040 480 22070
rect 1393 22067 1459 22070
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21450 480 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 480 21390
rect 1577 21387 1643 21390
rect 2405 21450 2471 21453
rect 12709 21450 12775 21453
rect 2405 21448 12775 21450
rect 2405 21392 2410 21448
rect 2466 21392 12714 21448
rect 12770 21392 12775 21448
rect 2405 21390 12775 21392
rect 2405 21387 2471 21390
rect 12709 21387 12775 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 20770 480 20800
rect 4061 20770 4127 20773
rect 0 20768 4127 20770
rect 0 20712 4066 20768
rect 4122 20712 4127 20768
rect 0 20710 4127 20712
rect 0 20680 480 20710
rect 4061 20707 4127 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 1669 20362 1735 20365
rect 12065 20362 12131 20365
rect 1669 20360 12131 20362
rect 1669 20304 1674 20360
rect 1730 20304 12070 20360
rect 12126 20304 12131 20360
rect 1669 20302 12131 20304
rect 1669 20299 1735 20302
rect 12065 20299 12131 20302
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 3325 20090 3391 20093
rect 0 20088 3391 20090
rect 0 20032 3330 20088
rect 3386 20032 3391 20088
rect 0 20030 3391 20032
rect 0 20000 480 20030
rect 3325 20027 3391 20030
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19410 480 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 480 19350
rect 1577 19347 1643 19350
rect 4061 19274 4127 19277
rect 8293 19274 8359 19277
rect 4061 19272 8359 19274
rect 4061 19216 4066 19272
rect 4122 19216 8298 19272
rect 8354 19216 8359 19272
rect 4061 19214 8359 19216
rect 4061 19211 4127 19214
rect 8293 19211 8359 19214
rect 1669 19138 1735 19141
rect 6729 19138 6795 19141
rect 1669 19136 6795 19138
rect 1669 19080 1674 19136
rect 1730 19080 6734 19136
rect 6790 19080 6795 19136
rect 1669 19078 6795 19080
rect 1669 19075 1735 19078
rect 6729 19075 6795 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 3325 19002 3391 19005
rect 7741 19002 7807 19005
rect 3325 19000 7807 19002
rect 3325 18944 3330 19000
rect 3386 18944 7746 19000
rect 7802 18944 7807 19000
rect 3325 18942 7807 18944
rect 3325 18939 3391 18942
rect 7741 18939 7807 18942
rect 2497 18866 2563 18869
rect 14549 18866 14615 18869
rect 2497 18864 14615 18866
rect 2497 18808 2502 18864
rect 2558 18808 14554 18864
rect 14610 18808 14615 18864
rect 2497 18806 14615 18808
rect 2497 18803 2563 18806
rect 14549 18803 14615 18806
rect 0 18730 480 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 480 18670
rect 1485 18667 1551 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 0 18050 480 18080
rect 0 17990 3986 18050
rect 0 17960 480 17990
rect 3926 17914 3986 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 7465 17914 7531 17917
rect 3926 17912 7531 17914
rect 3926 17856 7470 17912
rect 7526 17856 7531 17912
rect 3926 17854 7531 17856
rect 7465 17851 7531 17854
rect 9673 17778 9739 17781
rect 12617 17778 12683 17781
rect 9673 17776 12683 17778
rect 9673 17720 9678 17776
rect 9734 17720 12622 17776
rect 12678 17720 12683 17776
rect 9673 17718 12683 17720
rect 9673 17715 9739 17718
rect 12617 17715 12683 17718
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 5441 17370 5507 17373
rect 0 17368 5507 17370
rect 0 17312 5446 17368
rect 5502 17312 5507 17368
rect 0 17310 5507 17312
rect 0 17280 480 17310
rect 5441 17307 5507 17310
rect 3049 16962 3115 16965
rect 5717 16962 5783 16965
rect 3049 16960 5783 16962
rect 3049 16904 3054 16960
rect 3110 16904 5722 16960
rect 5778 16904 5783 16960
rect 3049 16902 5783 16904
rect 3049 16899 3115 16902
rect 5717 16899 5783 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 2037 16826 2103 16829
rect 7005 16826 7071 16829
rect 2037 16824 7071 16826
rect 2037 16768 2042 16824
rect 2098 16768 7010 16824
rect 7066 16768 7071 16824
rect 2037 16766 7071 16768
rect 2037 16763 2103 16766
rect 7005 16763 7071 16766
rect 0 16690 480 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 480 16630
rect 1577 16627 1643 16630
rect 6729 16690 6795 16693
rect 10685 16690 10751 16693
rect 6729 16688 10751 16690
rect 6729 16632 6734 16688
rect 6790 16632 10690 16688
rect 10746 16632 10751 16688
rect 6729 16630 10751 16632
rect 6729 16627 6795 16630
rect 10685 16627 10751 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 1669 16146 1735 16149
rect 11697 16146 11763 16149
rect 1669 16144 11763 16146
rect 1669 16088 1674 16144
rect 1730 16088 11702 16144
rect 11758 16088 11763 16144
rect 1669 16086 11763 16088
rect 1669 16083 1735 16086
rect 11697 16083 11763 16086
rect 0 16010 480 16040
rect 1485 16010 1551 16013
rect 0 16008 1551 16010
rect 0 15952 1490 16008
rect 1546 15952 1551 16008
rect 0 15950 1551 15952
rect 0 15920 480 15950
rect 1485 15947 1551 15950
rect 5901 16010 5967 16013
rect 6361 16010 6427 16013
rect 8109 16010 8175 16013
rect 24117 16010 24183 16013
rect 5901 16008 24183 16010
rect 5901 15952 5906 16008
rect 5962 15952 6366 16008
rect 6422 15952 8114 16008
rect 8170 15952 24122 16008
rect 24178 15952 24183 16008
rect 5901 15950 24183 15952
rect 5901 15947 5967 15950
rect 6361 15947 6427 15950
rect 8109 15947 8175 15950
rect 24117 15947 24183 15950
rect 5165 15874 5231 15877
rect 7097 15874 7163 15877
rect 5165 15872 7163 15874
rect 5165 15816 5170 15872
rect 5226 15816 7102 15872
rect 7158 15816 7163 15872
rect 5165 15814 7163 15816
rect 5165 15811 5231 15814
rect 7097 15811 7163 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 0 15330 480 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 480 15270
rect 1577 15267 1643 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1393 14650 1459 14653
rect 0 14648 1459 14650
rect 0 14592 1398 14648
rect 1454 14592 1459 14648
rect 0 14590 1459 14592
rect 0 14560 480 14590
rect 1393 14587 1459 14590
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13970 480 14000
rect 1577 13970 1643 13973
rect 27520 13970 28000 14000
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 480 13910
rect 1577 13907 1643 13910
rect 27478 13880 28000 13970
rect 2037 13834 2103 13837
rect 5349 13834 5415 13837
rect 2037 13832 5415 13834
rect 2037 13776 2042 13832
rect 2098 13776 5354 13832
rect 5410 13776 5415 13832
rect 2037 13774 5415 13776
rect 2037 13771 2103 13774
rect 5349 13771 5415 13774
rect 12249 13834 12315 13837
rect 27478 13834 27538 13880
rect 12249 13832 27538 13834
rect 12249 13776 12254 13832
rect 12310 13776 27538 13832
rect 12249 13774 27538 13776
rect 12249 13771 12315 13774
rect 8201 13698 8267 13701
rect 9397 13698 9463 13701
rect 8201 13696 9463 13698
rect 8201 13640 8206 13696
rect 8262 13640 9402 13696
rect 9458 13640 9463 13696
rect 8201 13638 9463 13640
rect 8201 13635 8267 13638
rect 9397 13635 9463 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 0 13290 480 13320
rect 3141 13290 3207 13293
rect 0 13288 3207 13290
rect 0 13232 3146 13288
rect 3202 13232 3207 13288
rect 0 13230 3207 13232
rect 0 13200 480 13230
rect 3141 13227 3207 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 4153 12882 4219 12885
rect 6637 12882 6703 12885
rect 4153 12880 6703 12882
rect 4153 12824 4158 12880
rect 4214 12824 6642 12880
rect 6698 12824 6703 12880
rect 4153 12822 6703 12824
rect 4153 12819 4219 12822
rect 6637 12819 6703 12822
rect 0 12610 480 12640
rect 3417 12610 3483 12613
rect 0 12608 3483 12610
rect 0 12552 3422 12608
rect 3478 12552 3483 12608
rect 0 12550 3483 12552
rect 0 12520 480 12550
rect 3417 12547 3483 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 3969 11930 4035 11933
rect 0 11928 4035 11930
rect 0 11872 3974 11928
rect 4030 11872 4035 11928
rect 0 11870 4035 11872
rect 0 11840 480 11870
rect 3969 11867 4035 11870
rect 3417 11794 3483 11797
rect 12801 11794 12867 11797
rect 3417 11792 12867 11794
rect 3417 11736 3422 11792
rect 3478 11736 12806 11792
rect 12862 11736 12867 11792
rect 3417 11734 12867 11736
rect 3417 11731 3483 11734
rect 12801 11731 12867 11734
rect 3141 11658 3207 11661
rect 14089 11658 14155 11661
rect 3141 11656 14155 11658
rect 3141 11600 3146 11656
rect 3202 11600 14094 11656
rect 14150 11600 14155 11656
rect 3141 11598 14155 11600
rect 3141 11595 3207 11598
rect 14089 11595 14155 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 0 11250 480 11280
rect 7741 11250 7807 11253
rect 0 11248 7807 11250
rect 0 11192 7746 11248
rect 7802 11192 7807 11248
rect 0 11190 7807 11192
rect 0 11160 480 11190
rect 7741 11187 7807 11190
rect 1669 10978 1735 10981
rect 4797 10978 4863 10981
rect 1669 10976 4863 10978
rect 1669 10920 1674 10976
rect 1730 10920 4802 10976
rect 4858 10920 4863 10976
rect 1669 10918 4863 10920
rect 1669 10915 1735 10918
rect 4797 10915 4863 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 2405 10706 2471 10709
rect 13997 10706 14063 10709
rect 2405 10704 14063 10706
rect 2405 10648 2410 10704
rect 2466 10648 14002 10704
rect 14058 10648 14063 10704
rect 2405 10646 14063 10648
rect 2405 10643 2471 10646
rect 13997 10643 14063 10646
rect 0 10570 480 10600
rect 6085 10570 6151 10573
rect 0 10568 6151 10570
rect 0 10512 6090 10568
rect 6146 10512 6151 10568
rect 0 10510 6151 10512
rect 0 10480 480 10510
rect 6085 10507 6151 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5349 10026 5415 10029
rect 5993 10026 6059 10029
rect 5349 10024 6059 10026
rect 5349 9968 5354 10024
rect 5410 9968 5998 10024
rect 6054 9968 6059 10024
rect 5349 9966 6059 9968
rect 5349 9963 5415 9966
rect 5993 9963 6059 9966
rect 6177 10026 6243 10029
rect 18321 10026 18387 10029
rect 6177 10024 18387 10026
rect 6177 9968 6182 10024
rect 6238 9968 18326 10024
rect 18382 9968 18387 10024
rect 6177 9966 18387 9968
rect 6177 9963 6243 9966
rect 18321 9963 18387 9966
rect 0 9890 480 9920
rect 3509 9890 3575 9893
rect 0 9888 3575 9890
rect 0 9832 3514 9888
rect 3570 9832 3575 9888
rect 0 9830 3575 9832
rect 0 9800 480 9830
rect 3509 9827 3575 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 5441 9618 5507 9621
rect 13445 9618 13511 9621
rect 5441 9616 13511 9618
rect 5441 9560 5446 9616
rect 5502 9560 13450 9616
rect 13506 9560 13511 9616
rect 5441 9558 13511 9560
rect 5441 9555 5507 9558
rect 13445 9555 13511 9558
rect 3693 9482 3759 9485
rect 15653 9482 15719 9485
rect 22185 9482 22251 9485
rect 3693 9480 15719 9482
rect 3693 9424 3698 9480
rect 3754 9424 15658 9480
rect 15714 9424 15719 9480
rect 3693 9422 15719 9424
rect 3693 9419 3759 9422
rect 15653 9419 15719 9422
rect 17174 9480 22251 9482
rect 17174 9424 22190 9480
rect 22246 9424 22251 9480
rect 17174 9422 22251 9424
rect 12525 9346 12591 9349
rect 17174 9346 17234 9422
rect 22185 9419 22251 9422
rect 12525 9344 17234 9346
rect 12525 9288 12530 9344
rect 12586 9288 17234 9344
rect 12525 9286 17234 9288
rect 12525 9283 12591 9286
rect 10277 9280 10597 9281
rect 0 9210 480 9240
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3785 9210 3851 9213
rect 0 9208 3851 9210
rect 0 9152 3790 9208
rect 3846 9152 3851 9208
rect 0 9150 3851 9152
rect 0 9120 480 9150
rect 3785 9147 3851 9150
rect 3969 9210 4035 9213
rect 9765 9210 9831 9213
rect 3969 9208 9831 9210
rect 3969 9152 3974 9208
rect 4030 9152 9770 9208
rect 9826 9152 9831 9208
rect 3969 9150 9831 9152
rect 3969 9147 4035 9150
rect 9765 9147 9831 9150
rect 1209 9074 1275 9077
rect 12206 9074 12450 9108
rect 16205 9074 16271 9077
rect 1209 9072 16271 9074
rect 1209 9016 1214 9072
rect 1270 9048 16210 9072
rect 1270 9016 12266 9048
rect 1209 9014 12266 9016
rect 12390 9016 16210 9048
rect 16266 9016 16271 9072
rect 12390 9014 16271 9016
rect 1209 9011 1275 9014
rect 16205 9011 16271 9014
rect 9673 8938 9739 8941
rect 21633 8938 21699 8941
rect 9673 8936 21699 8938
rect 9673 8880 9678 8936
rect 9734 8880 21638 8936
rect 21694 8880 21699 8936
rect 9673 8878 21699 8880
rect 9673 8875 9739 8878
rect 21633 8875 21699 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 8477 8666 8543 8669
rect 8477 8664 14842 8666
rect 8477 8608 8482 8664
rect 8538 8608 14842 8664
rect 8477 8606 14842 8608
rect 8477 8603 8543 8606
rect 0 8530 480 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 480 8470
rect 1209 8467 1275 8470
rect 1393 8530 1459 8533
rect 14181 8530 14247 8533
rect 1393 8528 14247 8530
rect 1393 8472 1398 8528
rect 1454 8472 14186 8528
rect 14242 8472 14247 8528
rect 1393 8470 14247 8472
rect 14782 8530 14842 8606
rect 16849 8530 16915 8533
rect 14782 8528 16915 8530
rect 14782 8472 16854 8528
rect 16910 8472 16915 8528
rect 14782 8470 16915 8472
rect 1393 8467 1459 8470
rect 14181 8467 14247 8470
rect 16849 8467 16915 8470
rect 9998 8334 10794 8394
rect 3877 8258 3943 8261
rect 9998 8258 10058 8334
rect 3877 8256 10058 8258
rect 3877 8200 3882 8256
rect 3938 8200 10058 8256
rect 3877 8198 10058 8200
rect 10734 8258 10794 8334
rect 17217 8258 17283 8261
rect 10734 8256 17283 8258
rect 10734 8200 17222 8256
rect 17278 8200 17283 8256
rect 10734 8198 17283 8200
rect 3877 8195 3943 8198
rect 17217 8195 17283 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 3785 8122 3851 8125
rect 9305 8122 9371 8125
rect 3785 8120 9371 8122
rect 3785 8064 3790 8120
rect 3846 8064 9310 8120
rect 9366 8064 9371 8120
rect 3785 8062 9371 8064
rect 3785 8059 3851 8062
rect 9305 8059 9371 8062
rect 11329 8122 11395 8125
rect 15653 8122 15719 8125
rect 11329 8120 15719 8122
rect 11329 8064 11334 8120
rect 11390 8064 15658 8120
rect 15714 8064 15719 8120
rect 11329 8062 15719 8064
rect 11329 8059 11395 8062
rect 15653 8059 15719 8062
rect 5073 7986 5139 7989
rect 20529 7986 20595 7989
rect 5073 7984 20595 7986
rect 5073 7928 5078 7984
rect 5134 7928 20534 7984
rect 20590 7928 20595 7984
rect 5073 7926 20595 7928
rect 5073 7923 5139 7926
rect 20529 7923 20595 7926
rect 0 7850 480 7880
rect 3693 7850 3759 7853
rect 0 7848 3759 7850
rect 0 7792 3698 7848
rect 3754 7792 3759 7848
rect 0 7790 3759 7792
rect 0 7760 480 7790
rect 3693 7787 3759 7790
rect 7557 7850 7623 7853
rect 21081 7850 21147 7853
rect 7557 7848 21147 7850
rect 7557 7792 7562 7848
rect 7618 7792 21086 7848
rect 21142 7792 21147 7848
rect 7557 7790 21147 7792
rect 7557 7787 7623 7790
rect 21081 7787 21147 7790
rect 7925 7714 7991 7717
rect 13721 7714 13787 7717
rect 7925 7712 13787 7714
rect 7925 7656 7930 7712
rect 7986 7656 13726 7712
rect 13782 7656 13787 7712
rect 7925 7654 13787 7656
rect 7925 7651 7991 7654
rect 13721 7651 13787 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 4613 7442 4679 7445
rect 6913 7442 6979 7445
rect 4613 7440 6979 7442
rect 4613 7384 4618 7440
rect 4674 7384 6918 7440
rect 6974 7384 6979 7440
rect 4613 7382 6979 7384
rect 4613 7379 4679 7382
rect 6913 7379 6979 7382
rect 8569 7442 8635 7445
rect 11053 7442 11119 7445
rect 8569 7440 11119 7442
rect 8569 7384 8574 7440
rect 8630 7384 11058 7440
rect 11114 7384 11119 7440
rect 8569 7382 11119 7384
rect 8569 7379 8635 7382
rect 11053 7379 11119 7382
rect 12985 7442 13051 7445
rect 17309 7442 17375 7445
rect 12985 7440 17375 7442
rect 12985 7384 12990 7440
rect 13046 7384 17314 7440
rect 17370 7384 17375 7440
rect 12985 7382 17375 7384
rect 12985 7379 13051 7382
rect 17309 7379 17375 7382
rect 5533 7306 5599 7309
rect 12157 7306 12223 7309
rect 5533 7304 12223 7306
rect 5533 7248 5538 7304
rect 5594 7248 12162 7304
rect 12218 7248 12223 7304
rect 5533 7246 12223 7248
rect 5533 7243 5599 7246
rect 12157 7243 12223 7246
rect 13629 7306 13695 7309
rect 23841 7306 23907 7309
rect 13629 7304 23907 7306
rect 13629 7248 13634 7304
rect 13690 7248 23846 7304
rect 23902 7248 23907 7304
rect 13629 7246 23907 7248
rect 13629 7243 13695 7246
rect 23841 7243 23907 7246
rect 0 7170 480 7200
rect 3877 7170 3943 7173
rect 0 7168 3943 7170
rect 0 7112 3882 7168
rect 3938 7112 3943 7168
rect 0 7110 3943 7112
rect 0 7080 480 7110
rect 3877 7107 3943 7110
rect 15285 7170 15351 7173
rect 19149 7170 19215 7173
rect 15285 7168 19215 7170
rect 15285 7112 15290 7168
rect 15346 7112 19154 7168
rect 19210 7112 19215 7168
rect 15285 7110 19215 7112
rect 15285 7107 15351 7110
rect 19149 7107 19215 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 10961 7034 11027 7037
rect 19425 7034 19491 7037
rect 10961 7032 19491 7034
rect 10961 6976 10966 7032
rect 11022 6976 19430 7032
rect 19486 6976 19491 7032
rect 10961 6974 19491 6976
rect 10961 6971 11027 6974
rect 19425 6971 19491 6974
rect 2497 6898 2563 6901
rect 5533 6898 5599 6901
rect 2497 6896 5599 6898
rect 2497 6840 2502 6896
rect 2558 6840 5538 6896
rect 5594 6840 5599 6896
rect 2497 6838 5599 6840
rect 2497 6835 2563 6838
rect 5533 6835 5599 6838
rect 6729 6898 6795 6901
rect 11053 6898 11119 6901
rect 6729 6896 11119 6898
rect 6729 6840 6734 6896
rect 6790 6840 11058 6896
rect 11114 6840 11119 6896
rect 6729 6838 11119 6840
rect 6729 6835 6795 6838
rect 11053 6835 11119 6838
rect 13077 6898 13143 6901
rect 15929 6898 15995 6901
rect 13077 6896 15995 6898
rect 13077 6840 13082 6896
rect 13138 6840 15934 6896
rect 15990 6840 15995 6896
rect 13077 6838 15995 6840
rect 13077 6835 13143 6838
rect 15929 6835 15995 6838
rect 3233 6762 3299 6765
rect 9305 6762 9371 6765
rect 3233 6760 9371 6762
rect 3233 6704 3238 6760
rect 3294 6704 9310 6760
rect 9366 6704 9371 6760
rect 3233 6702 9371 6704
rect 3233 6699 3299 6702
rect 9305 6699 9371 6702
rect 13721 6762 13787 6765
rect 19977 6762 20043 6765
rect 13721 6760 20043 6762
rect 13721 6704 13726 6760
rect 13782 6704 19982 6760
rect 20038 6704 20043 6760
rect 13721 6702 20043 6704
rect 13721 6699 13787 6702
rect 19977 6699 20043 6702
rect 8385 6626 8451 6629
rect 9765 6626 9831 6629
rect 8385 6624 9831 6626
rect 8385 6568 8390 6624
rect 8446 6568 9770 6624
rect 9826 6568 9831 6624
rect 8385 6566 9831 6568
rect 8385 6563 8451 6566
rect 9765 6563 9831 6566
rect 5610 6560 5930 6561
rect 0 6490 480 6520
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 21265 6490 21331 6493
rect 0 6430 1824 6490
rect 0 6400 480 6430
rect 1764 6218 1824 6430
rect 15702 6488 21331 6490
rect 15702 6432 21270 6488
rect 21326 6432 21331 6488
rect 15702 6430 21331 6432
rect 11605 6354 11671 6357
rect 15702 6354 15762 6430
rect 21265 6427 21331 6430
rect 11605 6352 15762 6354
rect 11605 6296 11610 6352
rect 11666 6296 15762 6352
rect 11605 6294 15762 6296
rect 15837 6354 15903 6357
rect 18505 6354 18571 6357
rect 15837 6352 18571 6354
rect 15837 6296 15842 6352
rect 15898 6296 18510 6352
rect 18566 6296 18571 6352
rect 15837 6294 18571 6296
rect 11605 6291 11671 6294
rect 15837 6291 15903 6294
rect 18505 6291 18571 6294
rect 12157 6218 12223 6221
rect 1764 6216 12223 6218
rect 1764 6160 12162 6216
rect 12218 6160 12223 6216
rect 1764 6158 12223 6160
rect 12157 6155 12223 6158
rect 13813 6218 13879 6221
rect 16941 6218 17007 6221
rect 13813 6216 17007 6218
rect 13813 6160 13818 6216
rect 13874 6160 16946 6216
rect 17002 6160 17007 6216
rect 13813 6158 17007 6160
rect 13813 6155 13879 6158
rect 16941 6155 17007 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 13629 5946 13695 5949
rect 17309 5946 17375 5949
rect 13629 5944 17375 5946
rect 13629 5888 13634 5944
rect 13690 5888 17314 5944
rect 17370 5888 17375 5944
rect 13629 5886 17375 5888
rect 13629 5883 13695 5886
rect 17309 5883 17375 5886
rect 0 5810 480 5840
rect 10041 5810 10107 5813
rect 0 5808 10107 5810
rect 0 5752 10046 5808
rect 10102 5752 10107 5808
rect 0 5750 10107 5752
rect 0 5720 480 5750
rect 10041 5747 10107 5750
rect 14365 5810 14431 5813
rect 18137 5810 18203 5813
rect 14365 5808 18203 5810
rect 14365 5752 14370 5808
rect 14426 5752 18142 5808
rect 18198 5752 18203 5808
rect 14365 5750 18203 5752
rect 14365 5747 14431 5750
rect 18137 5747 18203 5750
rect 18321 5810 18387 5813
rect 24669 5810 24735 5813
rect 18321 5808 24735 5810
rect 18321 5752 18326 5808
rect 18382 5752 24674 5808
rect 24730 5752 24735 5808
rect 18321 5750 24735 5752
rect 18321 5747 18387 5750
rect 24669 5747 24735 5750
rect 7005 5674 7071 5677
rect 11329 5674 11395 5677
rect 7005 5672 11395 5674
rect 7005 5616 7010 5672
rect 7066 5616 11334 5672
rect 11390 5616 11395 5672
rect 7005 5614 11395 5616
rect 7005 5611 7071 5614
rect 11329 5611 11395 5614
rect 11513 5674 11579 5677
rect 15009 5674 15075 5677
rect 11513 5672 15075 5674
rect 11513 5616 11518 5672
rect 11574 5616 15014 5672
rect 15070 5616 15075 5672
rect 11513 5614 15075 5616
rect 11513 5611 11579 5614
rect 15009 5611 15075 5614
rect 19241 5674 19307 5677
rect 21081 5674 21147 5677
rect 19241 5672 21147 5674
rect 19241 5616 19246 5672
rect 19302 5616 21086 5672
rect 21142 5616 21147 5672
rect 19241 5614 21147 5616
rect 19241 5611 19307 5614
rect 21081 5611 21147 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 6821 5402 6887 5405
rect 8477 5402 8543 5405
rect 19425 5402 19491 5405
rect 6821 5400 8543 5402
rect 6821 5344 6826 5400
rect 6882 5344 8482 5400
rect 8538 5344 8543 5400
rect 6821 5342 8543 5344
rect 6821 5339 6887 5342
rect 8477 5339 8543 5342
rect 16070 5400 19491 5402
rect 16070 5344 19430 5400
rect 19486 5344 19491 5400
rect 16070 5342 19491 5344
rect 10133 5266 10199 5269
rect 16070 5266 16130 5342
rect 19425 5339 19491 5342
rect 10133 5264 16130 5266
rect 10133 5208 10138 5264
rect 10194 5208 16130 5264
rect 10133 5206 16130 5208
rect 16205 5266 16271 5269
rect 20897 5266 20963 5269
rect 16205 5264 20963 5266
rect 16205 5208 16210 5264
rect 16266 5208 20902 5264
rect 20958 5208 20963 5264
rect 16205 5206 20963 5208
rect 10133 5203 10199 5206
rect 16205 5203 16271 5206
rect 20897 5203 20963 5206
rect 0 5130 480 5160
rect 8385 5130 8451 5133
rect 0 5128 8451 5130
rect 0 5072 8390 5128
rect 8446 5072 8451 5128
rect 0 5070 8451 5072
rect 0 5040 480 5070
rect 8385 5067 8451 5070
rect 8569 5130 8635 5133
rect 11237 5130 11303 5133
rect 8569 5128 11303 5130
rect 8569 5072 8574 5128
rect 8630 5072 11242 5128
rect 11298 5072 11303 5128
rect 8569 5070 11303 5072
rect 8569 5067 8635 5070
rect 11237 5067 11303 5070
rect 18045 5130 18111 5133
rect 22093 5130 22159 5133
rect 18045 5128 22159 5130
rect 18045 5072 18050 5128
rect 18106 5072 22098 5128
rect 22154 5072 22159 5128
rect 18045 5070 22159 5072
rect 18045 5067 18111 5070
rect 22093 5067 22159 5070
rect 4981 4994 5047 4997
rect 6637 4994 6703 4997
rect 10041 4994 10107 4997
rect 4981 4992 10107 4994
rect 4981 4936 4986 4992
rect 5042 4936 6642 4992
rect 6698 4936 10046 4992
rect 10102 4936 10107 4992
rect 4981 4934 10107 4936
rect 4981 4931 5047 4934
rect 6637 4931 6703 4934
rect 10041 4931 10107 4934
rect 11329 4994 11395 4997
rect 17769 4994 17835 4997
rect 11329 4992 17835 4994
rect 11329 4936 11334 4992
rect 11390 4936 17774 4992
rect 17830 4936 17835 4992
rect 11329 4934 17835 4936
rect 11329 4931 11395 4934
rect 17769 4931 17835 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 5349 4858 5415 4861
rect 8753 4858 8819 4861
rect 5349 4856 8819 4858
rect 5349 4800 5354 4856
rect 5410 4800 8758 4856
rect 8814 4800 8819 4856
rect 5349 4798 8819 4800
rect 5349 4795 5415 4798
rect 8753 4795 8819 4798
rect 14825 4858 14891 4861
rect 17953 4858 18019 4861
rect 14825 4856 18019 4858
rect 14825 4800 14830 4856
rect 14886 4800 17958 4856
rect 18014 4800 18019 4856
rect 14825 4798 18019 4800
rect 14825 4795 14891 4798
rect 17953 4795 18019 4798
rect 2681 4722 2747 4725
rect 5625 4722 5691 4725
rect 2681 4720 5691 4722
rect 2681 4664 2686 4720
rect 2742 4664 5630 4720
rect 5686 4664 5691 4720
rect 2681 4662 5691 4664
rect 2681 4659 2747 4662
rect 5625 4659 5691 4662
rect 10041 4722 10107 4725
rect 16849 4722 16915 4725
rect 10041 4720 16915 4722
rect 10041 4664 10046 4720
rect 10102 4664 16854 4720
rect 16910 4664 16915 4720
rect 10041 4662 16915 4664
rect 10041 4659 10107 4662
rect 16849 4659 16915 4662
rect 24669 4722 24735 4725
rect 27520 4722 28000 4752
rect 24669 4720 28000 4722
rect 24669 4664 24674 4720
rect 24730 4664 28000 4720
rect 24669 4662 28000 4664
rect 24669 4659 24735 4662
rect 27520 4632 28000 4662
rect 2405 4586 2471 4589
rect 13077 4586 13143 4589
rect 22185 4586 22251 4589
rect 2405 4584 12266 4586
rect 2405 4528 2410 4584
rect 2466 4528 12266 4584
rect 2405 4526 12266 4528
rect 2405 4523 2471 4526
rect 0 4450 480 4480
rect 4705 4450 4771 4453
rect 0 4448 4771 4450
rect 0 4392 4710 4448
rect 4766 4392 4771 4448
rect 0 4390 4771 4392
rect 0 4360 480 4390
rect 4705 4387 4771 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 1393 4314 1459 4317
rect 4981 4314 5047 4317
rect 1393 4312 5047 4314
rect 1393 4256 1398 4312
rect 1454 4256 4986 4312
rect 5042 4256 5047 4312
rect 1393 4254 5047 4256
rect 1393 4251 1459 4254
rect 4981 4251 5047 4254
rect 1761 4178 1827 4181
rect 4889 4178 4955 4181
rect 1761 4176 4955 4178
rect 1761 4120 1766 4176
rect 1822 4120 4894 4176
rect 4950 4120 4955 4176
rect 1761 4118 4955 4120
rect 1761 4115 1827 4118
rect 4889 4115 4955 4118
rect 8017 4178 8083 4181
rect 11329 4178 11395 4181
rect 8017 4176 11395 4178
rect 8017 4120 8022 4176
rect 8078 4120 11334 4176
rect 11390 4120 11395 4176
rect 8017 4118 11395 4120
rect 12206 4178 12266 4526
rect 13077 4584 22251 4586
rect 13077 4528 13082 4584
rect 13138 4528 22190 4584
rect 22246 4528 22251 4584
rect 13077 4526 22251 4528
rect 13077 4523 13143 4526
rect 22185 4523 22251 4526
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 15745 4178 15811 4181
rect 12206 4176 15811 4178
rect 12206 4120 15750 4176
rect 15806 4120 15811 4176
rect 12206 4118 15811 4120
rect 8017 4115 8083 4118
rect 11329 4115 11395 4118
rect 15745 4115 15811 4118
rect 20161 4178 20227 4181
rect 22553 4178 22619 4181
rect 20161 4176 22619 4178
rect 20161 4120 20166 4176
rect 20222 4120 22558 4176
rect 22614 4120 22619 4176
rect 20161 4118 22619 4120
rect 20161 4115 20227 4118
rect 22553 4115 22619 4118
rect 4337 4042 4403 4045
rect 9673 4042 9739 4045
rect 4337 4040 9739 4042
rect 4337 3984 4342 4040
rect 4398 3984 9678 4040
rect 9734 3984 9739 4040
rect 4337 3982 9739 3984
rect 4337 3979 4403 3982
rect 9673 3979 9739 3982
rect 10777 4042 10843 4045
rect 11145 4042 11211 4045
rect 10777 4040 11211 4042
rect 10777 3984 10782 4040
rect 10838 3984 11150 4040
rect 11206 3984 11211 4040
rect 10777 3982 11211 3984
rect 10777 3979 10843 3982
rect 11145 3979 11211 3982
rect 15837 4042 15903 4045
rect 17401 4042 17467 4045
rect 15837 4040 17467 4042
rect 15837 3984 15842 4040
rect 15898 3984 17406 4040
rect 17462 3984 17467 4040
rect 15837 3982 17467 3984
rect 15837 3979 15903 3982
rect 17401 3979 17467 3982
rect 19793 4042 19859 4045
rect 22093 4042 22159 4045
rect 19793 4040 22159 4042
rect 19793 3984 19798 4040
rect 19854 3984 22098 4040
rect 22154 3984 22159 4040
rect 19793 3982 22159 3984
rect 19793 3979 19859 3982
rect 22093 3979 22159 3982
rect 24117 4042 24183 4045
rect 25957 4042 26023 4045
rect 24117 4040 26023 4042
rect 24117 3984 24122 4040
rect 24178 3984 25962 4040
rect 26018 3984 26023 4040
rect 24117 3982 26023 3984
rect 24117 3979 24183 3982
rect 25957 3979 26023 3982
rect 4245 3906 4311 3909
rect 7005 3906 7071 3909
rect 4245 3904 7071 3906
rect 4245 3848 4250 3904
rect 4306 3848 7010 3904
rect 7066 3848 7071 3904
rect 4245 3846 7071 3848
rect 4245 3843 4311 3846
rect 7005 3843 7071 3846
rect 10777 3906 10843 3909
rect 12893 3906 12959 3909
rect 10777 3904 12959 3906
rect 10777 3848 10782 3904
rect 10838 3848 12898 3904
rect 12954 3848 12959 3904
rect 10777 3846 12959 3848
rect 10777 3843 10843 3846
rect 12893 3843 12959 3846
rect 14457 3906 14523 3909
rect 17677 3906 17743 3909
rect 19241 3906 19307 3909
rect 14457 3904 19307 3906
rect 14457 3848 14462 3904
rect 14518 3848 17682 3904
rect 17738 3848 19246 3904
rect 19302 3848 19307 3904
rect 14457 3846 19307 3848
rect 14457 3843 14523 3846
rect 17677 3843 17743 3846
rect 19241 3843 19307 3846
rect 23841 3906 23907 3909
rect 25313 3906 25379 3909
rect 23841 3904 25379 3906
rect 23841 3848 23846 3904
rect 23902 3848 25318 3904
rect 25374 3848 25379 3904
rect 23841 3846 25379 3848
rect 23841 3843 23907 3846
rect 25313 3843 25379 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2313 3770 2379 3773
rect 0 3768 2379 3770
rect 0 3712 2318 3768
rect 2374 3712 2379 3768
rect 0 3710 2379 3712
rect 0 3680 480 3710
rect 2313 3707 2379 3710
rect 3693 3770 3759 3773
rect 8293 3770 8359 3773
rect 3693 3768 8359 3770
rect 3693 3712 3698 3768
rect 3754 3712 8298 3768
rect 8354 3712 8359 3768
rect 3693 3710 8359 3712
rect 3693 3707 3759 3710
rect 8293 3707 8359 3710
rect 11145 3770 11211 3773
rect 19333 3770 19399 3773
rect 11145 3768 19399 3770
rect 11145 3712 11150 3768
rect 11206 3712 19338 3768
rect 19394 3712 19399 3768
rect 11145 3710 19399 3712
rect 11145 3707 11211 3710
rect 19333 3707 19399 3710
rect 22369 3770 22435 3773
rect 24209 3770 24275 3773
rect 22369 3768 24275 3770
rect 22369 3712 22374 3768
rect 22430 3712 24214 3768
rect 24270 3712 24275 3768
rect 22369 3710 24275 3712
rect 22369 3707 22435 3710
rect 24209 3707 24275 3710
rect 3325 3634 3391 3637
rect 4245 3634 4311 3637
rect 3325 3632 4311 3634
rect 3325 3576 3330 3632
rect 3386 3576 4250 3632
rect 4306 3576 4311 3632
rect 3325 3574 4311 3576
rect 3325 3571 3391 3574
rect 4245 3571 4311 3574
rect 8109 3634 8175 3637
rect 12157 3634 12223 3637
rect 8109 3632 12223 3634
rect 8109 3576 8114 3632
rect 8170 3576 12162 3632
rect 12218 3576 12223 3632
rect 8109 3574 12223 3576
rect 8109 3571 8175 3574
rect 12157 3571 12223 3574
rect 15653 3634 15719 3637
rect 20897 3634 20963 3637
rect 15653 3632 20963 3634
rect 15653 3576 15658 3632
rect 15714 3576 20902 3632
rect 20958 3576 20963 3632
rect 15653 3574 20963 3576
rect 15653 3571 15719 3574
rect 20897 3571 20963 3574
rect 22921 3634 22987 3637
rect 24669 3634 24735 3637
rect 22921 3632 24735 3634
rect 22921 3576 22926 3632
rect 22982 3576 24674 3632
rect 24730 3576 24735 3632
rect 22921 3574 24735 3576
rect 22921 3571 22987 3574
rect 24669 3571 24735 3574
rect 8937 3498 9003 3501
rect 14457 3498 14523 3501
rect 21081 3498 21147 3501
rect 8937 3496 14523 3498
rect 8937 3440 8942 3496
rect 8998 3440 14462 3496
rect 14518 3440 14523 3496
rect 8937 3438 14523 3440
rect 8937 3435 9003 3438
rect 14457 3435 14523 3438
rect 14782 3496 21147 3498
rect 14782 3440 21086 3496
rect 21142 3440 21147 3496
rect 14782 3438 21147 3440
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 6085 3226 6151 3229
rect 14457 3226 14523 3229
rect 6085 3224 14523 3226
rect 6085 3168 6090 3224
rect 6146 3168 14462 3224
rect 14518 3168 14523 3224
rect 6085 3166 14523 3168
rect 6085 3163 6151 3166
rect 14457 3163 14523 3166
rect 0 3090 480 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 480 3030
rect 1577 3027 1643 3030
rect 8753 3090 8819 3093
rect 14782 3090 14842 3438
rect 21081 3435 21147 3438
rect 21265 3498 21331 3501
rect 22461 3498 22527 3501
rect 21265 3496 22527 3498
rect 21265 3440 21270 3496
rect 21326 3440 22466 3496
rect 22522 3440 22527 3496
rect 21265 3438 22527 3440
rect 21265 3435 21331 3438
rect 22461 3435 22527 3438
rect 15469 3362 15535 3365
rect 20713 3362 20779 3365
rect 15469 3360 20779 3362
rect 15469 3304 15474 3360
rect 15530 3304 20718 3360
rect 20774 3304 20779 3360
rect 15469 3302 20779 3304
rect 15469 3299 15535 3302
rect 20713 3299 20779 3302
rect 21173 3362 21239 3365
rect 23105 3362 23171 3365
rect 21173 3360 23171 3362
rect 21173 3304 21178 3360
rect 21234 3304 23110 3360
rect 23166 3304 23171 3360
rect 21173 3302 23171 3304
rect 21173 3299 21239 3302
rect 23105 3299 23171 3302
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 15745 3226 15811 3229
rect 21265 3226 21331 3229
rect 15745 3224 21331 3226
rect 15745 3168 15750 3224
rect 15806 3168 21270 3224
rect 21326 3168 21331 3224
rect 15745 3166 21331 3168
rect 15745 3163 15811 3166
rect 21265 3163 21331 3166
rect 21909 3226 21975 3229
rect 23657 3226 23723 3229
rect 21909 3224 23723 3226
rect 21909 3168 21914 3224
rect 21970 3168 23662 3224
rect 23718 3168 23723 3224
rect 21909 3166 23723 3168
rect 21909 3163 21975 3166
rect 23657 3163 23723 3166
rect 8753 3088 14842 3090
rect 8753 3032 8758 3088
rect 8814 3032 14842 3088
rect 8753 3030 14842 3032
rect 15285 3090 15351 3093
rect 23289 3090 23355 3093
rect 27613 3090 27679 3093
rect 15285 3088 23355 3090
rect 15285 3032 15290 3088
rect 15346 3032 23294 3088
rect 23350 3032 23355 3088
rect 15285 3030 23355 3032
rect 8753 3027 8819 3030
rect 15285 3027 15351 3030
rect 23289 3027 23355 3030
rect 24350 3088 27679 3090
rect 24350 3032 27618 3088
rect 27674 3032 27679 3088
rect 24350 3030 27679 3032
rect 4061 2954 4127 2957
rect 10409 2954 10475 2957
rect 4061 2952 10475 2954
rect 4061 2896 4066 2952
rect 4122 2896 10414 2952
rect 10470 2896 10475 2952
rect 4061 2894 10475 2896
rect 4061 2891 4127 2894
rect 10409 2891 10475 2894
rect 14273 2954 14339 2957
rect 16757 2954 16823 2957
rect 14273 2952 16823 2954
rect 14273 2896 14278 2952
rect 14334 2896 16762 2952
rect 16818 2896 16823 2952
rect 14273 2894 16823 2896
rect 14273 2891 14339 2894
rect 16757 2891 16823 2894
rect 20069 2954 20135 2957
rect 24350 2954 24410 3030
rect 27613 3027 27679 3030
rect 20069 2952 24410 2954
rect 20069 2896 20074 2952
rect 20130 2896 24410 2952
rect 20069 2894 24410 2896
rect 24577 2954 24643 2957
rect 26509 2954 26575 2957
rect 24577 2952 26575 2954
rect 24577 2896 24582 2952
rect 24638 2896 26514 2952
rect 26570 2896 26575 2952
rect 24577 2894 26575 2896
rect 20069 2891 20135 2894
rect 24577 2891 24643 2894
rect 26509 2891 26575 2894
rect 14457 2818 14523 2821
rect 15929 2818 15995 2821
rect 16205 2818 16271 2821
rect 14457 2816 16271 2818
rect 14457 2760 14462 2816
rect 14518 2760 15934 2816
rect 15990 2760 16210 2816
rect 16266 2760 16271 2816
rect 14457 2758 16271 2760
rect 14457 2755 14523 2758
rect 15929 2755 15995 2758
rect 16205 2755 16271 2758
rect 16389 2818 16455 2821
rect 18505 2818 18571 2821
rect 16389 2816 18571 2818
rect 16389 2760 16394 2816
rect 16450 2760 18510 2816
rect 18566 2760 18571 2816
rect 16389 2758 18571 2760
rect 16389 2755 16455 2758
rect 18505 2755 18571 2758
rect 24761 2818 24827 2821
rect 27061 2818 27127 2821
rect 24761 2816 27127 2818
rect 24761 2760 24766 2816
rect 24822 2760 27066 2816
rect 27122 2760 27127 2816
rect 24761 2758 27127 2760
rect 24761 2755 24827 2758
rect 27061 2755 27127 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 10777 2682 10843 2685
rect 18045 2682 18111 2685
rect 10777 2680 18111 2682
rect 10777 2624 10782 2680
rect 10838 2624 18050 2680
rect 18106 2624 18111 2680
rect 10777 2622 18111 2624
rect 10777 2619 10843 2622
rect 18045 2619 18111 2622
rect 6361 2546 6427 2549
rect 14273 2546 14339 2549
rect 6361 2544 14339 2546
rect 6361 2488 6366 2544
rect 6422 2488 14278 2544
rect 14334 2488 14339 2544
rect 6361 2486 14339 2488
rect 6361 2483 6427 2486
rect 14273 2483 14339 2486
rect 18413 2546 18479 2549
rect 21173 2546 21239 2549
rect 18413 2544 21239 2546
rect 18413 2488 18418 2544
rect 18474 2488 21178 2544
rect 21234 2488 21239 2544
rect 18413 2486 21239 2488
rect 18413 2483 18479 2486
rect 21173 2483 21239 2486
rect 0 2410 480 2440
rect 17677 2410 17743 2413
rect 0 2408 17743 2410
rect 0 2352 17682 2408
rect 17738 2352 17743 2408
rect 0 2350 17743 2352
rect 0 2320 480 2350
rect 17677 2347 17743 2350
rect 18229 2410 18295 2413
rect 22921 2410 22987 2413
rect 18229 2408 22987 2410
rect 18229 2352 18234 2408
rect 18290 2352 22926 2408
rect 22982 2352 22987 2408
rect 18229 2350 22987 2352
rect 18229 2347 18295 2350
rect 22921 2347 22987 2350
rect 11329 2274 11395 2277
rect 14365 2274 14431 2277
rect 11329 2272 14431 2274
rect 11329 2216 11334 2272
rect 11390 2216 14370 2272
rect 14426 2216 14431 2272
rect 11329 2214 14431 2216
rect 11329 2211 11395 2214
rect 14365 2211 14431 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 1945 2002 2011 2005
rect 10777 2002 10843 2005
rect 1945 2000 10843 2002
rect 1945 1944 1950 2000
rect 2006 1944 10782 2000
rect 10838 1944 10843 2000
rect 1945 1942 10843 1944
rect 1945 1939 2011 1942
rect 10777 1939 10843 1942
rect 14641 2002 14707 2005
rect 19885 2002 19951 2005
rect 14641 2000 19951 2002
rect 14641 1944 14646 2000
rect 14702 1944 19890 2000
rect 19946 1944 19951 2000
rect 14641 1942 19951 1944
rect 14641 1939 14707 1942
rect 19885 1939 19951 1942
rect 3141 1866 3207 1869
rect 10409 1866 10475 1869
rect 3141 1864 10475 1866
rect 3141 1808 3146 1864
rect 3202 1808 10414 1864
rect 10470 1808 10475 1864
rect 3141 1806 10475 1808
rect 3141 1803 3207 1806
rect 10409 1803 10475 1806
rect 11145 1866 11211 1869
rect 19425 1866 19491 1869
rect 11145 1864 19491 1866
rect 11145 1808 11150 1864
rect 11206 1808 19430 1864
rect 19486 1808 19491 1864
rect 11145 1806 19491 1808
rect 11145 1803 11211 1806
rect 19425 1803 19491 1806
rect 0 1730 480 1760
rect 2221 1730 2287 1733
rect 0 1728 2287 1730
rect 0 1672 2226 1728
rect 2282 1672 2287 1728
rect 0 1670 2287 1672
rect 0 1640 480 1670
rect 2221 1667 2287 1670
rect 8385 1730 8451 1733
rect 18321 1730 18387 1733
rect 8385 1728 18387 1730
rect 8385 1672 8390 1728
rect 8446 1672 18326 1728
rect 18382 1672 18387 1728
rect 8385 1670 18387 1672
rect 8385 1667 8451 1670
rect 18321 1667 18387 1670
rect 9857 1594 9923 1597
rect 22369 1594 22435 1597
rect 9857 1592 22435 1594
rect 9857 1536 9862 1592
rect 9918 1536 22374 1592
rect 22430 1536 22435 1592
rect 9857 1534 22435 1536
rect 9857 1531 9923 1534
rect 22369 1531 22435 1534
rect 10041 1458 10107 1461
rect 16205 1458 16271 1461
rect 10041 1456 16271 1458
rect 10041 1400 10046 1456
rect 10102 1400 16210 1456
rect 16266 1400 16271 1456
rect 10041 1398 16271 1400
rect 10041 1395 10107 1398
rect 16205 1395 16271 1398
rect 0 1050 480 1080
rect 4061 1050 4127 1053
rect 0 1048 4127 1050
rect 0 992 4066 1048
rect 4122 992 4127 1048
rect 0 990 4127 992
rect 0 960 480 990
rect 4061 987 4127 990
rect 0 370 480 400
rect 0 310 4906 370
rect 0 280 480 310
rect 4846 98 4906 310
rect 15837 98 15903 101
rect 4846 96 15903 98
rect 4846 40 15842 96
rect 15898 40 15903 96
rect 4846 38 15903 40
rect 15837 35 15903 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _29_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_11
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_66 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_70
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_0_82
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_86
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__87__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _87_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_99
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_148
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_152
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_39.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_162
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_39.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _83_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__82__A
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__83__A
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 406 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_3.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_233
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_39.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_221 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_245 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_249 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_261
timestamp 1586364061
transform 1 0 25116 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_273
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1472 0 -1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_37
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_54
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_58
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_85
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_133
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _86_
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_37.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _82_
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 406 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21344 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_222
timestamp 1586364061
transform 1 0 21528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_234
timestamp 1586364061
transform 1 0 22632 0 -1 3808
box -38 -48 590 592
use scs8hd_buf_1  mux_bottom_track_37.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_240
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_244
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_256
timestamp 1586364061
transform 1 0 24656 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_268
timestamp 1586364061
transform 1 0 25760 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_conb_1  _46_
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_33
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_37
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_50
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_54
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_79
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 1786 592
use scs8hd_buf_1  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_170
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _84_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__81__A
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__84__A
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_188
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_192
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _78_
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_200
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_228
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _36_
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_37
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 314 592
use scs8hd_conb_1  _38_
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_112
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_37.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__86__A
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _81_
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_192
timestamp 1586364061
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_204
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_253
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_265
timestamp 1586364061
transform 1 0 25484 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_273
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _37_
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_106
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _40_
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_129
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 590 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_209
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_213
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_235
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_76
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_137
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_152
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__85__A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _85_
timestamp 1586364061
transform 1 0 15364 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_188
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_192
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19136 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_212
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 20976 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_220
timestamp 1586364061
transform 1 0 21344 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_244
timestamp 1586364061
transform 1 0 23552 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_256
timestamp 1586364061
transform 1 0 24656 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_250
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_268
timestamp 1586364061
transform 1 0 25760 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_262
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_274
timestamp 1586364061
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_9
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_13
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_28
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_169
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_173
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 22172 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_233
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_252
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_264
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_20
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_68
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_72
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _39_
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_35.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12512 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_133
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _41_
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_27.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_237
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 590 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_35
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _44_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_112
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_35.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _42_
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_180
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_195
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_29.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_207
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_220
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_35.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_262
timestamp 1586364061
transform 1 0 25208 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_11_58
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use scs8hd_conb_1  _45_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_65
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_96
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_165
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_31.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_242
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_14
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_31.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_114
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22172 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_244
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_256
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_268
timestamp 1586364061
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_31.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_77
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _43_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 314 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_126
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_191
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_203
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 590 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _47_
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_79
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_25
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_127
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_139
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_151
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_163
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_14
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_14
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_26
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_51
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_107
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use scs8hd_conb_1  _34_
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_37
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_13
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_21
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_23_29
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_48
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 1142 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_24_48
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_52
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_78
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_90
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 406 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 5244 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_65
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_18
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 406 592
use scs8hd_buf_1  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 1142 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_6  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 8096 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_96
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_108
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_120
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_19
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_43
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_55
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_31
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_55
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_35
timestamp 1586364061
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_47
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3698 0 3754 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 4250 0 4306 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 27618 0 27674 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_head
port 9 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 960 480 1080 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 1640 480 1760 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 2320 480 2440 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 24080 480 24200 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 25440 480 25560 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 26120 480 26240 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 26800 480 26920 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 15240 480 15360 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 23110 0 23166 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 23662 0 23718 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal3 s 0 27480 480 27600 6 left_top_grid_pin_1_
port 91 nsew default input
rlabel metal3 s 27520 4632 28000 4752 6 prog_clk
port 92 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 93 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27600
<< end >>
