* NGSPICE file created from sb_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt sb_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] data_in enable left_bottom_grid_pin_12_
+ left_top_grid_pin_11_ left_top_grid_pin_13_ left_top_grid_pin_15_ left_top_grid_pin_1_
+ left_top_grid_pin_3_ left_top_grid_pin_5_ left_top_grid_pin_7_ left_top_grid_pin_9_
+ right_bottom_grid_pin_12_ right_top_grid_pin_11_ right_top_grid_pin_13_ right_top_grid_pin_15_
+ right_top_grid_pin_1_ right_top_grid_pin_3_ right_top_grid_pin_5_ right_top_grid_pin_7_
+ right_top_grid_pin_9_ vpwr vgnd
XFILLER_22_199 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_74 vgnd vpwr scs8hd_decap_6
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_166 vpwr vgnd scs8hd_fill_2
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
XFILLER_3_12 vpwr vgnd scs8hd_fill_2
XFILLER_3_78 vpwr vgnd scs8hd_fill_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_107 vgnd vpwr scs8hd_decap_3
XFILLER_6_129 vgnd vpwr scs8hd_decap_4
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XFILLER_12_65 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XANTENNA__108__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__124__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_23_272 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
X_131_ _131_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_97 vgnd vpwr scs8hd_fill_1
XFILLER_2_176 vpwr vgnd scs8hd_fill_2
XFILLER_0_68 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_11 vpwr vgnd scs8hd_fill_2
XFILLER_9_88 vgnd vpwr scs8hd_decap_4
XFILLER_14_250 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
XFILLER_12_209 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _188_/Y mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_11_275 vpwr vgnd scs8hd_fill_2
X_114_ _113_/Y address[4] _089_/C _114_/X vgnd vpwr scs8hd_or3_4
XANTENNA__105__C _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_7 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_106 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_3
XANTENNA__222__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__116__B _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _150_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_172 vpwr vgnd scs8hd_fill_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_109 vgnd vpwr scs8hd_fill_1
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__127__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_186 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_123 vpwr vgnd scs8hd_fill_2
XFILLER_26_20 vgnd vpwr scs8hd_decap_8
XFILLER_13_156 vgnd vpwr scs8hd_fill_1
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_119 vgnd vpwr scs8hd_decap_4
XFILLER_10_115 vgnd vpwr scs8hd_decap_3
XANTENNA__230__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_259 vgnd vpwr scs8hd_decap_12
XFILLER_18_248 vgnd vpwr scs8hd_decap_8
XFILLER_18_226 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _184_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_130_ _119_/A _131_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_43 vpwr vgnd scs8hd_fill_2
XFILLER_23_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_218 vpwr vgnd scs8hd_fill_2
XANTENNA__225__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_133 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_34 vgnd vpwr scs8hd_decap_4
XFILLER_9_56 vgnd vpwr scs8hd_decap_3
XFILLER_20_210 vgnd vpwr scs8hd_decap_4
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_87 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd
+ vpwr scs8hd_diode_2
X_113_ address[3] _113_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_232 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_7_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vgnd vpwr scs8hd_decap_4
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_20_44 vgnd vpwr scs8hd_decap_3
XFILLER_20_22 vgnd vpwr scs8hd_decap_8
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_4_228 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_151 vpwr vgnd scs8hd_fill_2
XFILLER_6_24 vgnd vpwr scs8hd_fill_1
XFILLER_6_46 vgnd vpwr scs8hd_decap_4
XANTENNA__116__C _182_/C vgnd vpwr scs8hd_diode_2
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_4
XFILLER_19_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_198 vgnd vpwr scs8hd_decap_12
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_176 vgnd vpwr scs8hd_decap_6
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_22 vpwr vgnd scs8hd_fill_2
XFILLER_31_43 vgnd vpwr scs8hd_decap_12
XFILLER_31_32 vpwr vgnd scs8hd_fill_2
XFILLER_31_21 vgnd vpwr scs8hd_decap_4
XFILLER_31_10 vpwr vgnd scs8hd_fill_2
XFILLER_15_88 vgnd vpwr scs8hd_decap_4
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_231 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_5_ mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__127__B address[5] vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_157 vgnd vpwr scs8hd_decap_6
XFILLER_22_146 vgnd vpwr scs8hd_decap_6
XFILLER_7_9 vpwr vgnd scs8hd_fill_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_102 vpwr vgnd scs8hd_fill_2
XFILLER_13_113 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_138 vpwr vgnd scs8hd_fill_2
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_205 vgnd vpwr scs8hd_decap_8
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_241 vgnd vpwr scs8hd_decap_3
XFILLER_23_77 vgnd vpwr scs8hd_decap_4
XFILLER_23_55 vgnd vpwr scs8hd_decap_4
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XFILLER_2_101 vpwr vgnd scs8hd_fill_2
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_226 vpwr vgnd scs8hd_fill_2
X_112_ address[5] _162_/A vgnd vpwr scs8hd_buf_1
XANTENNA__236__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__146__A _145_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_29_10 vpwr vgnd scs8hd_fill_2
XFILLER_29_54 vgnd vpwr scs8hd_decap_6
XFILLER_29_32 vpwr vgnd scs8hd_fill_2
XFILLER_29_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XFILLER_31_55 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _217_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_133 vgnd vpwr scs8hd_decap_3
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _127_/C vgnd vpwr scs8hd_diode_2
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__244__A _244_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_180 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_106 vgnd vpwr scs8hd_decap_6
XFILLER_5_7 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _131_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _203_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_253 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_205 vpwr vgnd scs8hd_fill_2
XFILLER_7_249 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
X_111_ address[6] _161_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_245 vgnd vpwr scs8hd_decap_3
XFILLER_11_267 vgnd vpwr scs8hd_decap_8
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_260 vgnd vpwr scs8hd_decap_12
XFILLER_20_35 vpwr vgnd scs8hd_fill_2
XFILLER_29_66 vpwr vgnd scs8hd_fill_2
XFILLER_28_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_197 vgnd vpwr scs8hd_decap_4
XANTENNA__157__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_25_156 vgnd vpwr scs8hd_decap_4
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_244 vgnd vpwr scs8hd_fill_1
XFILLER_16_112 vpwr vgnd scs8hd_fill_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_6
XFILLER_16_167 vgnd vpwr scs8hd_decap_6
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_4
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_89 vgnd vpwr scs8hd_decap_3
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_108 vgnd vpwr scs8hd_decap_4
XFILLER_3_38 vgnd vpwr scs8hd_decap_4
XFILLER_3_16 vpwr vgnd scs8hd_fill_2
XFILLER_8_174 vpwr vgnd scs8hd_fill_2
XANTENNA__170__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_14 vpwr vgnd scs8hd_fill_2
XFILLER_12_36 vgnd vpwr scs8hd_decap_4
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_69 vpwr vgnd scs8hd_fill_2
XFILLER_18_218 vgnd vpwr scs8hd_decap_8
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _146_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_81 vgnd vpwr scs8hd_decap_4
XFILLER_23_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_221 vgnd vpwr scs8hd_fill_1
XFILLER_14_254 vgnd vpwr scs8hd_decap_4
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_79 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_68 vpwr vgnd scs8hd_fill_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_202 vpwr vgnd scs8hd_fill_2
XFILLER_11_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd
+ vpwr scs8hd_diode_2
X_110_ _104_/A _123_/A _110_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_239_ _239_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_250 vgnd vpwr scs8hd_fill_1
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_20_58 vpwr vgnd scs8hd_fill_2
XFILLER_29_45 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_28_143 vgnd vpwr scs8hd_decap_8
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_19_132 vgnd vpwr scs8hd_decap_4
XFILLER_20_8 vgnd vpwr scs8hd_decap_3
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_176 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA__083__A address[2] vgnd vpwr scs8hd_diode_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_127 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_26_46 vgnd vpwr scs8hd_decap_12
XFILLER_26_35 vgnd vpwr scs8hd_decap_4
XFILLER_13_149 vgnd vpwr scs8hd_decap_4
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vgnd vpwr scs8hd_decap_8
XFILLER_21_171 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__170__B _169_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_9_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_112 vgnd vpwr scs8hd_decap_4
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_252 vpwr vgnd scs8hd_fill_2
XFILLER_17_263 vpwr vgnd scs8hd_fill_2
XANTENNA__181__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_3
XFILLER_23_233 vgnd vpwr scs8hd_decap_8
XFILLER_23_222 vpwr vgnd scs8hd_fill_2
XFILLER_23_14 vgnd vpwr scs8hd_decap_3
XFILLER_23_47 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_2_137 vpwr vgnd scs8hd_fill_2
XFILLER_0_18 vgnd vpwr scs8hd_decap_12
XFILLER_9_38 vgnd vpwr scs8hd_fill_1
XFILLER_14_233 vgnd vpwr scs8hd_decap_8
X_186_ _178_/A _162_/A _164_/X _167_/A _186_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__176__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_258 vgnd vpwr scs8hd_decap_12
XFILLER_20_247 vgnd vpwr scs8hd_decap_8
XFILLER_20_236 vgnd vpwr scs8hd_decap_8
XFILLER_9_270 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_58 vgnd vpwr scs8hd_decap_4
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_236 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd
+ vpwr scs8hd_diode_2
X_169_ _169_/A _169_/X vgnd vpwr scs8hd_buf_1
X_238_ _238_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_240 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_7.LATCH_0_.latch data_in _194_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_254 vpwr vgnd scs8hd_fill_2
XFILLER_10_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_155 vpwr vgnd scs8hd_fill_2
XFILLER_19_90 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__173__B _169_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_136 vgnd vpwr scs8hd_decap_3
XFILLER_15_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_235 vgnd vpwr scs8hd_fill_1
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__168__B _162_/X vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__184__A _178_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XFILLER_26_58 vgnd vpwr scs8hd_fill_1
XFILLER_13_106 vpwr vgnd scs8hd_fill_2
XFILLER_13_117 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_29 vgnd vpwr scs8hd_decap_3
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
XANTENNA__170__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__089__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_17_231 vgnd vpwr scs8hd_decap_12
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__181__B _162_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_245 vgnd vpwr scs8hd_fill_1
XFILLER_23_26 vpwr vgnd scs8hd_fill_2
XFILLER_2_116 vpwr vgnd scs8hd_fill_2
XFILLER_2_105 vpwr vgnd scs8hd_fill_2
XANTENNA__091__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
XFILLER_9_28 vgnd vpwr scs8hd_decap_4
X_185_ _178_/A _162_/A _164_/X _165_/A _185_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
XFILLER_1_182 vgnd vpwr scs8hd_fill_1
XANTENNA__176__B _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XANTENNA__086__B _083_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_259 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _201_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_168_ _161_/X _162_/X _164_/X _167_/X _168_/Y vgnd vpwr scs8hd_nor4_4
X_237_ _237_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_270 vgnd vpwr scs8hd_decap_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_3
X_099_ _102_/A address[2] _165_/A _099_/X vgnd vpwr scs8hd_or3_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XANTENNA__097__A _104_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_0_.latch data_in _202_/A _184_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_266 vpwr vgnd scs8hd_fill_2
XFILLER_3_222 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__173__C _182_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_38 vpwr vgnd scs8hd_fill_2
XFILLER_0_269 vpwr vgnd scs8hd_fill_2
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XFILLER_0_203 vpwr vgnd scs8hd_fill_2
XFILLER_16_104 vgnd vpwr scs8hd_decap_8
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__C _164_/X vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__184__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_94 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_70 vgnd vpwr scs8hd_decap_3
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_133 vgnd vpwr scs8hd_decap_3
XANTENNA__170__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_199 vpwr vgnd scs8hd_fill_2
XANTENNA__179__B _162_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XANTENNA__089__B address[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _244_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_210 vgnd vpwr scs8hd_decap_4
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_27_91 vgnd vpwr scs8hd_fill_1
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
XANTENNA__181__C _182_/C vgnd vpwr scs8hd_diode_2
XFILLER_23_213 vgnd vpwr scs8hd_decap_6
XFILLER_23_202 vgnd vpwr scs8hd_decap_4
XANTENNA__091__C _137_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_11_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_184_ _178_/X _162_/A _127_/C _167_/A _184_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_71 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__176__C _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA__086__C _165_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_167_ _167_/A _167_/X vgnd vpwr scs8hd_buf_1
X_098_ address[1] _102_/A vgnd vpwr scs8hd_inv_8
X_236_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_39 vgnd vpwr scs8hd_decap_3
XANTENNA__097__B _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_168 vpwr vgnd scs8hd_fill_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__173__D _167_/X vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_3.LATCH_0_.latch data_in _190_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_160 vgnd vpwr scs8hd_decap_3
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XFILLER_22_108 vpwr vgnd scs8hd_fill_2
XANTENNA__168__D _167_/X vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA__184__C _127_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
XFILLER_15_193 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _204_/A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_152 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _215_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_145 vpwr vgnd scs8hd_fill_2
XFILLER_8_178 vpwr vgnd scs8hd_fill_2
XANTENNA__179__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_12_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XANTENNA__089__C _089_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XANTENNA__181__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_85 vgnd vpwr scs8hd_fill_1
XFILLER_4_74 vgnd vpwr scs8hd_decap_4
XFILLER_4_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _178_/X _162_/A _127_/C _165_/A _183_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA__176__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_206 vpwr vgnd scs8hd_fill_2
XFILLER_11_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
X_235_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_166_ _161_/X _162_/X _164_/X _165_/X _166_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_097_ _104_/A _119_/A _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_34_6 vgnd vpwr scs8hd_decap_8
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_103 vpwr vgnd scs8hd_fill_2
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ _131_/A _146_/X _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_117 vgnd vpwr scs8hd_decap_3
XFILLER_31_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_39 vpwr vgnd scs8hd_fill_2
XFILLER_31_28 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_227 vpwr vgnd scs8hd_fill_2
XFILLER_24_172 vgnd vpwr scs8hd_decap_8
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_11.LATCH_0_.latch data_in _198_/A _180_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XANTENNA__184__D _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_71 vgnd vpwr scs8hd_decap_12
XFILLER_8_113 vgnd vpwr scs8hd_fill_1
XFILLER_12_175 vgnd vpwr scs8hd_decap_3
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA__179__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_105 vgnd vpwr scs8hd_decap_4
XFILLER_5_138 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_267 vgnd vpwr scs8hd_decap_8
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_20 vpwr vgnd scs8hd_fill_2
XFILLER_4_171 vpwr vgnd scs8hd_fill_2
XFILLER_4_53 vgnd vpwr scs8hd_fill_1
XFILLER_23_226 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _178_/X _162_/X _182_/C _167_/A _182_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_215 vgnd vpwr scs8hd_decap_6
XFILLER_1_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__100__A _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
XFILLER_13_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
X_165_ _165_/A _165_/X vgnd vpwr scs8hd_buf_1
X_234_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_211 vgnd vpwr scs8hd_decap_3
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _095_/X _119_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_4
XFILLER_29_28 vpwr vgnd scs8hd_fill_2
XFILLER_29_17 vpwr vgnd scs8hd_fill_2
XFILLER_3_258 vgnd vpwr scs8hd_decap_4
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_10_41 vgnd vpwr scs8hd_decap_8
XFILLER_10_85 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XFILLER_27_170 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _199_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_148_ _119_/A _146_/X _148_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_3 vgnd vpwr scs8hd_fill_1
XFILLER_18_192 vgnd vpwr scs8hd_decap_4
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _156_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_73 vpwr vgnd scs8hd_fill_2
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_84 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_3_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_51 vpwr vgnd scs8hd_fill_2
XFILLER_16_84 vgnd vpwr scs8hd_decap_6
XFILLER_32_83 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _185_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_7_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _203_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_83 vpwr vgnd scs8hd_fill_2
XFILLER_27_72 vgnd vpwr scs8hd_decap_4
XFILLER_4_183 vpwr vgnd scs8hd_fill_2
XFILLER_4_98 vgnd vpwr scs8hd_decap_3
XFILLER_23_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_181_ _178_/X _162_/X _182_/C _165_/A _181_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_85 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_153 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_260 vpwr vgnd scs8hd_fill_2
XFILLER_18_19 vpwr vgnd scs8hd_fill_2
XFILLER_34_29 vpwr vgnd scs8hd_fill_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_164_ _163_/X _164_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_84 vgnd vpwr scs8hd_decap_3
XFILLER_24_62 vpwr vgnd scs8hd_fill_2
X_233_ _233_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_201 vpwr vgnd scs8hd_fill_2
XFILLER_6_223 vpwr vgnd scs8hd_fill_2
X_095_ address[1] _083_/Y _167_/A _095_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_241 vgnd vpwr scs8hd_decap_8
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_11 vpwr vgnd scs8hd_fill_2
XFILLER_1_99 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_64 vpwr vgnd scs8hd_fill_2
XFILLER_10_75 vgnd vpwr scs8hd_decap_4
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_51 vpwr vgnd scs8hd_fill_2
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_147_ _147_/A _146_/X _147_/Y vgnd vpwr scs8hd_nor2_4
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A _105_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
XFILLER_18_171 vgnd vpwr scs8hd_decap_6
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_207 vgnd vpwr scs8hd_decap_4
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_152 vpwr vgnd scs8hd_fill_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_98 vgnd vpwr scs8hd_decap_4
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_133 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_7_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _202_/A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_95 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XFILLER_17_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A _113_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_180_ _178_/X _162_/X _137_/C _167_/X _180_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_75 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_180 vgnd vpwr scs8hd_decap_3
XFILLER_24_74 vgnd vpwr scs8hd_fill_1
XFILLER_24_41 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_232_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_163_ _113_/Y _163_/B _089_/C _163_/X vgnd vpwr scs8hd_or3_4
X_094_ address[0] _167_/A vgnd vpwr scs8hd_buf_1
XFILLER_1_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_205 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
X_146_ _145_/X _146_/X vgnd vpwr scs8hd_buf_1
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_6 vgnd vpwr scs8hd_decap_8
XFILLER_18_161 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_24_197 vpwr vgnd scs8hd_fill_2
XFILLER_24_131 vpwr vgnd scs8hd_fill_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_120 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
X_129_ _147_/A _131_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_167 vpwr vgnd scs8hd_fill_2
XFILLER_21_145 vgnd vpwr scs8hd_decap_4
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _195_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_7.LATCH_1_.latch data_in _193_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_116 vpwr vgnd scs8hd_fill_2
XFILLER_8_138 vpwr vgnd scs8hd_fill_2
XFILLER_8_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_270 vgnd vpwr scs8hd_decap_4
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_26_204 vgnd vpwr scs8hd_decap_8
XFILLER_27_30 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__220__A _220_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_17_248 vpwr vgnd scs8hd_fill_2
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_78 vgnd vpwr scs8hd_fill_1
XFILLER_4_45 vgnd vpwr scs8hd_decap_8
XFILLER_22_251 vgnd vpwr scs8hd_decap_8
XFILLER_22_240 vgnd vpwr scs8hd_decap_8
XFILLER_22_262 vgnd vpwr scs8hd_decap_12
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XFILLER_9_222 vpwr vgnd scs8hd_fill_2
XFILLER_9_266 vpwr vgnd scs8hd_fill_2
XFILLER_13_240 vgnd vpwr scs8hd_fill_1
XANTENNA__125__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_162_ _162_/A _162_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_97 vgnd vpwr scs8hd_fill_1
XFILLER_24_20 vpwr vgnd scs8hd_fill_2
X_231_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _147_/A _104_/A _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_79 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_107 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_11 vgnd vpwr scs8hd_fill_1
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_19_86 vpwr vgnd scs8hd_fill_2
XFILLER_19_75 vgnd vpwr scs8hd_decap_6
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _178_/A _169_/A _182_/C _145_/X vgnd vpwr scs8hd_or3_4
XANTENNA__122__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _205_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XFILLER_21_21 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_32 vpwr vgnd scs8hd_fill_2
XANTENNA__223__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _122_/A vgnd vpwr scs8hd_diode_2
X_128_ _127_/X _131_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _197_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_16_10 vgnd vpwr scs8hd_fill_1
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_1_.latch data_in _201_/A _183_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_109 vgnd vpwr scs8hd_fill_1
XFILLER_17_227 vpwr vgnd scs8hd_fill_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_24 vgnd vpwr scs8hd_decap_4
XANTENNA__114__C _089_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_175 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_57 vgnd vpwr scs8hd_decap_6
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _201_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_22 vpwr vgnd scs8hd_fill_2
XFILLER_1_178 vpwr vgnd scs8hd_fill_2
XFILLER_1_156 vgnd vpwr scs8hd_fill_1
XFILLER_1_112 vpwr vgnd scs8hd_fill_2
XANTENNA__231__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _131_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_160 vgnd vpwr scs8hd_decap_12
X_161_ _161_/A _161_/X vgnd vpwr scs8hd_buf_1
XANTENNA__226__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
X_230_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_092_ _091_/X _104_/A vgnd vpwr scs8hd_buf_1
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_28_119 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_218 vpwr vgnd scs8hd_fill_2
XFILLER_10_23 vgnd vpwr scs8hd_decap_8
XFILLER_10_89 vgnd vpwr scs8hd_fill_1
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
X_144_ _123_/A _138_/X _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_130 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_111 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_90 vpwr vgnd scs8hd_fill_2
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_88 vgnd vpwr scs8hd_decap_3
XFILLER_21_77 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_133 vpwr vgnd scs8hd_fill_2
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_24 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_79 vpwr vgnd scs8hd_fill_2
X_127_ address[6] address[5] _127_/C _127_/X vgnd vpwr scs8hd_or3_4
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _246_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vgnd vpwr scs8hd_decap_6
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_20_191 vgnd vpwr scs8hd_decap_4
XANTENNA__234__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_129 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_87 vgnd vpwr scs8hd_decap_4
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_217 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_3.LATCH_1_.latch data_in _189_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_187 vpwr vgnd scs8hd_fill_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_209 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XFILLER_13_89 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _200_/A mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__125__C _089_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_235 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_172 vgnd vpwr scs8hd_decap_8
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_66 vgnd vpwr scs8hd_decap_8
X_160_ _123_/A _154_/X _160_/Y vgnd vpwr scs8hd_nor2_4
X_091_ address[6] address[5] _137_/C _091_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_205 vgnd vpwr scs8hd_decap_4
XFILLER_6_227 vpwr vgnd scs8hd_fill_2
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_fill_1
XANTENNA__152__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_55 vgnd vpwr scs8hd_decap_4
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_143_ _122_/A _138_/X _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_2_241 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _204_/Y mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_189 vgnd vpwr scs8hd_decap_8
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_1_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_126_ _125_/X _127_/C vgnd vpwr scs8hd_buf_1
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_6 vgnd vpwr scs8hd_decap_8
XFILLER_21_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_23 vgnd vpwr scs8hd_decap_4
XFILLER_12_104 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_174 vgnd vpwr scs8hd_decap_3
XANTENNA__144__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _123_/A vgnd vpwr scs8hd_diode_2
X_109_ _108_/X _123_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_99 vpwr vgnd scs8hd_fill_2
XFILLER_27_44 vpwr vgnd scs8hd_fill_2
XFILLER_25_262 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _193_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__245__A _245_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_133 vpwr vgnd scs8hd_fill_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_11.LATCH_1_.latch data_in _197_/A _179_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_79 vgnd vpwr scs8hd_decap_3
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_203 vpwr vgnd scs8hd_fill_2
XFILLER_13_221 vgnd vpwr scs8hd_decap_3
XFILLER_13_243 vgnd vpwr scs8hd_fill_1
XFILLER_13_254 vgnd vpwr scs8hd_decap_4
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_258 vgnd vpwr scs8hd_decap_4
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_24_89 vgnd vpwr scs8hd_decap_3
X_090_ _089_/X _137_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__152__B _146_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_261 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ _190_/A mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_58 vgnd vpwr scs8hd_decap_4
XFILLER_27_154 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_27_110 vgnd vpwr scs8hd_decap_12
XFILLER_19_34 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
X_142_ _150_/A _138_/X _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_8 vpwr vgnd scs8hd_fill_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B _146_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_4
XANTENNA__163__A _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XFILLER_24_135 vgnd vpwr scs8hd_fill_1
XFILLER_24_124 vgnd vpwr scs8hd_decap_4
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_113 vgnd vpwr scs8hd_fill_1
XFILLER_15_146 vgnd vpwr scs8hd_decap_4
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
X_125_ address[3] _163_/B _089_/C _125_/X vgnd vpwr scs8hd_or3_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_90 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_23_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_149 vgnd vpwr scs8hd_fill_1
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_190 vpwr vgnd scs8hd_fill_2
XFILLER_16_13 vgnd vpwr scs8hd_fill_1
XFILLER_12_149 vpwr vgnd scs8hd_fill_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd
+ vpwr scs8hd_diode_2
X_108_ address[1] address[2] address[0] _108_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_153 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_4
XANTENNA__160__B _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_34 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_56 vgnd vpwr scs8hd_decap_4
XFILLER_25_274 vgnd vpwr scs8hd_decap_3
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _155_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_112 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _206_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_92 vgnd vpwr scs8hd_fill_1
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_24_24 vpwr vgnd scs8hd_fill_2
XFILLER_10_203 vgnd vpwr scs8hd_decap_4
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _207_/HI _199_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _196_/A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _131_/A _138_/X _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_188 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_114 vgnd vpwr scs8hd_fill_1
XFILLER_2_60 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_36 vpwr vgnd scs8hd_fill_2
XFILLER_21_25 vpwr vgnd scs8hd_fill_2
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_191 vgnd vpwr scs8hd_decap_4
X_124_ address[4] _163_/B vgnd vpwr scs8hd_inv_8
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_6 vgnd vpwr scs8hd_decap_4
XANTENNA__174__A _161_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_36 vpwr vgnd scs8hd_fill_2
XFILLER_16_47 vpwr vgnd scs8hd_fill_2
XFILLER_32_35 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_139 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_150 vpwr vgnd scs8hd_fill_2
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
X_107_ _104_/A _122_/A _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_6
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_68 vpwr vgnd scs8hd_fill_2
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XFILLER_25_242 vpwr vgnd scs8hd_fill_2
XFILLER_4_28 vgnd vpwr scs8hd_fill_1
XFILLER_16_220 vpwr vgnd scs8hd_fill_2
XFILLER_16_231 vgnd vpwr scs8hd_decap_12
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__171__B _169_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_26 vpwr vgnd scs8hd_fill_2
XFILLER_1_149 vgnd vpwr scs8hd_decap_4
XFILLER_1_116 vgnd vpwr scs8hd_decap_4
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _162_/X vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_219 vpwr vgnd scs8hd_fill_2
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_90 vpwr vgnd scs8hd_fill_2
XFILLER_5_241 vgnd vpwr scs8hd_fill_1
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _161_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _198_/A mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_6
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_140_ _119_/A _138_/X _140_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_211 vgnd vpwr scs8hd_decap_3
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _089_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_83 vgnd vpwr scs8hd_fill_1
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_123_ _123_/A _118_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_28 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__174__B _169_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _202_/Y mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_262 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_129 vpwr vgnd scs8hd_fill_2
XFILLER_32_47 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
X_106_ _105_/X _122_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_166 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_fill_1
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_82 vgnd vpwr scs8hd_fill_1
XFILLER_25_210 vgnd vpwr scs8hd_decap_12
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_243 vgnd vpwr scs8hd_fill_1
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _137_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_38 vgnd vpwr scs8hd_decap_4
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_202 vpwr vgnd scs8hd_fill_2
XFILLER_9_239 vgnd vpwr scs8hd_decap_3
XFILLER_0_161 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_3_ mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C _164_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _191_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__182__B _162_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_19 vpwr vgnd scs8hd_fill_2
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XANTENNA__177__B _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_245 vgnd vpwr scs8hd_decap_4
XFILLER_2_201 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_149 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _195_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
XFILLER_15_116 vpwr vgnd scs8hd_fill_2
XFILLER_23_182 vgnd vpwr scs8hd_fill_1
XFILLER_23_171 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ _188_/A mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_122_ _122_/A _118_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_108 vgnd vpwr scs8hd_decap_4
XANTENNA__174__C _127_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_182 vpwr vgnd scs8hd_fill_2
XFILLER_37_274 vgnd vpwr scs8hd_decap_3
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_fill_1
XFILLER_32_59 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_174 vpwr vgnd scs8hd_fill_2
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_105_ address[1] address[2] _085_/A _105_/X vgnd vpwr scs8hd_or3_4
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XANTENNA__185__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_61 vpwr vgnd scs8hd_fill_2
XFILLER_27_48 vgnd vpwr scs8hd_decap_6
XFILLER_27_37 vgnd vpwr scs8hd_decap_4
XFILLER_27_26 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vpwr vgnd scs8hd_fill_2
XFILLER_25_222 vgnd vpwr scs8hd_decap_12
XANTENNA__095__B _083_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_137 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_211 vgnd vpwr scs8hd_decap_3
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__171__D _167_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_15_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_203 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_236 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XANTENNA__166__D _165_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_51 vpwr vgnd scs8hd_fill_2
XANTENNA__182__C _182_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_95 vgnd vpwr scs8hd_fill_1
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_228 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_70 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_210 vpwr vgnd scs8hd_fill_2
XFILLER_5_265 vgnd vpwr scs8hd_decap_12
XANTENNA__177__C _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_158 vgnd vpwr scs8hd_decap_12
XFILLER_27_136 vgnd vpwr scs8hd_decap_12
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_224 vgnd vpwr scs8hd_decap_3
XFILLER_26_180 vgnd vpwr scs8hd_decap_12
XFILLER_18_158 vgnd vpwr scs8hd_fill_1
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_96 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _206_/HI _197_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_128 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _194_/A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_121_ _150_/A _118_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA__174__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_194 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_102 vgnd vpwr scs8hd_fill_1
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_120 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
X_104_ _104_/A _150_/A _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_7 vgnd vpwr scs8hd_fill_1
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__185__C _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
XFILLER_25_234 vgnd vpwr scs8hd_decap_8
XANTENNA__095__C _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_116 vpwr vgnd scs8hd_fill_2
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _216_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_226 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _207_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__182__D _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_6
XFILLER_24_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_50 vgnd vpwr scs8hd_fill_1
XFILLER_14_83 vgnd vpwr scs8hd_decap_6
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_82 vgnd vpwr scs8hd_decap_8
XFILLER_5_233 vpwr vgnd scs8hd_fill_2
XANTENNA__177__D _167_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_5_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_148 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_104 vpwr vgnd scs8hd_fill_2
XFILLER_2_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_192 vgnd vpwr scs8hd_decap_12
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_107 vgnd vpwr scs8hd_decap_4
XFILLER_2_86 vpwr vgnd scs8hd_fill_2
XFILLER_2_64 vgnd vpwr scs8hd_fill_1
XFILLER_15_129 vpwr vgnd scs8hd_fill_2
X_120_ _131_/A _118_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_17 vgnd vpwr scs8hd_decap_12
XFILLER_20_198 vgnd vpwr scs8hd_decap_12
XFILLER_20_187 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vgnd vpwr scs8hd_decap_3
XFILLER_22_72 vgnd vpwr scs8hd_fill_1
X_103_ _102_/X _150_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_154 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_221 vpwr vgnd scs8hd_fill_2
XFILLER_8_41 vpwr vgnd scs8hd_fill_2
XFILLER_8_85 vgnd vpwr scs8hd_decap_4
XANTENNA__185__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _200_/Y mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_142 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_220 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_62 vpwr vgnd scs8hd_fill_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_4
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _189_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_149 vgnd vpwr scs8hd_decap_4
XFILLER_18_138 vgnd vpwr scs8hd_decap_4
XFILLER_18_116 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_25_83 vpwr vgnd scs8hd_fill_2
XFILLER_25_72 vgnd vpwr scs8hd_decap_4
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_43 vpwr vgnd scs8hd_fill_2
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
XFILLER_1_270 vgnd vpwr scs8hd_decap_6
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_152 vgnd vpwr scs8hd_fill_1
XFILLER_14_163 vpwr vgnd scs8hd_fill_2
X_179_ _178_/X _162_/X _137_/C _165_/X _179_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _193_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
X_102_ _102_/A address[2] _167_/A _102_/X vgnd vpwr scs8hd_or3_4
XFILLER_34_258 vgnd vpwr scs8hd_decap_12
XFILLER_8_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_258 vpwr vgnd scs8hd_fill_2
XFILLER_4_129 vpwr vgnd scs8hd_fill_2
XFILLER_16_203 vpwr vgnd scs8hd_fill_2
XFILLER_16_247 vgnd vpwr scs8hd_decap_8
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_173 vgnd vpwr scs8hd_decap_4
XFILLER_3_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_206 vpwr vgnd scs8hd_fill_2
XFILLER_21_250 vgnd vpwr scs8hd_decap_4
XFILLER_28_50 vgnd vpwr scs8hd_decap_4
XFILLER_0_187 vgnd vpwr scs8hd_fill_1
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_243 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in _196_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_136 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _190_/Y mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_209 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__101__B _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_106 vpwr vgnd scs8hd_fill_2
XFILLER_19_19 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_205 vgnd vpwr scs8hd_decap_4
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_175 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_109 vgnd vpwr scs8hd_decap_4
XFILLER_11_42 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_86 vpwr vgnd scs8hd_fill_2
XFILLER_14_131 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_142 vpwr vgnd scs8hd_fill_2
XFILLER_14_186 vpwr vgnd scs8hd_fill_2
X_178_ _178_/A _178_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_145 vgnd vpwr scs8hd_decap_8
XFILLER_22_52 vgnd vpwr scs8hd_fill_1
XFILLER_22_41 vgnd vpwr scs8hd_decap_3
X_101_ _104_/A _131_/A _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_149 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _192_/A mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_19 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_3
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XFILLER_17_41 vgnd vpwr scs8hd_decap_3
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _150_/A vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_229 vgnd vpwr scs8hd_decap_8
XFILLER_22_218 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_15_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _186_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_1_ mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_262 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_211 vgnd vpwr scs8hd_fill_1
XFILLER_12_240 vgnd vpwr scs8hd_fill_1
XFILLER_12_262 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _114_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_11 vgnd vpwr scs8hd_decap_3
XFILLER_5_44 vgnd vpwr scs8hd_decap_4
XFILLER_5_55 vgnd vpwr scs8hd_decap_4
XFILLER_39_148 vgnd vpwr scs8hd_decap_12
XFILLER_5_88 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _196_/Y mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _204_/A _186_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_20 vpwr vgnd scs8hd_fill_2
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_151 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XFILLER_25_52 vgnd vpwr scs8hd_decap_6
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_67 vgnd vpwr scs8hd_fill_1
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_162 vpwr vgnd scs8hd_fill_2
XFILLER_17_173 vpwr vgnd scs8hd_fill_2
XFILLER_23_198 vpwr vgnd scs8hd_fill_2
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _183_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_110 vgnd vpwr scs8hd_fill_1
X_246_ _246_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B _122_/A vgnd vpwr scs8hd_diode_2
X_177_ _161_/A _169_/A _164_/X _167_/X _177_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
XFILLER_22_64 vgnd vpwr scs8hd_decap_8
XFILLER_11_113 vgnd vpwr scs8hd_fill_1
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
X_100_ _099_/X _131_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _147_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_172 vpwr vgnd scs8hd_fill_2
X_229_ _229_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_13_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_20 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_21_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_fill_1
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XANTENNA__221__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_96 vgnd vpwr scs8hd_decap_8
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _198_/Y mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_11_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_237 vgnd vpwr scs8hd_decap_4
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A _125_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_0_.latch data_in _192_/A _173_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_229 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_18_108 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_79 vgnd vpwr scs8hd_decap_4
XFILLER_2_13 vgnd vpwr scs8hd_decap_3
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_141 vgnd vpwr scs8hd_fill_1
XFILLER_23_100 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_133 vgnd vpwr scs8hd_decap_3
XFILLER_11_22 vgnd vpwr scs8hd_decap_4
XFILLER_11_66 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _187_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_245_ _245_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_176_ _161_/A _169_/A _164_/X _165_/X _176_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__123__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_258 vpwr vgnd scs8hd_fill_2
XFILLER_20_158 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_21 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA__224__A _224_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_19_225 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_45 vgnd vpwr scs8hd_decap_3
XANTENNA__134__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr
+ scs8hd_diode_2
X_228_ _228_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
X_159_ _122_/A _154_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_78 vgnd vpwr scs8hd_decap_4
XFILLER_8_89 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _147_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_261 vgnd vpwr scs8hd_decap_12
XANTENNA__129__A _147_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _191_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_102 vpwr vgnd scs8hd_fill_2
XFILLER_8_224 vpwr vgnd scs8hd_fill_2
XFILLER_8_257 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_66 vgnd vpwr scs8hd_decap_4
XFILLER_5_249 vgnd vpwr scs8hd_fill_1
XANTENNA__232__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _150_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_131 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _205_/HI _188_/Y mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmem_bottom_track_13.LATCH_0_.latch data_in _200_/A _182_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_2_47 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_fill_1
XFILLER_23_178 vpwr vgnd scs8hd_fill_2
XFILLER_23_167 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _219_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_7 vgnd vpwr scs8hd_decap_4
X_244_ _244_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_14_167 vgnd vpwr scs8hd_decap_4
X_175_ _161_/A _169_/X _127_/C _167_/X _175_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_137 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_204 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_24 vgnd vpwr scs8hd_decap_4
X_227_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__134__B _131_/B vgnd vpwr scs8hd_diode_2
X_089_ address[3] address[4] _089_/C _089_/X vgnd vpwr scs8hd_or3_4
X_158_ _150_/A _154_/X _158_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_207 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_33_21 vpwr vgnd scs8hd_fill_2
XFILLER_33_10 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_273 vpwr vgnd scs8hd_fill_2
XANTENNA__235__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _178_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _190_/A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_254 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_65 vgnd vpwr scs8hd_fill_1
XFILLER_28_32 vgnd vpwr scs8hd_decap_3
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_8_203 vpwr vgnd scs8hd_fill_2
XFILLER_8_247 vgnd vpwr scs8hd_fill_1
XFILLER_8_269 vgnd vpwr scs8hd_decap_6
XFILLER_12_232 vgnd vpwr scs8hd_decap_8
XFILLER_12_243 vpwr vgnd scs8hd_fill_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_25 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_89 vgnd vpwr scs8hd_fill_1
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA__142__B _138_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _218_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _194_/Y mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_121 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_143 vgnd vpwr scs8hd_decap_8
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA__137__B _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__153__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_46 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_0_.latch data_in _188_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_102 vpwr vgnd scs8hd_fill_2
X_243_ _243_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_14_135 vpwr vgnd scs8hd_fill_2
XFILLER_14_146 vgnd vpwr scs8hd_decap_6
X_174_ _161_/A _169_/X _127_/C _165_/X _174_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__148__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_161 vpwr vgnd scs8hd_fill_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_11_105 vpwr vgnd scs8hd_fill_2
XFILLER_11_116 vpwr vgnd scs8hd_fill_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_19_249 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_226_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
X_157_ _131_/A _154_/X _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_182 vpwr vgnd scs8hd_fill_2
XANTENNA__150__B _146_/X vgnd vpwr scs8hd_diode_2
X_088_ enable _089_/C vgnd vpwr scs8hd_inv_8
XFILLER_6_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XFILLER_18_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_123 vgnd vpwr scs8hd_fill_1
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_115 vpwr vgnd scs8hd_fill_2
XANTENNA__246__A _246_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_215 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_48 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_7 vpwr vgnd scs8hd_fill_2
XANTENNA__156__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XFILLER_14_24 vgnd vpwr scs8hd_decap_4
XFILLER_5_229 vpwr vgnd scs8hd_fill_2
XFILLER_14_46 vpwr vgnd scs8hd_fill_2
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_262 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_254 vpwr vgnd scs8hd_fill_2
XFILLER_1_221 vpwr vgnd scs8hd_fill_2
XFILLER_17_144 vgnd vpwr scs8hd_decap_4
XFILLER_17_166 vpwr vgnd scs8hd_fill_2
XFILLER_17_177 vgnd vpwr scs8hd_decap_4
XANTENNA__137__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _169_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_15_ mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_191 vgnd vpwr scs8hd_decap_8
X_173_ _161_/X _169_/X _182_/C _167_/X _173_/Y vgnd vpwr scs8hd_nor4_4
X_242_ _242_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_128 vgnd vpwr scs8hd_decap_8
XANTENNA__148__B _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_46 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_225_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_154 vgnd vpwr scs8hd_fill_1
XFILLER_6_176 vpwr vgnd scs8hd_fill_2
X_156_ _119_/A _154_/X _156_/Y vgnd vpwr scs8hd_nor2_4
X_087_ _087_/A _147_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_24 vpwr vgnd scs8hd_fill_2
XFILLER_17_46 vpwr vgnd scs8hd_fill_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__145__C _182_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
X_139_ _147_/A _138_/X _139_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_245 vgnd vpwr scs8hd_decap_3
XFILLER_21_234 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__172__A _161_/X vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _189_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _245_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_46 vgnd vpwr scs8hd_decap_12
XFILLER_30_35 vgnd vpwr scs8hd_decap_8
XFILLER_39_22 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_241 vpwr vgnd scs8hd_fill_2
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_24 vpwr vgnd scs8hd_fill_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_68 vpwr vgnd scs8hd_fill_2
XFILLER_1_266 vpwr vgnd scs8hd_fill_2
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XANTENNA__153__C _127_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_26 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_9.LATCH_1_.latch data_in _195_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
X_172_ _161_/X _169_/X _182_/C _165_/X _172_/Y vgnd vpwr scs8hd_nor4_4
X_241_ _241_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_107 vgnd vpwr scs8hd_decap_12
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XANTENNA__180__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_82 vpwr vgnd scs8hd_fill_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_25 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_7 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _089_/X vgnd vpwr scs8hd_diode_2
X_224_ _224_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
X_086_ address[1] _083_/Y _165_/A _087_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_133 vgnd vpwr scs8hd_fill_1
X_155_ _147_/A _154_/X _155_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _161_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_221 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_169 vpwr vgnd scs8hd_fill_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
X_207_ _207_/HI _207_/LO vgnd vpwr scs8hd_conb_1
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_138_ _137_/X _138_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
XFILLER_9_92 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_57 vgnd vpwr scs8hd_decap_8
XFILLER_8_239 vpwr vgnd scs8hd_fill_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _169_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_261 vpwr vgnd scs8hd_fill_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_30_58 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _188_/A mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_39_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__183__A _178_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_168 vgnd vpwr scs8hd_decap_12
XFILLER_26_157 vgnd vpwr scs8hd_decap_6
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XFILLER_25_58 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_201 vpwr vgnd scs8hd_fill_2
XFILLER_2_18 vpwr vgnd scs8hd_fill_2
XFILLER_17_113 vpwr vgnd scs8hd_fill_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_138 vgnd vpwr scs8hd_decap_3
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_16_190 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A enable vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
X_171_ _161_/X _169_/X _137_/C _167_/X _171_/Y vgnd vpwr scs8hd_nor4_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _192_/Y mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in _203_/A _185_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_153 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XANTENNA__180__B _162_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_19_208 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_223_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_8_28 vgnd vpwr scs8hd_fill_1
X_154_ _154_/A _154_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
X_085_ _085_/A _165_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
XFILLER_10_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__175__B _169_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_37 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_25 vgnd vpwr scs8hd_decap_12
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_148 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_266 vpwr vgnd scs8hd_fill_2
X_206_ _206_/HI _206_/LO vgnd vpwr scs8hd_conb_1
X_137_ _178_/A _169_/A _137_/C _137_/X vgnd vpwr scs8hd_or3_4
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XFILLER_21_258 vpwr vgnd scs8hd_fill_2
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XANTENNA__186__A _178_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _220_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_69 vgnd vpwr scs8hd_decap_8
XANTENNA__096__A _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_207 vgnd vpwr scs8hd_decap_4
XFILLER_12_247 vpwr vgnd scs8hd_fill_2
XFILLER_12_258 vpwr vgnd scs8hd_fill_2
XFILLER_5_29 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__172__C _182_/C vgnd vpwr scs8hd_diode_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_46 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _224_/A vgnd vpwr scs8hd_inv_1
XANTENNA__183__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_72 vgnd vpwr scs8hd_fill_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_125 vgnd vpwr scs8hd_decap_4
XFILLER_25_48 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__093__B _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_191 vgnd vpwr scs8hd_decap_4
XFILLER_15_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_170_ _161_/X _169_/X _137_/C _165_/X _170_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_106 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_9_165 vgnd vpwr scs8hd_fill_1
XANTENNA__180__C _137_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_4
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_109 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_1_.latch data_in _191_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_102 vgnd vpwr scs8hd_decap_3
X_222_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_10_120 vgnd vpwr scs8hd_decap_3
X_153_ _178_/A _169_/A _127_/C _154_/A vgnd vpwr scs8hd_or3_4
X_084_ address[0] _085_/A vgnd vpwr scs8hd_inv_8
XFILLER_26_8 vgnd vpwr scs8hd_decap_3
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
XANTENNA__175__C _127_/C vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_37 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
X_205_ _205_/HI _205_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_81 vgnd vpwr scs8hd_fill_1
X_136_ address[5] _169_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_171 vgnd vpwr scs8hd_decap_3
XFILLER_0_30 vgnd vpwr scs8hd_fill_1
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA__186__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_226 vpwr vgnd scs8hd_fill_2
XFILLER_21_215 vpwr vgnd scs8hd_fill_2
XFILLER_21_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_15 vpwr vgnd scs8hd_fill_2
XFILLER_0_119 vgnd vpwr scs8hd_decap_3
XFILLER_12_215 vgnd vpwr scs8hd_decap_4
XFILLER_20_270 vgnd vpwr scs8hd_decap_4
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ _119_/A _118_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__172__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_230 vpwr vgnd scs8hd_fill_2
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_28 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__183__C _127_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _187_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_1_258 vgnd vpwr scs8hd_decap_4
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_1_225 vpwr vgnd scs8hd_fill_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_137 vgnd vpwr scs8hd_decap_4
XFILLER_17_148 vgnd vpwr scs8hd_fill_1
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_18 vpwr vgnd scs8hd_fill_2
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_262 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_188 vpwr vgnd scs8hd_fill_2
XFILLER_9_199 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__180__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
X_083_ address[2] _083_/Y vgnd vpwr scs8hd_inv_8
X_152_ _123_/A _146_/X _152_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_125 vpwr vgnd scs8hd_fill_2
X_221_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_232 vgnd vpwr scs8hd_decap_12
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA__175__D _167_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_13.LATCH_1_.latch data_in _199_/A _181_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_33_49 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_235 vgnd vpwr scs8hd_decap_3
XFILLER_23_93 vgnd vpwr scs8hd_decap_4
XFILLER_23_71 vgnd vpwr scs8hd_decap_4
X_135_ address[6] _178_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__186__C _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_95 vpwr vgnd scs8hd_fill_2
XFILLER_28_38 vgnd vpwr scs8hd_decap_12
XFILLER_12_205 vpwr vgnd scs8hd_fill_2
XFILLER_7_220 vgnd vpwr scs8hd_decap_4
X_118_ _147_/A _118_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_4
XFILLER_30_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_9_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_4_245 vgnd vpwr scs8hd_decap_4
XFILLER_29_70 vgnd vpwr scs8hd_decap_12
XFILLER_35_127 vgnd vpwr scs8hd_fill_1
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vgnd vpwr scs8hd_decap_3
XFILLER_6_52 vgnd vpwr scs8hd_fill_1
XANTENNA__183__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_138 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_28 vgnd vpwr scs8hd_decap_4
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_13_ mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_7 vpwr vgnd scs8hd_fill_2
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_25_160 vgnd vpwr scs8hd_fill_1
XFILLER_17_105 vgnd vpwr scs8hd_decap_4
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_174 vgnd vpwr scs8hd_decap_8
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_174 vgnd vpwr scs8hd_decap_3
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XANTENNA__099__C _165_/A vgnd vpwr scs8hd_diode_2
X_220_ _220_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
X_151_ _122_/A _146_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_40 vgnd vpwr scs8hd_fill_1
XFILLER_12_84 vgnd vpwr scs8hd_decap_6
XFILLER_18_244 vgnd vpwr scs8hd_fill_1
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _190_/Y mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_33_17 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_225 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _214_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_214 vpwr vgnd scs8hd_fill_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_258 vgnd vpwr scs8hd_decap_4
X_134_ _123_/A _131_/B _134_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_7 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in _187_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
XANTENNA__186__D _167_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_52 vpwr vgnd scs8hd_fill_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_117_ _117_/A _118_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_265 vgnd vpwr scs8hd_decap_12
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XFILLER_30_29 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
XFILLER_4_202 vpwr vgnd scs8hd_fill_2
XFILLER_4_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_82 vgnd vpwr scs8hd_decap_12
XFILLER_29_60 vgnd vpwr scs8hd_fill_1
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_20 vgnd vpwr scs8hd_decap_4
XFILLER_6_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_106 vgnd vpwr scs8hd_decap_6
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_205 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_117 vgnd vpwr scs8hd_decap_3
XFILLER_25_172 vpwr vgnd scs8hd_fill_2
XFILLER_25_150 vgnd vpwr scs8hd_decap_4
XFILLER_15_95 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
XFILLER_22_142 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_83 vgnd vpwr scs8hd_decap_4
XFILLER_9_157 vpwr vgnd scs8hd_fill_2
XFILLER_13_153 vgnd vpwr scs8hd_fill_1
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _150_/A _146_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_167 vpwr vgnd scs8hd_fill_2
XFILLER_10_178 vpwr vgnd scs8hd_fill_2
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_12_52 vpwr vgnd scs8hd_fill_2
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XFILLER_24_237 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_51 vpwr vgnd scs8hd_fill_2
X_133_ _122_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_11 vgnd vpwr scs8hd_decap_4
XANTENNA__110__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__105__A address[1] vgnd vpwr scs8hd_diode_2
X_116_ _161_/A _162_/A _182_/C _117_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_20_30 vgnd vpwr scs8hd_fill_1
XFILLER_4_258 vpwr vgnd scs8hd_fill_2
XFILLER_29_94 vgnd vpwr scs8hd_decap_12
XFILLER_29_50 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_13_121 vgnd vpwr scs8hd_fill_1
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_99 vpwr vgnd scs8hd_fill_2
XFILLER_3_66 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_102 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_249 vgnd vpwr scs8hd_decap_12
X_132_ _150_/A _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_260 vgnd vpwr scs8hd_decap_12
XFILLER_23_30 vpwr vgnd scs8hd_fill_2
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_197 vpwr vgnd scs8hd_fill_2
XFILLER_2_120 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _123_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_219 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_19 vgnd vpwr scs8hd_decap_12
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_20_230 vgnd vpwr scs8hd_decap_3
XFILLER_18_41 vgnd vpwr scs8hd_decap_6
X_115_ _114_/X _182_/C vgnd vpwr scs8hd_buf_1
XANTENNA__105__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_201 vpwr vgnd scs8hd_fill_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_4
XFILLER_11_263 vpwr vgnd scs8hd_fill_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__121__A _150_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vgnd vpwr scs8hd_fill_1
XFILLER_20_97 vgnd vpwr scs8hd_fill_1
XFILLER_20_75 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_270 vgnd vpwr scs8hd_decap_6
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_3
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_229 vgnd vpwr scs8hd_decap_3
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_42 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_273 vpwr vgnd scs8hd_fill_2
XFILLER_0_262 vpwr vgnd scs8hd_fill_2
XFILLER_0_240 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__C _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
.ends

