VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_right
  CLASS BLOCK ;
  FOREIGN grid_io_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 187.920 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 2.400 ;
    END
  END ccff_tail
  PIN gfpga_pad_GPIO_A
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 24.520 80.000 25.120 ;
    END
  END gfpga_pad_GPIO_A
  PIN gfpga_pad_GPIO_IE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 74.160 80.000 74.760 ;
    END
  END gfpga_pad_GPIO_IE
  PIN gfpga_pad_GPIO_OE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 124.480 80.000 125.080 ;
    END
  END gfpga_pad_GPIO_OE
  PIN gfpga_pad_GPIO_Y
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 174.120 80.000 174.720 ;
    END
  END gfpga_pad_GPIO_Y
  PIN left_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END left_width_0_height_0__pin_0_
  PIN left_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END left_width_0_height_0__pin_1_lower
  PIN left_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.400 167.240 ;
    END
  END left_width_0_height_0__pin_1_upper
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 2.400 ;
    END
  END prog_clk
  PIN vpwr
    USE POWER ; 
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ; 
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 74.060 187.920 ;
      LAYER met2 ;
        RECT 6.990 2.680 72.925 187.920 ;
        RECT 6.990 2.400 13.150 2.680 ;
        RECT 13.990 2.400 39.830 2.680 ;
        RECT 40.670 2.400 66.510 2.680 ;
        RECT 67.350 2.400 72.925 2.680 ;
      LAYER met3 ;
        RECT 2.400 175.120 77.600 187.845 ;
        RECT 2.400 173.720 77.200 175.120 ;
        RECT 2.400 167.640 77.600 173.720 ;
        RECT 2.800 166.240 77.600 167.640 ;
        RECT 2.400 125.480 77.600 166.240 ;
        RECT 2.400 124.080 77.200 125.480 ;
        RECT 2.400 101.000 77.600 124.080 ;
        RECT 2.800 99.600 77.600 101.000 ;
        RECT 2.400 75.160 77.600 99.600 ;
        RECT 2.400 73.760 77.200 75.160 ;
        RECT 2.400 34.360 77.600 73.760 ;
        RECT 2.800 32.960 77.600 34.360 ;
        RECT 2.400 25.520 77.600 32.960 ;
        RECT 2.400 24.120 77.200 25.520 ;
        RECT 2.400 9.695 77.600 24.120 ;
      LAYER met4 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END grid_io_right
END LIBRARY

