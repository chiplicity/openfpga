* NGSPICE file created from sb_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

.subckt sb_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_11_ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ left_top_grid_pin_10_ right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_
+ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_
+ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ vpwr vgnd
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_30 vgnd vpwr scs8hd_fill_1
XFILLER_13_100 vpwr vgnd scs8hd_fill_2
XFILLER_9_104 vgnd vpwr scs8hd_decap_4
XFILLER_9_115 vpwr vgnd scs8hd_fill_2
XFILLER_9_126 vpwr vgnd scs8hd_fill_2
XFILLER_9_148 vgnd vpwr scs8hd_decap_6
XFILLER_13_188 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _115_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_114 vgnd vpwr scs8hd_decap_3
XFILLER_10_147 vgnd vpwr scs8hd_decap_6
XFILLER_10_158 vpwr vgnd scs8hd_fill_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_33_217 vgnd vpwr scs8hd_decap_12
XFILLER_33_206 vpwr vgnd scs8hd_fill_2
XANTENNA__108__B _097_/X vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _103_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_206 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_261 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_200_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_131_ _101_/X _128_/X _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_42 vpwr vgnd scs8hd_fill_2
XFILLER_23_53 vgnd vpwr scs8hd_decap_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_9 vpwr vgnd scs8hd_fill_2
XFILLER_9_33 vpwr vgnd scs8hd_fill_2
XFILLER_9_11 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_21_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_64 vgnd vpwr scs8hd_decap_3
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_114_ _103_/X _115_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__121__B _126_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vgnd vpwr scs8hd_decap_4
XFILLER_29_85 vgnd vpwr scs8hd_decap_3
XFILLER_28_150 vgnd vpwr scs8hd_decap_3
XANTENNA__116__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA__132__A _103_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_19_150 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vpwr vgnd scs8hd_fill_2
XFILLER_31_97 vgnd vpwr scs8hd_decap_3
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_0_252 vpwr vgnd scs8hd_fill_2
XFILLER_0_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__127__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_142 vpwr vgnd scs8hd_fill_2
XFILLER_16_186 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_112 vgnd vpwr scs8hd_decap_4
XFILLER_22_134 vpwr vgnd scs8hd_fill_2
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
XFILLER_26_97 vgnd vpwr scs8hd_fill_1
XFILLER_13_167 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_13_178 vpwr vgnd scs8hd_fill_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
XFILLER_27_248 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_77 vgnd vpwr scs8hd_decap_4
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XFILLER_18_248 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_229 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XANTENNA__140__A _103_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_270 vgnd vpwr scs8hd_decap_6
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_273 vgnd vpwr scs8hd_decap_4
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
X_130_ _099_/X _128_/X _130_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__119__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_4
XANTENNA__135__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_265 vgnd vpwr scs8hd_decap_8
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_76 vgnd vpwr scs8hd_decap_8
XFILLER_18_87 vpwr vgnd scs8hd_fill_2
X_113_ _101_/X _115_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_7 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_5_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_162 vpwr vgnd scs8hd_fill_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_88 vgnd vpwr scs8hd_fill_1
XFILLER_29_53 vgnd vpwr scs8hd_decap_4
XFILLER_28_184 vpwr vgnd scs8hd_fill_2
XFILLER_28_173 vgnd vpwr scs8hd_decap_4
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XANTENNA__132__B _128_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_140 vgnd vpwr scs8hd_fill_1
XFILLER_19_173 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_176 vgnd vpwr scs8hd_decap_4
XFILLER_25_132 vgnd vpwr scs8hd_decap_4
XFILLER_15_66 vpwr vgnd scs8hd_fill_2
XFILLER_40_179 vgnd vpwr scs8hd_decap_12
XFILLER_40_168 vpwr vgnd scs8hd_fill_2
XFILLER_31_10 vgnd vpwr scs8hd_decap_12
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XFILLER_31_157 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__127__B _163_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_235 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _144_/Y mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_4
XFILLER_26_65 vpwr vgnd scs8hd_fill_2
XFILLER_13_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_219 vpwr vgnd scs8hd_fill_2
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_23_99 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XANTENNA__119__C address[5] vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
X_189_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__135__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _144_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_18_22 vgnd vpwr scs8hd_decap_6
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
X_112_ _099_/X _115_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_266 vgnd vpwr scs8hd_decap_8
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_108 vgnd vpwr scs8hd_decap_4
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_141 vpwr vgnd scs8hd_fill_2
XFILLER_34_133 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_199 vpwr vgnd scs8hd_fill_2
XFILLER_25_155 vpwr vgnd scs8hd_fill_2
XFILLER_25_111 vpwr vgnd scs8hd_fill_2
XFILLER_15_23 vpwr vgnd scs8hd_fill_2
XFILLER_31_22 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _176_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_136 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vgnd vpwr scs8hd_decap_3
XFILLER_31_103 vgnd vpwr scs8hd_decap_3
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C address[5] vgnd vpwr scs8hd_diode_2
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_199 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_191 vgnd vpwr scs8hd_decap_4
XFILLER_22_169 vpwr vgnd scs8hd_fill_2
XFILLER_26_22 vpwr vgnd scs8hd_fill_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__138__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _101_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_239 vgnd vpwr scs8hd_decap_4
XFILLER_27_228 vpwr vgnd scs8hd_fill_2
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _157_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__119__D _119_/D vgnd vpwr scs8hd_diode_2
XANTENNA__135__C address[5] vgnd vpwr scs8hd_diode_2
X_188_ _188_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_12 vgnd vpwr scs8hd_fill_1
XFILLER_18_45 vgnd vpwr scs8hd_fill_1
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_234 vpwr vgnd scs8hd_fill_2
XFILLER_11_245 vgnd vpwr scs8hd_decap_8
X_111_ _076_/A _115_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _144_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_7 vgnd vpwr scs8hd_decap_3
XFILLER_34_189 vpwr vgnd scs8hd_fill_2
XFILLER_34_112 vgnd vpwr scs8hd_decap_8
XFILLER_34_101 vpwr vgnd scs8hd_fill_2
XANTENNA__157__A _126_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vgnd vpwr scs8hd_fill_1
XANTENNA__067__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_67 vpwr vgnd scs8hd_fill_2
XFILLER_31_34 vgnd vpwr scs8hd_decap_12
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_167 vpwr vgnd scs8hd_fill_2
XFILLER_31_126 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _119_/D vgnd vpwr scs8hd_diode_2
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_204 vgnd vpwr scs8hd_decap_12
XFILLER_22_104 vgnd vpwr scs8hd_decap_6
XFILLER_30_170 vgnd vpwr scs8hd_decap_6
XFILLER_7_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XFILLER_13_148 vpwr vgnd scs8hd_fill_2
XFILLER_21_192 vpwr vgnd scs8hd_fill_2
XFILLER_36_229 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B _151_/X vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_207 vpwr vgnd scs8hd_fill_2
XFILLER_12_36 vgnd vpwr scs8hd_fill_1
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__080__A _093_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XANTENNA__149__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_221 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _074_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vgnd vpwr scs8hd_fill_1
XFILLER_0_17 vpwr vgnd scs8hd_fill_2
XFILLER_9_37 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_243 vgnd vpwr scs8hd_fill_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__135__D _119_/D vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_202 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _109_/X _115_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _160_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_37_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_47 vgnd vpwr scs8hd_decap_12
XFILLER_28_154 vgnd vpwr scs8hd_decap_6
XFILLER_28_110 vgnd vpwr scs8hd_decap_8
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_154 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _151_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_198 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_168 vpwr vgnd scs8hd_fill_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XANTENNA__067__B _065_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_46 vgnd vpwr scs8hd_decap_12
XFILLER_0_256 vgnd vpwr scs8hd_decap_4
XFILLER_0_267 vgnd vpwr scs8hd_decap_8
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_146 vpwr vgnd scs8hd_fill_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_216 vgnd vpwr scs8hd_decap_12
XFILLER_39_249 vpwr vgnd scs8hd_fill_2
XANTENNA__168__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_116 vgnd vpwr scs8hd_fill_1
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
XFILLER_7_92 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_260 vgnd vpwr scs8hd_decap_12
XFILLER_26_46 vpwr vgnd scs8hd_fill_2
XANTENNA__078__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_160 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__170__B _171_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_59 vgnd vpwr scs8hd_decap_3
XANTENNA__080__B _099_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _090_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_1_.latch data_in _145_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__C address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_23_25 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_29 vpwr vgnd scs8hd_fill_2
X_186_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_236 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_58 vgnd vpwr scs8hd_decap_4
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_203 vgnd vpwr scs8hd_decap_3
XFILLER_11_258 vpwr vgnd scs8hd_fill_2
XANTENNA__162__C _160_/C vgnd vpwr scs8hd_diode_2
X_169_ _083_/X _171_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_188 vgnd vpwr scs8hd_decap_4
XFILLER_28_177 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_17 vgnd vpwr scs8hd_decap_12
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_177 vgnd vpwr scs8hd_decap_4
XFILLER_19_188 vgnd vpwr scs8hd_fill_1
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XANTENNA__067__C _159_/C vgnd vpwr scs8hd_diode_2
XFILLER_33_180 vgnd vpwr scs8hd_fill_1
XFILLER_31_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_191 vpwr vgnd scs8hd_fill_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_239 vgnd vpwr scs8hd_decap_4
XFILLER_39_228 vgnd vpwr scs8hd_decap_4
XANTENNA__168__B _171_/B vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_128 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_272 vgnd vpwr scs8hd_decap_3
XANTENNA__078__B _065_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_69 vpwr vgnd scs8hd_fill_2
XFILLER_26_36 vgnd vpwr scs8hd_fill_1
XANTENNA__094__A address[4] vgnd vpwr scs8hd_diode_2
Xmem_top_track_14.LATCH_0_.latch data_in _148_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XFILLER_8_143 vgnd vpwr scs8hd_decap_8
XFILLER_8_110 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _143_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A _088_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__C _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vgnd vpwr scs8hd_decap_3
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
X_185_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_215 vpwr vgnd scs8hd_fill_2
XFILLER_20_248 vpwr vgnd scs8hd_fill_2
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_48 vgnd vpwr scs8hd_fill_1
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XFILLER_11_226 vpwr vgnd scs8hd_fill_2
X_168_ _099_/A _171_/B _168_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
XFILLER_10_270 vgnd vpwr scs8hd_decap_4
X_099_ _099_/A _099_/X vgnd vpwr scs8hd_buf_1
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XANTENNA__187__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_47 vgnd vpwr scs8hd_fill_1
XFILLER_28_145 vgnd vpwr scs8hd_decap_3
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_29 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_148 vpwr vgnd scs8hd_fill_2
XFILLER_19_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_115 vgnd vpwr scs8hd_decap_4
XFILLER_16_104 vpwr vgnd scs8hd_fill_2
XFILLER_24_170 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_81 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_26 vgnd vpwr scs8hd_decap_4
XANTENNA__078__C _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_35_243 vgnd vpwr scs8hd_fill_1
XANTENNA__195__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_12_39 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_221 vpwr vgnd scs8hd_fill_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_27_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_254 vpwr vgnd scs8hd_fill_2
XFILLER_17_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_202 vpwr vgnd scs8hd_fill_2
XFILLER_23_257 vpwr vgnd scs8hd_fill_2
XFILLER_23_38 vpwr vgnd scs8hd_fill_2
XFILLER_23_49 vpwr vgnd scs8hd_fill_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA__091__C _160_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_9_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
XFILLER_14_235 vgnd vpwr scs8hd_decap_8
X_184_ _184_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _179_/HI mem_top_track_0.LATCH_5_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_238 vgnd vpwr scs8hd_decap_6
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_167_ _068_/X _171_/B _167_/Y vgnd vpwr scs8hd_nor2_4
X_098_ _076_/A _097_/X _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_179 vgnd vpwr scs8hd_decap_4
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_105 vgnd vpwr scs8hd_decap_4
XANTENNA__198__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_119 vgnd vpwr scs8hd_decap_3
XFILLER_31_108 vgnd vpwr scs8hd_decap_3
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_7 vgnd vpwr scs8hd_decap_4
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_62 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_152 vpwr vgnd scs8hd_fill_2
XFILLER_29_241 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _174_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_12_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_17_200 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_266 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _192_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vpwr vgnd scs8hd_fill_2
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XFILLER_9_19 vgnd vpwr scs8hd_decap_3
XFILLER_14_247 vpwr vgnd scs8hd_fill_2
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_50 vgnd vpwr scs8hd_decap_3
XFILLER_13_83 vpwr vgnd scs8hd_fill_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_28 vgnd vpwr scs8hd_fill_1
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _175_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_71 vgnd vpwr scs8hd_decap_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ _165_/X _171_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_097_ _097_/A _097_/X vgnd vpwr scs8hd_buf_1
XFILLER_37_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_51 vgnd vpwr scs8hd_decap_4
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
XFILLER_19_169 vpwr vgnd scs8hd_fill_2
X_149_ _149_/A address[6] address[5] _158_/A vgnd vpwr scs8hd_or3_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_172 vpwr vgnd scs8hd_fill_2
XFILLER_33_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_50 vgnd vpwr scs8hd_fill_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_38_231 vgnd vpwr scs8hd_fill_1
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_142 vgnd vpwr scs8hd_fill_1
XFILLER_21_164 vpwr vgnd scs8hd_fill_2
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XFILLER_8_102 vgnd vpwr scs8hd_decap_8
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XFILLER_35_201 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_259 vpwr vgnd scs8hd_fill_2
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _099_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
X_165_ address[4] address[3] _074_/B _165_/X vgnd vpwr scs8hd_or3_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _074_/B _162_/A _097_/A vgnd vpwr scs8hd_or2_4
XFILLER_1_10 vgnd vpwr scs8hd_decap_12
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _156_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_19 vpwr vgnd scs8hd_fill_2
XFILLER_29_39 vgnd vpwr scs8hd_decap_8
XFILLER_28_137 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_50 vgnd vpwr scs8hd_decap_4
XFILLER_19_83 vgnd vpwr scs8hd_decap_3
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_129 vpwr vgnd scs8hd_fill_2
XFILLER_27_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ _148_/A _148_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_079_ _078_/X _099_/A vgnd vpwr scs8hd_buf_1
XFILLER_15_19 vpwr vgnd scs8hd_fill_2
XFILLER_18_181 vgnd vpwr scs8hd_fill_1
XFILLER_33_195 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_187 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vpwr vgnd scs8hd_fill_2
XFILLER_30_121 vpwr vgnd scs8hd_fill_2
XFILLER_30_110 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_1_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_140 vpwr vgnd scs8hd_fill_2
XFILLER_15_151 vpwr vgnd scs8hd_fill_2
XFILLER_15_173 vpwr vgnd scs8hd_fill_2
XFILLER_15_184 vgnd vpwr scs8hd_decap_3
XFILLER_7_42 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_18 vpwr vgnd scs8hd_fill_2
XFILLER_21_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _144_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_114 vgnd vpwr scs8hd_decap_3
XFILLER_12_165 vgnd vpwr scs8hd_decap_12
XFILLER_16_73 vpwr vgnd scs8hd_fill_2
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _170_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XFILLER_35_213 vgnd vpwr scs8hd_decap_12
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_246 vgnd vpwr scs8hd_decap_8
XFILLER_26_235 vgnd vpwr scs8hd_decap_8
XFILLER_26_224 vgnd vpwr scs8hd_decap_8
XFILLER_26_257 vgnd vpwr scs8hd_decap_12
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_83 vgnd vpwr scs8hd_fill_1
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XANTENNA__100__B _097_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_219 vpwr vgnd scs8hd_fill_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_51 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_164_ _163_/A _163_/B _160_/B _160_/C _164_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
X_095_ _163_/A address[3] _162_/A vgnd vpwr scs8hd_or2_4
XFILLER_27_7 vgnd vpwr scs8hd_decap_3
XFILLER_1_22 vgnd vpwr scs8hd_decap_12
XANTENNA__111__A _076_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_147_ _147_/A _147_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_078_ address[1] _065_/Y _160_/C _078_/X vgnd vpwr scs8hd_or3_4
XANTENNA__106__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
XFILLER_33_141 vgnd vpwr scs8hd_decap_6
XFILLER_25_119 vgnd vpwr scs8hd_fill_1
XFILLER_18_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_16_108 vgnd vpwr scs8hd_decap_6
XFILLER_24_174 vgnd vpwr scs8hd_decap_4
XFILLER_24_141 vpwr vgnd scs8hd_fill_2
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_85 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_98 vgnd vpwr scs8hd_fill_1
XFILLER_38_211 vgnd vpwr scs8hd_decap_3
XFILLER_21_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_188 vpwr vgnd scs8hd_fill_2
XFILLER_12_177 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_269 vgnd vpwr scs8hd_decap_6
XANTENNA__204__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _103_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_4
XFILLER_14_228 vgnd vpwr scs8hd_decap_4
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
XANTENNA__109__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_163_ _163_/A _163_/B _160_/B _159_/C _163_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_10_242 vgnd vpwr scs8hd_fill_1
X_094_ address[4] _163_/A vgnd vpwr scs8hd_inv_8
XANTENNA__111__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_106 vpwr vgnd scs8hd_fill_2
XFILLER_10_10 vpwr vgnd scs8hd_fill_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_6
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XFILLER_10_76 vgnd vpwr scs8hd_decap_8
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_146_ _146_/A _146_/Y vgnd vpwr scs8hd_inv_8
X_077_ address[0] _160_/C vgnd vpwr scs8hd_buf_1
XANTENNA__106__B _097_/X vgnd vpwr scs8hd_diode_2
XANTENNA__122__A _099_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__207__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_24_131 vgnd vpwr scs8hd_fill_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_31 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_145 vgnd vpwr scs8hd_decap_3
XFILLER_7_77 vgnd vpwr scs8hd_fill_1
XFILLER_7_66 vgnd vpwr scs8hd_fill_1
XFILLER_7_11 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A enable vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
X_129_ _076_/A _128_/X _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XFILLER_21_156 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
XFILLER_29_212 vgnd vpwr scs8hd_decap_3
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_112 vgnd vpwr scs8hd_decap_3
XFILLER_12_134 vpwr vgnd scs8hd_fill_2
XFILLER_12_145 vpwr vgnd scs8hd_fill_2
XFILLER_12_189 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_17_215 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XANTENNA__114__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XFILLER_31_262 vgnd vpwr scs8hd_decap_12
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_14.LATCH_1_.latch data_in _147_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__109__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vgnd vpwr scs8hd_decap_12
X_162_ _162_/A _160_/B _160_/C _162_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
X_093_ _093_/A _093_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_254 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_46 vgnd vpwr scs8hd_decap_12
XFILLER_36_140 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_173 vpwr vgnd scs8hd_fill_2
XFILLER_10_55 vgnd vpwr scs8hd_fill_1
XFILLER_10_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_42 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_173 vgnd vpwr scs8hd_decap_4
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_19_97 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/A _145_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_076_ _076_/A _093_/A _076_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__B _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_176 vgnd vpwr scs8hd_decap_4
XFILLER_33_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_173 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_187 vpwr vgnd scs8hd_fill_2
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_45 vgnd vpwr scs8hd_decap_12
XFILLER_7_34 vgnd vpwr scs8hd_decap_8
X_128_ _127_/X _128_/X vgnd vpwr scs8hd_buf_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_3
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_2_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__130__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_31_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_13_55 vpwr vgnd scs8hd_fill_2
XFILLER_13_66 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_223 vgnd vpwr scs8hd_decap_12
XFILLER_9_245 vpwr vgnd scs8hd_fill_2
XFILLER_13_263 vgnd vpwr scs8hd_decap_12
XANTENNA__109__C _074_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _156_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_161_ _162_/A _160_/B _159_/C _161_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_24_54 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_6
XFILLER_24_10 vgnd vpwr scs8hd_decap_4
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_200 vgnd vpwr scs8hd_decap_3
X_092_ _092_/A _093_/B vgnd vpwr scs8hd_buf_1
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_58 vgnd vpwr scs8hd_decap_3
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _135_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_19_54 vgnd vpwr scs8hd_fill_1
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _144_/A _144_/Y vgnd vpwr scs8hd_inv_8
X_075_ _074_/X _093_/A vgnd vpwr scs8hd_buf_1
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_33_199 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_11 vgnd vpwr scs8hd_decap_3
XFILLER_21_77 vpwr vgnd scs8hd_fill_2
XFILLER_30_158 vgnd vpwr scs8hd_fill_1
XFILLER_30_125 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vgnd vpwr scs8hd_decap_4
XFILLER_15_155 vpwr vgnd scs8hd_fill_2
XFILLER_15_177 vgnd vpwr scs8hd_decap_4
XANTENNA__133__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_57 vgnd vpwr scs8hd_decap_4
X_127_ address[4] _163_/B address[5] _119_/D _127_/X vgnd vpwr scs8hd_or4_4
XFILLER_38_236 vgnd vpwr scs8hd_decap_12
XFILLER_16_3 vgnd vpwr scs8hd_decap_4
XFILLER_21_114 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_16_22 vpwr vgnd scs8hd_fill_2
XFILLER_16_88 vpwr vgnd scs8hd_fill_2
XFILLER_32_98 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_239 vgnd vpwr scs8hd_decap_4
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_decap_3
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _147_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_87 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _101_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_272 vgnd vpwr scs8hd_decap_3
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_13_34 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_9_202 vgnd vpwr scs8hd_fill_1
XFILLER_9_235 vgnd vpwr scs8hd_decap_8
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_13_275 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_160_ _160_/A _160_/B _160_/C _160_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_24_88 vgnd vpwr scs8hd_decap_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_091_ address[1] address[2] _160_/C _092_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _068_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_35_10 vgnd vpwr scs8hd_decap_12
X_143_ _143_/A _143_/Y vgnd vpwr scs8hd_inv_8
X_074_ _160_/A _074_/B _074_/X vgnd vpwr scs8hd_or2_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_3
XFILLER_33_101 vpwr vgnd scs8hd_fill_2
XFILLER_18_197 vgnd vpwr scs8hd_decap_6
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_126_ _126_/A _126_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_69 vgnd vpwr scs8hd_decap_8
XFILLER_38_248 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_21_104 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_119 vgnd vpwr scs8hd_decap_12
XFILLER_12_104 vgnd vpwr scs8hd_decap_8
XFILLER_12_126 vpwr vgnd scs8hd_fill_2
XFILLER_16_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_170 vgnd vpwr scs8hd_decap_4
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
X_109_ _163_/A _163_/B _074_/B _109_/X vgnd vpwr scs8hd_or3_4
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vgnd vpwr scs8hd_decap_6
XFILLER_27_33 vgnd vpwr scs8hd_decap_4
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_31_243 vgnd vpwr scs8hd_fill_1
XFILLER_31_221 vpwr vgnd scs8hd_fill_2
XFILLER_31_210 vgnd vpwr scs8hd_decap_8
XANTENNA__155__A _103_/X vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_46 vpwr vgnd scs8hd_fill_2
XFILLER_13_79 vpwr vgnd scs8hd_fill_2
XFILLER_22_232 vgnd vpwr scs8hd_decap_6
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_232 vpwr vgnd scs8hd_fill_2
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_39_162 vpwr vgnd scs8hd_fill_2
XFILLER_39_151 vgnd vpwr scs8hd_fill_1
XFILLER_24_67 vpwr vgnd scs8hd_fill_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_8
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_10_246 vgnd vpwr scs8hd_decap_8
X_090_ _093_/A _171_/A _090_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__152__B _151_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_47 vpwr vgnd scs8hd_fill_2
XFILLER_10_69 vgnd vpwr scs8hd_decap_4
XFILLER_35_22 vgnd vpwr scs8hd_decap_12
XFILLER_27_154 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vgnd vpwr scs8hd_decap_3
XFILLER_27_110 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_23 vgnd vpwr scs8hd_decap_4
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_27_187 vgnd vpwr scs8hd_decap_3
X_142_ _126_/A _142_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_073_ enable _073_/B address[5] _074_/B vgnd vpwr scs8hd_nand3_4
XFILLER_18_8 vpwr vgnd scs8hd_fill_2
XFILLER_18_132 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__A enable vgnd vpwr scs8hd_diode_2
XFILLER_21_46 vgnd vpwr scs8hd_decap_4
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_168 vgnd vpwr scs8hd_decap_3
X_125_ _156_/A _126_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _155_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_149 vgnd vpwr scs8hd_decap_4
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
X_108_ _126_/A _097_/X _108_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__B _160_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_12 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_211 vgnd vpwr scs8hd_decap_3
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _151_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_252 vgnd vpwr scs8hd_decap_8
XANTENNA__171__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_266 vgnd vpwr scs8hd_decap_8
XANTENNA__081__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_6
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_211 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__076__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_177 vgnd vpwr scs8hd_decap_4
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_19_79 vpwr vgnd scs8hd_fill_2
X_210_ _210_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_141_ _156_/A _142_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_072_ address[6] _073_/B vgnd vpwr scs8hd_inv_8
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _145_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_147 vgnd vpwr scs8hd_fill_1
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_191 vgnd vpwr scs8hd_decap_8
XFILLER_24_158 vgnd vpwr scs8hd_fill_1
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
X_124_ _103_/X _126_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_217 vgnd vpwr scs8hd_decap_3
XFILLER_16_69 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _093_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_161 vgnd vpwr scs8hd_decap_4
XFILLER_20_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
X_107_ _093_/B _126_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_121 vgnd vpwr scs8hd_fill_1
XANTENNA__160__C _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XFILLER_26_209 vgnd vpwr scs8hd_decap_3
XANTENNA__169__A _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_81 vgnd vpwr scs8hd_decap_8
XFILLER_8_70 vgnd vpwr scs8hd_decap_8
XANTENNA__079__A _078_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_16_264 vgnd vpwr scs8hd_decap_8
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _146_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _171_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_201 vpwr vgnd scs8hd_fill_2
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_205 vgnd vpwr scs8hd_decap_12
XFILLER_9_249 vgnd vpwr scs8hd_decap_6
XFILLER_13_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_47 vgnd vpwr scs8hd_decap_4
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_226 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__076__B _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_46 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _093_/A vgnd vpwr scs8hd_diode_2
X_140_ _103_/X _142_/B _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ address[4] _163_/B _160_/A vgnd vpwr scs8hd_or2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XFILLER_33_137 vpwr vgnd scs8hd_fill_2
XFILLER_25_90 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _160_/B vgnd vpwr scs8hd_diode_2
XANTENNA__073__C address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_129 vgnd vpwr scs8hd_decap_3
XFILLER_15_115 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_123_ _101_/X _126_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_8 vpwr vgnd scs8hd_fill_2
XFILLER_14_170 vpwr vgnd scs8hd_fill_2
XFILLER_14_192 vgnd vpwr scs8hd_decap_3
XFILLER_21_118 vgnd vpwr scs8hd_fill_1
XANTENNA__190__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_229 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_26 vgnd vpwr scs8hd_decap_3
XFILLER_16_48 vgnd vpwr scs8hd_decap_8
XFILLER_20_140 vgnd vpwr scs8hd_decap_3
XANTENNA__084__B _083_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_184 vpwr vgnd scs8hd_fill_2
XFILLER_11_195 vpwr vgnd scs8hd_fill_2
X_106_ _156_/A _097_/X _106_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__B _171_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_265 vpwr vgnd scs8hd_fill_2
XFILLER_25_254 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_10_238 vgnd vpwr scs8hd_decap_4
XFILLER_6_6 vgnd vpwr scs8hd_decap_8
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_35_58 vgnd vpwr scs8hd_decap_3
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__087__B _170_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_070_ address[3] _163_/B vgnd vpwr scs8hd_inv_8
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_102 vgnd vpwr scs8hd_decap_12
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _148_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__163__D _159_/C vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_199_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_16 vpwr vgnd scs8hd_fill_2
XFILLER_21_27 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_18 vgnd vpwr scs8hd_decap_6
X_122_ _099_/X _126_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_29 vgnd vpwr scs8hd_decap_3
XFILLER_38_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_108 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_7_101 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_105_ _171_/A _156_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_200 vgnd vpwr scs8hd_decap_12
XFILLER_19_230 vpwr vgnd scs8hd_fill_2
XFILLER_19_241 vgnd vpwr scs8hd_decap_3
XFILLER_19_263 vpwr vgnd scs8hd_fill_2
XFILLER_40_203 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B address[3] vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_258 vpwr vgnd scs8hd_fill_2
XFILLER_31_225 vgnd vpwr scs8hd_decap_12
XFILLER_17_81 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__196__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_13_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_236 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_10_206 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_158 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_169 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_198_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_24_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__B _097_/X vgnd vpwr scs8hd_diode_2
X_121_ _076_/A _126_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_83 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__199__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_37_242 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_2.LATCH_0_.latch data_in _144_/A _160_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_7_113 vgnd vpwr scs8hd_decap_8
XFILLER_11_153 vgnd vpwr scs8hd_fill_1
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _103_/X _097_/X _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_71 vgnd vpwr scs8hd_decap_4
XFILLER_34_212 vpwr vgnd scs8hd_fill_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_234 vgnd vpwr scs8hd_decap_4
XFILLER_25_212 vpwr vgnd scs8hd_fill_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_237 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _175_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_215 vpwr vgnd scs8hd_fill_2
XFILLER_30_270 vgnd vpwr scs8hd_decap_4
XFILLER_13_29 vgnd vpwr scs8hd_decap_3
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_219 vpwr vgnd scs8hd_fill_2
XFILLER_13_215 vpwr vgnd scs8hd_fill_2
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _144_/A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_5_30 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_6
XFILLER_30_60 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_3_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_27_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
X_120_ _119_/X _126_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_51 vgnd vpwr scs8hd_decap_4
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _145_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _147_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_18 vpwr vgnd scs8hd_fill_2
XFILLER_20_110 vpwr vgnd scs8hd_fill_2
XFILLER_20_165 vgnd vpwr scs8hd_fill_1
XFILLER_20_198 vgnd vpwr scs8hd_decap_4
XFILLER_28_210 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
X_103_ _170_/A _103_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_11_176 vpwr vgnd scs8hd_fill_2
XFILLER_14_7 vpwr vgnd scs8hd_fill_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_3
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XFILLER_16_235 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_205 vpwr vgnd scs8hd_fill_2
XFILLER_22_249 vgnd vpwr scs8hd_decap_8
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_249 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _146_/A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_271 vgnd vpwr scs8hd_decap_4
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_42 vgnd vpwr scs8hd_decap_12
XFILLER_39_179 vgnd vpwr scs8hd_decap_4
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_62 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _197_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _083_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_193 vpwr vgnd scs8hd_fill_2
XFILLER_4_6 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_116 vgnd vpwr scs8hd_decap_3
XFILLER_18_149 vgnd vpwr scs8hd_decap_4
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_196_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_119 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_163 vgnd vpwr scs8hd_decap_3
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_152 vgnd vpwr scs8hd_fill_1
XFILLER_14_174 vgnd vpwr scs8hd_decap_4
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XFILLER_11_166 vpwr vgnd scs8hd_fill_2
XFILLER_11_199 vpwr vgnd scs8hd_fill_2
X_102_ _101_/X _097_/X _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_8_64 vgnd vpwr scs8hd_decap_3
XFILLER_27_29 vpwr vgnd scs8hd_fill_2
XFILLER_27_18 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_25_258 vgnd vpwr scs8hd_decap_4
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_16_203 vgnd vpwr scs8hd_fill_1
XFILLER_17_73 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _103_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_250 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_228 vpwr vgnd scs8hd_fill_2
XFILLER_28_61 vgnd vpwr scs8hd_fill_1
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _154_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_54 vgnd vpwr scs8hd_decap_6
XFILLER_39_158 vpwr vgnd scs8hd_fill_2
XFILLER_39_147 vgnd vpwr scs8hd_decap_4
XFILLER_40_18 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_52 vgnd vpwr scs8hd_fill_1
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XFILLER_29_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_106 vpwr vgnd scs8hd_fill_2
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XFILLER_35_172 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_128 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_161 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_40 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_172 vgnd vpwr scs8hd_decap_4
XFILLER_32_175 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _172_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_175 vgnd vpwr scs8hd_decap_3
XFILLER_23_153 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_97 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _093_/B vgnd vpwr scs8hd_diode_2
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_37_234 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_123 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_101_ _083_/X _101_/X vgnd vpwr scs8hd_buf_1
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XFILLER_11_112 vgnd vpwr scs8hd_decap_4
XFILLER_11_156 vgnd vpwr scs8hd_fill_1
XFILLER_19_234 vgnd vpwr scs8hd_decap_4
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_19_267 vgnd vpwr scs8hd_decap_8
XFILLER_8_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__210__A _210_/A vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XFILLER_17_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _097_/X vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _119_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_15_270 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_262 vpwr vgnd scs8hd_fill_2
XFILLER_21_273 vgnd vpwr scs8hd_decap_4
XANTENNA__205__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_40 vgnd vpwr scs8hd_decap_4
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _183_/HI _145_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_50 vgnd vpwr scs8hd_decap_8
XFILLER_36_129 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _146_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XFILLER_26_184 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XANTENNA__112__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_165 vpwr vgnd scs8hd_fill_2
XFILLER_32_132 vpwr vgnd scs8hd_fill_2
XFILLER_17_140 vpwr vgnd scs8hd_fill_2
XFILLER_23_198 vpwr vgnd scs8hd_fill_2
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_11_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_187 vgnd vpwr scs8hd_decap_3
X_177_ _177_/HI _177_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__123__A _101_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_102 vgnd vpwr scs8hd_decap_6
XFILLER_20_157 vpwr vgnd scs8hd_fill_2
XFILLER_28_235 vgnd vpwr scs8hd_decap_12
XFILLER_28_224 vgnd vpwr scs8hd_decap_8
XANTENNA__208__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_100_ _099_/X _097_/X _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_202 vgnd vpwr scs8hd_fill_1
XFILLER_19_213 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _149_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _148_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_11_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XFILLER_22_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_74 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_241 vgnd vpwr scs8hd_decap_12
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _101_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_87 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_top_track_16.LATCH_5_.latch/Q
+ mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _126_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_31 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_86 vpwr vgnd scs8hd_fill_2
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_1_262 vgnd vpwr scs8hd_decap_12
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_188 vgnd vpwr scs8hd_fill_1
XFILLER_11_77 vgnd vpwr scs8hd_decap_4
XFILLER_14_133 vpwr vgnd scs8hd_fill_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
XFILLER_14_166 vpwr vgnd scs8hd_fill_2
X_176_ _176_/HI _176_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_247 vgnd vpwr scs8hd_decap_12
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
X_159_ _160_/A _160_/B _159_/C _159_/Y vgnd vpwr scs8hd_nor3_4
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__134__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _174_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_6
XFILLER_16_228 vgnd vpwr scs8hd_decap_4
XFILLER_16_239 vgnd vpwr scs8hd_decap_4
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA__129__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_209 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_28_64 vgnd vpwr scs8hd_fill_1
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XFILLER_12_253 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _128_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_22 vgnd vpwr scs8hd_decap_4
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_29_172 vpwr vgnd scs8hd_fill_2
XFILLER_29_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _148_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__B _126_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_197 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_164 vgnd vpwr scs8hd_decap_3
XFILLER_26_120 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_1_274 vgnd vpwr scs8hd_decap_3
XFILLER_17_153 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vpwr vgnd scs8hd_fill_2
XFILLER_32_145 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_112 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _178_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_175_ _175_/HI _175_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_55 vgnd vpwr scs8hd_fill_1
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_46 vgnd vpwr scs8hd_decap_8
XFILLER_8_35 vpwr vgnd scs8hd_fill_2
XFILLER_8_13 vgnd vpwr scs8hd_fill_1
X_158_ _158_/A _160_/B vgnd vpwr scs8hd_buf_1
X_089_ _088_/X _171_/A vgnd vpwr scs8hd_buf_1
XANTENNA__134__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XFILLER_10_192 vgnd vpwr scs8hd_decap_8
XANTENNA__150__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_25_229 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_22 vgnd vpwr scs8hd_decap_4
XFILLER_17_33 vpwr vgnd scs8hd_fill_2
XFILLER_17_77 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_fill_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_30_254 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_4
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_210 vgnd vpwr scs8hd_decap_4
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _143_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_14 vpwr vgnd scs8hd_fill_2
XFILLER_10_6 vpwr vgnd scs8hd_fill_2
Xmem_top_track_2.LATCH_1_.latch data_in _143_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_77 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _177_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_176 vgnd vpwr scs8hd_fill_1
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_176 vgnd vpwr scs8hd_decap_8
XFILLER_26_132 vgnd vpwr scs8hd_decap_4
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_253 vpwr vgnd scs8hd_fill_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_113 vgnd vpwr scs8hd_decap_4
XFILLER_32_102 vgnd vpwr scs8hd_fill_1
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_17_176 vgnd vpwr scs8hd_fill_1
XANTENNA__137__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_13 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_102 vpwr vgnd scs8hd_fill_2
X_174_ _174_/HI _174_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_7 vgnd vpwr scs8hd_decap_3
XANTENNA__148__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_127 vpwr vgnd scs8hd_fill_2
XFILLER_20_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_109 vpwr vgnd scs8hd_fill_2
XFILLER_11_149 vgnd vpwr scs8hd_decap_4
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XFILLER_22_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_205 vgnd vpwr scs8hd_fill_1
XFILLER_19_238 vgnd vpwr scs8hd_fill_1
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_19_249 vgnd vpwr scs8hd_decap_4
X_157_ _126_/A _151_/X _157_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
XFILLER_10_182 vgnd vpwr scs8hd_decap_4
XFILLER_40_6 vgnd vpwr scs8hd_decap_12
XANTENNA__150__B address[3] vgnd vpwr scs8hd_diode_2
X_088_ address[1] address[2] _159_/C _088_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_4
XFILLER_33_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_230 vgnd vpwr scs8hd_decap_8
XFILLER_17_56 vgnd vpwr scs8hd_decap_3
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _182_/HI _144_/Y mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_30_222 vpwr vgnd scs8hd_fill_2
X_209_ _209_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__161__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _145_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_222 vpwr vgnd scs8hd_fill_2
XFILLER_21_233 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__071__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA__066__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_fill_1
XFILLER_14_46 vgnd vpwr scs8hd_decap_6
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vpwr vgnd scs8hd_fill_2
XFILLER_30_89 vgnd vpwr scs8hd_decap_3
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_155 vpwr vgnd scs8hd_fill_2
XFILLER_35_144 vgnd vpwr scs8hd_decap_6
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_188 vgnd vpwr scs8hd_decap_6
X_190_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_100 vgnd vpwr scs8hd_decap_4
XFILLER_40_191 vgnd vpwr scs8hd_decap_12
XFILLER_32_169 vgnd vpwr scs8hd_decap_6
XANTENNA__153__B _151_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _147_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_36 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_114 vpwr vgnd scs8hd_fill_2
X_173_ _173_/HI _173_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_217 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__164__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_140 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XFILLER_28_206 vpwr vgnd scs8hd_fill_2
XANTENNA__074__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_156_ _156_/A _151_/X _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_10_172 vgnd vpwr scs8hd_fill_1
X_087_ _093_/A _170_/A _087_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__C _158_/A vgnd vpwr scs8hd_diode_2
XANTENNA__159__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _068_/X vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _146_/Y mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_208_ chanx_right_in[4] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__161__B _160_/B vgnd vpwr scs8hd_diode_2
X_139_ _101_/X _142_/B _139_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_9_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _173_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_245 vpwr vgnd scs8hd_fill_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA__071__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_78 vgnd vpwr scs8hd_decap_12
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__156__B _151_/X vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _093_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_29_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_6
XANTENNA__167__A _068_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_8
XFILLER_26_101 vpwr vgnd scs8hd_fill_2
XFILLER_25_24 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[0] vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _153_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_159 vpwr vgnd scs8hd_fill_2
XFILLER_11_26 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_137 vpwr vgnd scs8hd_fill_2
XFILLER_14_148 vpwr vgnd scs8hd_fill_2
X_172_ _093_/B _171_/B _172_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_229 vgnd vpwr scs8hd_decap_3
XANTENNA__164__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_130 vgnd vpwr scs8hd_decap_4
XFILLER_13_192 vgnd vpwr scs8hd_decap_3
XFILLER_9_196 vgnd vpwr scs8hd_decap_6
XFILLER_36_273 vpwr vgnd scs8hd_fill_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__074__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_47 vgnd vpwr scs8hd_decap_8
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_8_16 vgnd vpwr scs8hd_decap_4
X_086_ _086_/A _170_/A vgnd vpwr scs8hd_buf_1
X_155_ _103_/X _151_/X _155_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_162 vpwr vgnd scs8hd_fill_2
XFILLER_33_210 vgnd vpwr scs8hd_decap_4
XANTENNA__159__B _160_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_273 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _171_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_207_ chanx_right_in[5] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
XANTENNA__161__C _159_/C vgnd vpwr scs8hd_diode_2
X_138_ _099_/X _142_/B _138_/Y vgnd vpwr scs8hd_nor2_4
X_069_ _068_/X _076_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_28_13 vgnd vpwr scs8hd_decap_12
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_57 vgnd vpwr scs8hd_decap_4
XFILLER_28_46 vpwr vgnd scs8hd_fill_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _171_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_187 vgnd vpwr scs8hd_decap_12
XFILLER_38_176 vgnd vpwr scs8hd_decap_8
XFILLER_38_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_14_26 vgnd vpwr scs8hd_fill_1
XANTENNA__082__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_176 vgnd vpwr scs8hd_decap_4
XFILLER_29_165 vpwr vgnd scs8hd_fill_2
XFILLER_20_80 vgnd vpwr scs8hd_fill_1
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XANTENNA__167__B _171_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _210_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_157 vgnd vpwr scs8hd_decap_4
XFILLER_26_124 vpwr vgnd scs8hd_fill_2
XFILLER_25_36 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_8
XFILLER_32_149 vgnd vpwr scs8hd_decap_4
XFILLER_32_105 vgnd vpwr scs8hd_fill_1
XFILLER_17_157 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_116 vgnd vpwr scs8hd_decap_4
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XFILLER_23_149 vpwr vgnd scs8hd_fill_2
XFILLER_39_260 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
X_171_ _171_/A _171_/B _171_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_182 vgnd vpwr scs8hd_decap_6
XANTENNA__164__C _160_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_15_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_241 vgnd vpwr scs8hd_decap_12
XFILLER_11_108 vpwr vgnd scs8hd_fill_2
XANTENNA__090__B _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_252 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_39 vpwr vgnd scs8hd_fill_2
X_154_ _101_/X _151_/X _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
X_085_ _082_/A address[2] _160_/C _086_/A vgnd vpwr scs8hd_or3_4
XFILLER_26_7 vgnd vpwr scs8hd_decap_8
XANTENNA__159__C _159_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__191__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_26 vgnd vpwr scs8hd_fill_1
XFILLER_17_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_15_266 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_30_258 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_137_ _076_/A _142_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_068_ _067_/X _068_/X vgnd vpwr scs8hd_buf_1
XFILLER_17_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__186__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XFILLER_21_258 vpwr vgnd scs8hd_fill_2
XFILLER_21_269 vpwr vgnd scs8hd_fill_2
XFILLER_9_82 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _184_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_36 vgnd vpwr scs8hd_fill_1
XFILLER_28_25 vgnd vpwr scs8hd_decap_6
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_18 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XANTENNA__082__C _159_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_144 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _148_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _188_/A vgnd vpwr scs8hd_inv_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _093_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_40_172 vgnd vpwr scs8hd_decap_4
XFILLER_32_128 vpwr vgnd scs8hd_fill_2
XFILLER_25_180 vgnd vpwr scs8hd_fill_1
XFILLER_15_81 vpwr vgnd scs8hd_fill_2
XFILLER_31_91 vgnd vpwr scs8hd_decap_4
XFILLER_31_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_161 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B address[2] vgnd vpwr scs8hd_diode_2
X_170_ _170_/A _171_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_106 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__164__D _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_154 vgnd vpwr scs8hd_fill_1
XFILLER_36_253 vgnd vpwr scs8hd_decap_12
XANTENNA__189__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_275 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _144_/A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_153_ _099_/X _151_/X _153_/Y vgnd vpwr scs8hd_nor2_4
X_084_ _093_/A _083_/X _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_231 vgnd vpwr scs8hd_decap_4
XFILLER_19_7 vgnd vpwr scs8hd_fill_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _177_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__085__C _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_226 vgnd vpwr scs8hd_decap_12
XFILLER_30_204 vpwr vgnd scs8hd_fill_2
XFILLER_15_223 vpwr vgnd scs8hd_fill_2
X_205_ chanx_left_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_81 vgnd vpwr scs8hd_decap_3
X_136_ _135_/X _142_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_6 vpwr vgnd scs8hd_fill_2
X_067_ address[1] _065_/Y _159_/C _067_/X vgnd vpwr scs8hd_or3_4
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_50 vgnd vpwr scs8hd_decap_4
XFILLER_21_226 vpwr vgnd scs8hd_fill_2
XFILLER_21_237 vgnd vpwr scs8hd_decap_3
XANTENNA__096__B _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_259 vgnd vpwr scs8hd_decap_12
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ address[4] address[3] address[5] _119_/D _119_/X vgnd vpwr scs8hd_or4_4
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_14 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_35_159 vpwr vgnd scs8hd_fill_2
XFILLER_29_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_258 vpwr vgnd scs8hd_fill_2
XFILLER_17_104 vgnd vpwr scs8hd_fill_1
XFILLER_40_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_60 vgnd vpwr scs8hd_fill_1
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_118 vgnd vpwr scs8hd_fill_1
XANTENNA__088__C _159_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _176_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _144_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_100 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_111 vpwr vgnd scs8hd_fill_2
XFILLER_9_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_36_265 vgnd vpwr scs8hd_decap_8
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_243 vgnd vpwr scs8hd_fill_1
X_083_ _083_/A _083_/X vgnd vpwr scs8hd_buf_1
X_152_ _068_/X _151_/X _152_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_143 vpwr vgnd scs8hd_fill_2
XFILLER_10_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_210 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_202 vgnd vpwr scs8hd_decap_6
X_204_ chanx_left_in[4] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_30_238 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_066_ address[0] _159_/C vgnd vpwr scs8hd_inv_8
XFILLER_23_71 vgnd vpwr scs8hd_decap_4
X_135_ _163_/A address[3] address[5] _119_/D _135_/X vgnd vpwr scs8hd_or4_4
XFILLER_23_60 vgnd vpwr scs8hd_fill_1
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_95 vpwr vgnd scs8hd_fill_2
XFILLER_21_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
X_118_ _149_/A _073_/B _119_/D vgnd vpwr scs8hd_or2_4
XFILLER_14_18 vpwr vgnd scs8hd_fill_2
XFILLER_14_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_26 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_7_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_72 vgnd vpwr scs8hd_decap_8
XFILLER_29_81 vpwr vgnd scs8hd_fill_2
XFILLER_26_105 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_34_193 vgnd vpwr scs8hd_decap_4
XFILLER_34_160 vgnd vpwr scs8hd_fill_1
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_7 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_71 vgnd vpwr scs8hd_decap_6
XFILLER_15_94 vpwr vgnd scs8hd_fill_2
XFILLER_31_130 vgnd vpwr scs8hd_decap_4
XFILLER_16_171 vpwr vgnd scs8hd_fill_2
XFILLER_16_182 vpwr vgnd scs8hd_fill_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vgnd vpwr scs8hd_fill_1
XFILLER_13_163 vpwr vgnd scs8hd_fill_2
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
XFILLER_27_211 vpwr vgnd scs8hd_fill_2
X_151_ _151_/A _151_/X vgnd vpwr scs8hd_buf_1
X_082_ _082_/A address[2] _159_/C _083_/A vgnd vpwr scs8hd_or3_4
XFILLER_10_166 vgnd vpwr scs8hd_decap_6
XFILLER_10_188 vpwr vgnd scs8hd_fill_2
XFILLER_12_51 vgnd vpwr scs8hd_decap_8
XFILLER_12_73 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
XFILLER_18_244 vpwr vgnd scs8hd_fill_2
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_29 vpwr vgnd scs8hd_fill_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_247 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _173_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_203_ _203_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _143_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_15_258 vpwr vgnd scs8hd_fill_2
X_065_ address[2] _065_/Y vgnd vpwr scs8hd_inv_8
X_134_ _126_/A _128_/X _134_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_10 vgnd vpwr scs8hd_decap_4
XFILLER_0_21 vgnd vpwr scs8hd_decap_8
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XFILLER_12_228 vgnd vpwr scs8hd_decap_4
XFILLER_34_93 vgnd vpwr scs8hd_decap_8
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
X_117_ enable _149_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_4
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_38 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_37_191 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_20_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_180 vgnd vpwr scs8hd_fill_1
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_128 vpwr vgnd scs8hd_fill_2
XFILLER_25_29 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_109 vpwr vgnd scs8hd_fill_2
XFILLER_25_172 vpwr vgnd scs8hd_fill_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _101_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_150 vgnd vpwr scs8hd_decap_3
XFILLER_31_197 vpwr vgnd scs8hd_fill_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_31_153 vpwr vgnd scs8hd_fill_2
XFILLER_39_264 vgnd vpwr scs8hd_decap_12
XFILLER_39_253 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_50 vpwr vgnd scs8hd_fill_2
XFILLER_9_157 vgnd vpwr scs8hd_decap_12
XFILLER_13_197 vgnd vpwr scs8hd_decap_3
XFILLER_9_179 vgnd vpwr scs8hd_decap_4
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_43 vgnd vpwr scs8hd_decap_12
XFILLER_36_223 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
X_150_ address[4] address[3] _158_/A _151_/A vgnd vpwr scs8hd_or3_4
X_081_ address[1] _082_/A vgnd vpwr scs8hd_inv_8
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_226 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vpwr vgnd scs8hd_fill_2
XANTENNA__200__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
X_202_ _202_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_30_218 vpwr vgnd scs8hd_fill_2
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
X_133_ _156_/A _128_/X _133_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _147_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _109_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_75 vgnd vpwr scs8hd_decap_4
XFILLER_9_86 vgnd vpwr scs8hd_decap_3
XFILLER_20_273 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vgnd vpwr scs8hd_fill_1
XFILLER_11_262 vpwr vgnd scs8hd_fill_2
X_116_ _126_/A _115_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _171_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_159 vgnd vpwr scs8hd_decap_8
XFILLER_28_192 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_34_140 vgnd vpwr scs8hd_decap_8
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in _146_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_107 vpwr vgnd scs8hd_fill_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_8
XFILLER_25_195 vpwr vgnd scs8hd_fill_2
XFILLER_25_184 vpwr vgnd scs8hd_fill_2
XFILLER_25_151 vpwr vgnd scs8hd_fill_2
XFILLER_31_84 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B _097_/X vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XFILLER_22_165 vpwr vgnd scs8hd_fill_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_6
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_169 vgnd vpwr scs8hd_decap_4
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_13_143 vgnd vpwr scs8hd_decap_3
XANTENNA__113__A _101_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_55 vgnd vpwr scs8hd_decap_6
XFILLER_27_235 vpwr vgnd scs8hd_fill_2
XFILLER_27_224 vpwr vgnd scs8hd_fill_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ _093_/A _099_/A _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_10_102 vgnd vpwr scs8hd_decap_12
XFILLER_10_124 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_208 vgnd vpwr scs8hd_decap_6
XFILLER_15_227 vgnd vpwr scs8hd_decap_4
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _152_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_132_ _103_/X _128_/X _132_/Y vgnd vpwr scs8hd_nor2_4
X_201_ _201_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _193_/A vgnd vpwr scs8hd_inv_1
XFILLER_9_54 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_230 vgnd vpwr scs8hd_decap_6
XFILLER_20_252 vgnd vpwr scs8hd_decap_4
XFILLER_18_41 vgnd vpwr scs8hd_decap_4
XFILLER_11_230 vpwr vgnd scs8hd_fill_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_11_274 vgnd vpwr scs8hd_decap_3
X_115_ _156_/A _115_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__121__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _143_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vgnd vpwr scs8hd_decap_4
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_53 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

