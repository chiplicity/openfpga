magic
tech EFS8A
magscale 1 2
timestamp 1602269293
<< locali >>
rect 9631 23137 9758 23171
rect 15335 23137 15462 23171
rect 24627 23137 24662 23171
rect 24627 22049 24662 22083
rect 7935 21097 7941 21131
rect 7935 21029 7969 21097
rect 1547 20213 1685 20247
rect 10787 20009 10793 20043
rect 10787 19941 10821 20009
rect 24627 19873 24662 19907
rect 12081 19295 12115 19397
rect 11655 18785 11690 18819
rect 3151 18071 3185 18139
rect 3151 18037 3157 18071
rect 10051 17833 10057 17867
rect 10051 17765 10085 17833
rect 24501 17119 24535 17153
rect 24501 17085 24615 17119
rect 5457 15487 5491 15657
rect 6929 15453 7055 15487
rect 7021 15351 7055 15453
rect 7205 14331 7239 14569
rect 6043 13345 6078 13379
rect 8861 13175 8895 13481
rect 1547 13141 1593 13175
rect 11891 10217 11897 10251
rect 11891 10149 11925 10217
rect 15663 8041 15669 8075
rect 15663 7973 15697 8041
rect 25455 6817 25490 6851
rect 15663 5865 15669 5899
rect 15663 5797 15697 5865
rect 15243 4641 15370 4675
rect 12771 2601 12909 2635
<< viali >>
rect 10977 24361 11011 24395
rect 1476 24225 1510 24259
rect 8652 24225 8686 24259
rect 10793 24225 10827 24259
rect 16472 24225 16506 24259
rect 24660 24225 24694 24259
rect 1547 24021 1581 24055
rect 8401 24021 8435 24055
rect 8723 24021 8757 24055
rect 10057 24021 10091 24055
rect 16543 24021 16577 24055
rect 24731 24021 24765 24055
rect 2237 23817 2271 23851
rect 4261 23817 4295 23851
rect 9413 23817 9447 23851
rect 10977 23817 11011 23851
rect 14473 23817 14507 23851
rect 15945 23817 15979 23851
rect 20453 23817 20487 23851
rect 25145 23817 25179 23851
rect 16497 23749 16531 23783
rect 25513 23749 25547 23783
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 3776 23613 3810 23647
rect 4629 23613 4663 23647
rect 5365 23613 5399 23647
rect 8309 23613 8343 23647
rect 8769 23613 8803 23647
rect 9873 23613 9907 23647
rect 9965 23613 9999 23647
rect 10517 23613 10551 23647
rect 14289 23613 14323 23647
rect 15444 23613 15478 23647
rect 16732 23613 16766 23647
rect 17233 23613 17267 23647
rect 19952 23613 19986 23647
rect 24660 23613 24694 23647
rect 1547 23545 1581 23579
rect 4721 23545 4755 23579
rect 15531 23545 15565 23579
rect 16819 23545 16853 23579
rect 20039 23545 20073 23579
rect 3847 23477 3881 23511
rect 8125 23477 8159 23511
rect 8585 23477 8619 23511
rect 10057 23477 10091 23511
rect 14933 23477 14967 23511
rect 24731 23477 24765 23511
rect 9827 23273 9861 23307
rect 16313 23273 16347 23307
rect 13737 23205 13771 23239
rect 1444 23137 1478 23171
rect 2824 23137 2858 23171
rect 5365 23137 5399 23171
rect 8217 23137 8251 23171
rect 9597 23137 9631 23171
rect 11345 23137 11379 23171
rect 15301 23137 15335 23171
rect 24593 23137 24627 23171
rect 13645 23069 13679 23103
rect 14565 23069 14599 23103
rect 14197 23001 14231 23035
rect 1547 22933 1581 22967
rect 2053 22933 2087 22967
rect 2927 22933 2961 22967
rect 4629 22933 4663 22967
rect 5181 22933 5215 22967
rect 8309 22933 8343 22967
rect 11529 22933 11563 22967
rect 15531 22933 15565 22967
rect 15853 22933 15887 22967
rect 24731 22933 24765 22967
rect 1593 22729 1627 22763
rect 2973 22729 3007 22763
rect 8217 22729 8251 22763
rect 11345 22729 11379 22763
rect 15485 22729 15519 22763
rect 18705 22729 18739 22763
rect 24685 22729 24719 22763
rect 3663 22661 3697 22695
rect 4629 22593 4663 22627
rect 9781 22593 9815 22627
rect 13461 22593 13495 22627
rect 13737 22593 13771 22627
rect 14381 22593 14415 22627
rect 15945 22593 15979 22627
rect 16221 22593 16255 22627
rect 2329 22525 2363 22559
rect 3560 22525 3594 22559
rect 3985 22525 4019 22559
rect 10425 22525 10459 22559
rect 13369 22525 13403 22559
rect 18220 22525 18254 22559
rect 4445 22457 4479 22491
rect 4721 22457 4755 22491
rect 5273 22457 5307 22491
rect 8861 22457 8895 22491
rect 8953 22457 8987 22491
rect 9505 22457 9539 22491
rect 10333 22457 10367 22491
rect 14473 22457 14507 22491
rect 15025 22457 15059 22491
rect 16037 22457 16071 22491
rect 2237 22389 2271 22423
rect 5549 22389 5583 22423
rect 7757 22389 7791 22423
rect 8677 22389 8711 22423
rect 10149 22389 10183 22423
rect 14105 22389 14139 22423
rect 18291 22389 18325 22423
rect 5181 22185 5215 22219
rect 9045 22185 9079 22219
rect 12817 22185 12851 22219
rect 13553 22185 13587 22219
rect 14105 22185 14139 22219
rect 2145 22117 2179 22151
rect 5457 22117 5491 22151
rect 6009 22117 6043 22151
rect 8217 22117 8251 22151
rect 9781 22117 9815 22151
rect 9873 22117 9907 22151
rect 11621 22117 11655 22151
rect 15393 22117 15427 22151
rect 15485 22117 15519 22151
rect 16037 22117 16071 22151
rect 6996 22049 7030 22083
rect 14289 22049 14323 22083
rect 24593 22049 24627 22083
rect 2053 21981 2087 22015
rect 4261 21981 4295 22015
rect 5365 21981 5399 22015
rect 8125 21981 8159 22015
rect 10057 21981 10091 22015
rect 11529 21981 11563 22015
rect 2605 21913 2639 21947
rect 7849 21913 7883 21947
rect 8677 21913 8711 21947
rect 12081 21913 12115 21947
rect 7067 21845 7101 21879
rect 10885 21845 10919 21879
rect 24731 21845 24765 21879
rect 2053 21641 2087 21675
rect 3525 21641 3559 21675
rect 3893 21641 3927 21675
rect 6101 21641 6135 21675
rect 7021 21641 7055 21675
rect 7941 21641 7975 21675
rect 10333 21641 10367 21675
rect 11805 21641 11839 21675
rect 13737 21641 13771 21675
rect 14473 21641 14507 21675
rect 15945 21641 15979 21675
rect 16635 21641 16669 21675
rect 24685 21641 24719 21675
rect 2789 21573 2823 21607
rect 7573 21573 7607 21607
rect 8677 21573 8711 21607
rect 2237 21505 2271 21539
rect 3157 21505 3191 21539
rect 5181 21505 5215 21539
rect 5549 21505 5583 21539
rect 8125 21505 8159 21539
rect 9919 21505 9953 21539
rect 10885 21505 10919 21539
rect 3709 21437 3743 21471
rect 4261 21437 4295 21471
rect 6837 21437 6871 21471
rect 9827 21437 9861 21471
rect 12449 21437 12483 21471
rect 12909 21437 12943 21471
rect 16532 21437 16566 21471
rect 1685 21369 1719 21403
rect 2329 21369 2363 21403
rect 4997 21369 5031 21403
rect 5273 21369 5307 21403
rect 8217 21369 8251 21403
rect 9045 21369 9079 21403
rect 10701 21369 10735 21403
rect 10977 21369 11011 21403
rect 11529 21369 11563 21403
rect 15025 21369 15059 21403
rect 15117 21369 15151 21403
rect 15669 21369 15703 21403
rect 16957 21369 16991 21403
rect 6653 21301 6687 21335
rect 9597 21301 9631 21335
rect 12173 21301 12207 21335
rect 12541 21301 12575 21335
rect 14749 21301 14783 21335
rect 5825 21097 5859 21131
rect 7205 21097 7239 21131
rect 7941 21097 7975 21131
rect 8493 21097 8527 21131
rect 8769 21097 8803 21131
rect 9873 21097 9907 21131
rect 11437 21097 11471 21131
rect 11805 21097 11839 21131
rect 13921 21097 13955 21131
rect 2053 21029 2087 21063
rect 5267 21029 5301 21063
rect 10879 21029 10913 21063
rect 13363 21029 13397 21063
rect 15485 21029 15519 21063
rect 16865 21029 16899 21063
rect 2973 20961 3007 20995
rect 10517 20961 10551 20995
rect 16957 20961 16991 20995
rect 1961 20893 1995 20927
rect 2605 20893 2639 20927
rect 4905 20893 4939 20927
rect 7573 20893 7607 20927
rect 13001 20893 13035 20927
rect 15393 20893 15427 20927
rect 15669 20893 15703 20927
rect 1685 20757 1719 20791
rect 6193 20757 6227 20791
rect 6929 20757 6963 20791
rect 12449 20757 12483 20791
rect 14933 20757 14967 20791
rect 3341 20553 3375 20587
rect 5825 20553 5859 20587
rect 9505 20553 9539 20587
rect 10241 20553 10275 20587
rect 14473 20553 14507 20587
rect 17233 20553 17267 20587
rect 4077 20485 4111 20519
rect 7941 20485 7975 20519
rect 8493 20485 8527 20519
rect 2421 20417 2455 20451
rect 8585 20417 8619 20451
rect 15761 20417 15795 20451
rect 16313 20417 16347 20451
rect 1476 20349 1510 20383
rect 1961 20349 1995 20383
rect 4905 20349 4939 20383
rect 6653 20349 6687 20383
rect 7113 20349 7147 20383
rect 7389 20349 7423 20383
rect 9873 20349 9907 20383
rect 10793 20349 10827 20383
rect 13553 20349 13587 20383
rect 2329 20281 2363 20315
rect 2783 20281 2817 20315
rect 4445 20281 4479 20315
rect 4721 20281 4755 20315
rect 5267 20281 5301 20315
rect 6193 20281 6227 20315
rect 8906 20281 8940 20315
rect 10609 20281 10643 20315
rect 13874 20281 13908 20315
rect 15025 20281 15059 20315
rect 16129 20281 16163 20315
rect 16405 20281 16439 20315
rect 16957 20281 16991 20315
rect 1685 20213 1719 20247
rect 6929 20213 6963 20247
rect 10977 20213 11011 20247
rect 12449 20213 12483 20247
rect 13093 20213 13127 20247
rect 13461 20213 13495 20247
rect 15301 20213 15335 20247
rect 6561 20009 6595 20043
rect 7573 20009 7607 20043
rect 8125 20009 8159 20043
rect 10241 20009 10275 20043
rect 10793 20009 10827 20043
rect 11345 20009 11379 20043
rect 13185 20009 13219 20043
rect 14197 20009 14231 20043
rect 2421 19941 2455 19975
rect 4997 19941 5031 19975
rect 5089 19941 5123 19975
rect 12357 19941 12391 19975
rect 15622 19941 15656 19975
rect 17233 19941 17267 19975
rect 18613 19941 18647 19975
rect 6469 19873 6503 19907
rect 7021 19873 7055 19907
rect 8033 19873 8067 19907
rect 8585 19873 8619 19907
rect 10425 19873 10459 19907
rect 18705 19873 18739 19907
rect 24593 19873 24627 19907
rect 2329 19805 2363 19839
rect 2605 19805 2639 19839
rect 7941 19805 7975 19839
rect 12265 19805 12299 19839
rect 12541 19805 12575 19839
rect 15301 19805 15335 19839
rect 17141 19805 17175 19839
rect 17601 19805 17635 19839
rect 5549 19737 5583 19771
rect 1869 19669 1903 19703
rect 3341 19669 3375 19703
rect 4445 19669 4479 19703
rect 13553 19669 13587 19703
rect 14013 19669 14047 19703
rect 16221 19669 16255 19703
rect 24731 19669 24765 19703
rect 1593 19465 1627 19499
rect 2421 19465 2455 19499
rect 5365 19465 5399 19499
rect 6469 19465 6503 19499
rect 8217 19465 8251 19499
rect 10517 19465 10551 19499
rect 11805 19465 11839 19499
rect 14933 19465 14967 19499
rect 17141 19465 17175 19499
rect 18705 19465 18739 19499
rect 24685 19465 24719 19499
rect 5733 19397 5767 19431
rect 6193 19397 6227 19431
rect 12081 19397 12115 19431
rect 12173 19397 12207 19431
rect 3801 19329 3835 19363
rect 4721 19329 4755 19363
rect 10793 19329 10827 19363
rect 11437 19329 11471 19363
rect 14013 19329 14047 19363
rect 1409 19261 1443 19295
rect 2605 19261 2639 19295
rect 6929 19261 6963 19295
rect 8401 19261 8435 19295
rect 8861 19261 8895 19295
rect 9413 19261 9447 19295
rect 12081 19261 12115 19295
rect 12449 19261 12483 19295
rect 12909 19261 12943 19295
rect 15761 19261 15795 19295
rect 16313 19261 16347 19295
rect 2145 19193 2179 19227
rect 2967 19193 3001 19227
rect 4445 19193 4479 19227
rect 4537 19193 4571 19227
rect 6837 19193 6871 19227
rect 10149 19193 10183 19227
rect 10885 19193 10919 19227
rect 13185 19193 13219 19227
rect 14375 19193 14409 19227
rect 15301 19193 15335 19227
rect 15577 19193 15611 19227
rect 3525 19125 3559 19159
rect 4169 19125 4203 19159
rect 7941 19125 7975 19159
rect 8493 19125 8527 19159
rect 13921 19125 13955 19159
rect 15853 19125 15887 19159
rect 17509 19125 17543 19159
rect 4353 18921 4387 18955
rect 8033 18921 8067 18955
rect 11069 18921 11103 18955
rect 12817 18921 12851 18955
rect 15117 18921 15151 18955
rect 2145 18853 2179 18887
rect 3341 18853 3375 18887
rect 6561 18853 6595 18887
rect 7389 18853 7423 18887
rect 13737 18853 13771 18887
rect 15577 18853 15611 18887
rect 16957 18853 16991 18887
rect 4169 18785 4203 18819
rect 7941 18785 7975 18819
rect 8401 18785 8435 18819
rect 10241 18785 10275 18819
rect 11621 18785 11655 18819
rect 13001 18785 13035 18819
rect 13461 18785 13495 18819
rect 2053 18717 2087 18751
rect 2329 18717 2363 18751
rect 5181 18717 5215 18751
rect 6469 18717 6503 18751
rect 7113 18717 7147 18751
rect 15485 18717 15519 18751
rect 16129 18717 16163 18751
rect 1685 18649 1719 18683
rect 11759 18649 11793 18683
rect 2973 18581 3007 18615
rect 6193 18581 6227 18615
rect 10333 18581 10367 18615
rect 12541 18581 12575 18615
rect 14105 18581 14139 18615
rect 16405 18581 16439 18615
rect 2053 18377 2087 18411
rect 7941 18377 7975 18411
rect 11713 18377 11747 18411
rect 1639 18309 1673 18343
rect 7481 18309 7515 18343
rect 12173 18309 12207 18343
rect 15025 18309 15059 18343
rect 5273 18241 5307 18275
rect 6285 18241 6319 18275
rect 6929 18241 6963 18275
rect 10149 18241 10183 18275
rect 13277 18241 13311 18275
rect 14105 18241 14139 18275
rect 15393 18241 15427 18275
rect 15945 18241 15979 18275
rect 16221 18241 16255 18275
rect 1568 18173 1602 18207
rect 2789 18173 2823 18207
rect 9045 18173 9079 18207
rect 9413 18173 9447 18207
rect 12541 18173 12575 18207
rect 13001 18173 13035 18207
rect 5365 18105 5399 18139
rect 5917 18105 5951 18139
rect 7021 18105 7055 18139
rect 8401 18105 8435 18139
rect 10241 18105 10275 18139
rect 10793 18105 10827 18139
rect 14426 18105 14460 18139
rect 16037 18105 16071 18139
rect 2697 18037 2731 18071
rect 3157 18037 3191 18071
rect 3709 18037 3743 18071
rect 4077 18037 4111 18071
rect 5089 18037 5123 18071
rect 6653 18037 6687 18071
rect 9965 18037 9999 18071
rect 11069 18037 11103 18071
rect 13553 18037 13587 18071
rect 14013 18037 14047 18071
rect 15761 18037 15795 18071
rect 16865 18037 16899 18071
rect 1409 17833 1443 17867
rect 6469 17833 6503 17867
rect 7573 17833 7607 17867
rect 8033 17833 8067 17867
rect 8401 17833 8435 17867
rect 10057 17833 10091 17867
rect 10609 17833 10643 17867
rect 13369 17833 13403 17867
rect 15117 17833 15151 17867
rect 15761 17833 15795 17867
rect 2605 17765 2639 17799
rect 5267 17765 5301 17799
rect 7015 17765 7049 17799
rect 10885 17765 10919 17799
rect 12265 17765 12299 17799
rect 12909 17765 12943 17799
rect 11529 17697 11563 17731
rect 13093 17697 13127 17731
rect 13553 17697 13587 17731
rect 15945 17697 15979 17731
rect 16865 17697 16899 17731
rect 17325 17697 17359 17731
rect 2329 17629 2363 17663
rect 2513 17629 2547 17663
rect 4905 17629 4939 17663
rect 6653 17629 6687 17663
rect 9689 17629 9723 17663
rect 11897 17629 11931 17663
rect 17417 17629 17451 17663
rect 3065 17561 3099 17595
rect 5825 17561 5859 17595
rect 1869 17493 1903 17527
rect 4353 17493 4387 17527
rect 8861 17493 8895 17527
rect 11345 17493 11379 17527
rect 11667 17493 11701 17527
rect 11805 17493 11839 17527
rect 12541 17493 12575 17527
rect 14105 17493 14139 17527
rect 8861 17289 8895 17323
rect 10149 17289 10183 17323
rect 13093 17289 13127 17323
rect 14657 17289 14691 17323
rect 16589 17289 16623 17323
rect 17233 17289 17267 17323
rect 5733 17221 5767 17255
rect 6653 17221 6687 17255
rect 8539 17221 8573 17255
rect 8677 17221 8711 17255
rect 11897 17221 11931 17255
rect 24777 17221 24811 17255
rect 1869 17153 1903 17187
rect 2697 17153 2731 17187
rect 4169 17153 4203 17187
rect 7205 17153 7239 17187
rect 7941 17153 7975 17187
rect 8769 17153 8803 17187
rect 9781 17153 9815 17187
rect 10425 17153 10459 17187
rect 16221 17153 16255 17187
rect 24501 17153 24535 17187
rect 25145 17153 25179 17187
rect 4537 17085 4571 17119
rect 5089 17085 5123 17119
rect 5273 17085 5307 17119
rect 8309 17085 8343 17119
rect 13461 17085 13495 17119
rect 14381 17085 14415 17119
rect 15117 17085 15151 17119
rect 15761 17085 15795 17119
rect 16808 17085 16842 17119
rect 16911 17085 16945 17119
rect 2421 17017 2455 17051
rect 2513 17017 2547 17051
rect 3801 17017 3835 17051
rect 6929 17017 6963 17051
rect 7021 17017 7055 17051
rect 8401 17017 8435 17051
rect 10517 17017 10551 17051
rect 11069 17017 11103 17051
rect 13823 17017 13857 17051
rect 2237 16949 2271 16983
rect 3341 16949 3375 16983
rect 5181 16949 5215 16983
rect 6193 16949 6227 16983
rect 11529 16949 11563 16983
rect 12449 16949 12483 16983
rect 15485 16949 15519 16983
rect 17601 16949 17635 16983
rect 3525 16745 3559 16779
rect 4353 16745 4387 16779
rect 5181 16745 5215 16779
rect 6193 16745 6227 16779
rect 6929 16745 6963 16779
rect 9505 16745 9539 16779
rect 10977 16745 11011 16779
rect 13277 16745 13311 16779
rect 14013 16745 14047 16779
rect 2599 16677 2633 16711
rect 4813 16677 4847 16711
rect 10609 16677 10643 16711
rect 12173 16677 12207 16711
rect 15393 16677 15427 16711
rect 15485 16677 15519 16711
rect 4169 16609 4203 16643
rect 5457 16609 5491 16643
rect 5733 16609 5767 16643
rect 6101 16609 6135 16643
rect 7297 16609 7331 16643
rect 9873 16609 9907 16643
rect 11253 16609 11287 16643
rect 11437 16609 11471 16643
rect 12449 16609 12483 16643
rect 13001 16609 13035 16643
rect 13553 16609 13587 16643
rect 24660 16609 24694 16643
rect 2237 16541 2271 16575
rect 10020 16541 10054 16575
rect 10241 16541 10275 16575
rect 11805 16541 11839 16575
rect 15669 16541 15703 16575
rect 3157 16473 3191 16507
rect 7481 16473 7515 16507
rect 8769 16473 8803 16507
rect 11575 16473 11609 16507
rect 12817 16473 12851 16507
rect 8493 16405 8527 16439
rect 10149 16405 10183 16439
rect 11713 16405 11747 16439
rect 24731 16405 24765 16439
rect 2329 16201 2363 16235
rect 4629 16201 4663 16235
rect 8217 16201 8251 16235
rect 8677 16201 8711 16235
rect 8861 16201 8895 16235
rect 9873 16201 9907 16235
rect 11805 16201 11839 16235
rect 13093 16201 13127 16235
rect 13461 16201 13495 16235
rect 15761 16201 15795 16235
rect 16129 16201 16163 16235
rect 24685 16201 24719 16235
rect 8539 16133 8573 16167
rect 12587 16133 12621 16167
rect 2697 16065 2731 16099
rect 7205 16065 7239 16099
rect 8769 16065 8803 16099
rect 12173 16065 12207 16099
rect 12817 16065 12851 16099
rect 15485 16065 15519 16099
rect 1460 15997 1494 16031
rect 1869 15997 1903 16031
rect 3065 15997 3099 16031
rect 3433 15997 3467 16031
rect 3617 15997 3651 16031
rect 4721 15997 4755 16031
rect 5273 15997 5307 16031
rect 12679 15997 12713 16031
rect 1547 15929 1581 15963
rect 6929 15929 6963 15963
rect 7021 15929 7055 15963
rect 8401 15929 8435 15963
rect 10333 15929 10367 15963
rect 10425 15929 10459 15963
rect 10977 15929 11011 15963
rect 12449 15929 12483 15963
rect 13829 15929 13863 15963
rect 14841 15929 14875 15963
rect 14933 15929 14967 15963
rect 2881 15861 2915 15895
rect 4261 15861 4295 15895
rect 4813 15861 4847 15895
rect 5733 15861 5767 15895
rect 6193 15861 6227 15895
rect 6653 15861 6687 15895
rect 7941 15861 7975 15895
rect 9505 15861 9539 15895
rect 11437 15861 11471 15895
rect 14657 15861 14691 15895
rect 1547 15657 1581 15691
rect 2329 15657 2363 15691
rect 3433 15657 3467 15691
rect 5273 15657 5307 15691
rect 5457 15657 5491 15691
rect 7205 15657 7239 15691
rect 10241 15657 10275 15691
rect 11897 15657 11931 15691
rect 13461 15657 13495 15691
rect 14841 15657 14875 15691
rect 15301 15657 15335 15691
rect 2421 15589 2455 15623
rect 4629 15589 4663 15623
rect 1444 15521 1478 15555
rect 2513 15521 2547 15555
rect 4776 15521 4810 15555
rect 6285 15589 6319 15623
rect 6377 15589 6411 15623
rect 11069 15589 11103 15623
rect 12449 15589 12483 15623
rect 8033 15521 8067 15555
rect 12817 15521 12851 15555
rect 16348 15521 16382 15555
rect 4997 15453 5031 15487
rect 5457 15453 5491 15487
rect 7757 15453 7791 15487
rect 10977 15453 11011 15487
rect 11345 15453 11379 15487
rect 9413 15385 9447 15419
rect 12265 15385 12299 15419
rect 4905 15317 4939 15351
rect 5641 15317 5675 15351
rect 6009 15317 6043 15351
rect 7021 15317 7055 15351
rect 7573 15317 7607 15351
rect 8861 15317 8895 15351
rect 9873 15317 9907 15351
rect 10701 15317 10735 15351
rect 16451 15317 16485 15351
rect 1593 15113 1627 15147
rect 2421 15113 2455 15147
rect 4353 15113 4387 15147
rect 4721 15113 4755 15147
rect 6653 15113 6687 15147
rect 8033 15113 8067 15147
rect 8493 15113 8527 15147
rect 9781 15113 9815 15147
rect 11161 15113 11195 15147
rect 11529 15113 11563 15147
rect 16313 15113 16347 15147
rect 10793 15045 10827 15079
rect 5273 14977 5307 15011
rect 11897 14977 11931 15011
rect 2053 14909 2087 14943
rect 2881 14909 2915 14943
rect 6837 14909 6871 14943
rect 9873 14909 9907 14943
rect 12265 14909 12299 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 2789 14841 2823 14875
rect 3243 14841 3277 14875
rect 5365 14841 5399 14875
rect 5917 14841 5951 14875
rect 6285 14841 6319 14875
rect 7199 14841 7233 14875
rect 8585 14841 8619 14875
rect 10194 14841 10228 14875
rect 3801 14773 3835 14807
rect 5089 14773 5123 14807
rect 7757 14773 7791 14807
rect 12541 14773 12575 14807
rect 4537 14569 4571 14603
rect 7113 14569 7147 14603
rect 7205 14569 7239 14603
rect 9965 14569 9999 14603
rect 12817 14569 12851 14603
rect 16865 14569 16899 14603
rect 2605 14501 2639 14535
rect 6514 14501 6548 14535
rect 4629 14433 4663 14467
rect 5181 14433 5215 14467
rect 5733 14433 5767 14467
rect 2513 14365 2547 14399
rect 3157 14365 3191 14399
rect 5365 14365 5399 14399
rect 6193 14365 6227 14399
rect 7941 14501 7975 14535
rect 10378 14501 10412 14535
rect 11989 14501 12023 14535
rect 8033 14433 8067 14467
rect 16681 14433 16715 14467
rect 10057 14365 10091 14399
rect 11897 14365 11931 14399
rect 12173 14365 12207 14399
rect 6101 14297 6135 14331
rect 7205 14297 7239 14331
rect 7389 14229 7423 14263
rect 8953 14229 8987 14263
rect 10977 14229 11011 14263
rect 11345 14229 11379 14263
rect 1777 14025 1811 14059
rect 6285 14025 6319 14059
rect 6561 14025 6595 14059
rect 7941 14025 7975 14059
rect 9229 14025 9263 14059
rect 11897 14025 11931 14059
rect 16681 14025 16715 14059
rect 7481 13957 7515 13991
rect 11161 13957 11195 13991
rect 2789 13889 2823 13923
rect 3801 13889 3835 13923
rect 5917 13889 5951 13923
rect 9321 13889 9355 13923
rect 9689 13889 9723 13923
rect 10149 13889 10183 13923
rect 10609 13889 10643 13923
rect 12449 13889 12483 13923
rect 3065 13821 3099 13855
rect 3709 13821 3743 13855
rect 4997 13821 5031 13855
rect 5181 13821 5215 13855
rect 5641 13821 5675 13855
rect 9100 13821 9134 13855
rect 4353 13753 4387 13787
rect 6929 13753 6963 13787
rect 7021 13753 7055 13787
rect 8953 13753 8987 13787
rect 10701 13753 10735 13787
rect 11529 13753 11563 13787
rect 1869 13685 1903 13719
rect 2421 13685 2455 13719
rect 2973 13685 3007 13719
rect 4721 13685 4755 13719
rect 8401 13685 8435 13719
rect 8769 13685 8803 13719
rect 2237 13481 2271 13515
rect 3525 13481 3559 13515
rect 5135 13481 5169 13515
rect 6561 13481 6595 13515
rect 8125 13481 8159 13515
rect 8861 13481 8895 13515
rect 9045 13481 9079 13515
rect 11897 13481 11931 13515
rect 2605 13413 2639 13447
rect 3157 13413 3191 13447
rect 1476 13345 1510 13379
rect 5032 13345 5066 13379
rect 6009 13345 6043 13379
rect 6929 13345 6963 13379
rect 7481 13345 7515 13379
rect 2513 13277 2547 13311
rect 7849 13277 7883 13311
rect 6147 13209 6181 13243
rect 7646 13209 7680 13243
rect 11345 13413 11379 13447
rect 10701 13345 10735 13379
rect 12208 13345 12242 13379
rect 1593 13141 1627 13175
rect 5549 13141 5583 13175
rect 7389 13141 7423 13175
rect 7757 13141 7791 13175
rect 8861 13141 8895 13175
rect 10057 13141 10091 13175
rect 12311 13141 12345 13175
rect 1685 12937 1719 12971
rect 2053 12937 2087 12971
rect 4997 12937 5031 12971
rect 6101 12937 6135 12971
rect 7941 12937 7975 12971
rect 10701 12937 10735 12971
rect 11621 12937 11655 12971
rect 12173 12937 12207 12971
rect 7619 12869 7653 12903
rect 7757 12869 7791 12903
rect 8493 12869 8527 12903
rect 2513 12801 2547 12835
rect 2789 12801 2823 12835
rect 7849 12801 7883 12835
rect 10057 12801 10091 12835
rect 2881 12733 2915 12767
rect 6653 12733 6687 12767
rect 9597 12733 9631 12767
rect 9965 12733 9999 12767
rect 11136 12733 11170 12767
rect 12817 12733 12851 12767
rect 13369 12733 13403 12767
rect 7481 12665 7515 12699
rect 8953 12665 8987 12699
rect 13553 12665 13587 12699
rect 7297 12597 7331 12631
rect 9413 12597 9447 12631
rect 11207 12597 11241 12631
rect 12633 12597 12667 12631
rect 2881 12393 2915 12427
rect 7205 12393 7239 12427
rect 9873 12393 9907 12427
rect 10149 12325 10183 12359
rect 1409 12257 1443 12291
rect 7792 12257 7826 12291
rect 10241 12257 10275 12291
rect 11713 12257 11747 12291
rect 13277 12257 13311 12291
rect 13829 12257 13863 12291
rect 12081 12189 12115 12223
rect 12449 12189 12483 12223
rect 12909 12189 12943 12223
rect 14013 12189 14047 12223
rect 7573 12121 7607 12155
rect 1593 12053 1627 12087
rect 7895 12053 7929 12087
rect 8309 12053 8343 12087
rect 11161 12053 11195 12087
rect 11529 12053 11563 12087
rect 11851 12053 11885 12087
rect 11989 12053 12023 12087
rect 14381 12053 14415 12087
rect 15853 12053 15887 12087
rect 2237 11849 2271 11883
rect 7757 11849 7791 11883
rect 9873 11849 9907 11883
rect 10793 11849 10827 11883
rect 12081 11849 12115 11883
rect 13829 11849 13863 11883
rect 24777 11849 24811 11883
rect 1547 11713 1581 11747
rect 10885 11713 10919 11747
rect 15853 11713 15887 11747
rect 16221 11713 16255 11747
rect 1444 11645 1478 11679
rect 1869 11645 1903 11679
rect 9321 11645 9355 11679
rect 10664 11645 10698 11679
rect 11713 11645 11747 11679
rect 12633 11645 12667 11679
rect 14381 11645 14415 11679
rect 14933 11645 14967 11679
rect 24593 11645 24627 11679
rect 25145 11645 25179 11679
rect 8677 11577 8711 11611
rect 10517 11577 10551 11611
rect 13185 11577 13219 11611
rect 15945 11577 15979 11611
rect 8493 11509 8527 11543
rect 10149 11509 10183 11543
rect 11161 11509 11195 11543
rect 13461 11509 13495 11543
rect 15577 11509 15611 11543
rect 10701 11305 10735 11339
rect 12633 11305 12667 11339
rect 14381 11305 14415 11339
rect 16865 11305 16899 11339
rect 13823 11237 13857 11271
rect 15485 11237 15519 11271
rect 9689 11169 9723 11203
rect 10241 11169 10275 11203
rect 11529 11169 11563 11203
rect 13461 11169 13495 11203
rect 10425 11101 10459 11135
rect 11253 11101 11287 11135
rect 15393 11101 15427 11135
rect 15761 11101 15795 11135
rect 11161 10965 11195 10999
rect 12265 10965 12299 10999
rect 16313 10965 16347 10999
rect 10149 10761 10183 10795
rect 11529 10761 11563 10795
rect 11805 10761 11839 10795
rect 12173 10761 12207 10795
rect 13553 10761 13587 10795
rect 14013 10761 14047 10795
rect 15485 10761 15519 10795
rect 15761 10761 15795 10795
rect 16957 10761 16991 10795
rect 24777 10761 24811 10795
rect 16589 10693 16623 10727
rect 10609 10625 10643 10659
rect 12541 10625 12575 10659
rect 12817 10625 12851 10659
rect 14197 10625 14231 10659
rect 16037 10625 16071 10659
rect 24593 10557 24627 10591
rect 10517 10489 10551 10523
rect 10971 10489 11005 10523
rect 12633 10489 12667 10523
rect 14559 10489 14593 10523
rect 16129 10489 16163 10523
rect 9689 10421 9723 10455
rect 15117 10421 15151 10455
rect 25237 10421 25271 10455
rect 10977 10217 11011 10251
rect 11897 10217 11931 10251
rect 12449 10217 12483 10251
rect 12725 10217 12759 10251
rect 14289 10217 14323 10251
rect 24777 10217 24811 10251
rect 13461 10149 13495 10183
rect 14657 10149 14691 10183
rect 15669 10149 15703 10183
rect 16221 10149 16255 10183
rect 10057 10081 10091 10115
rect 10425 10081 10459 10115
rect 17084 10081 17118 10115
rect 24593 10081 24627 10115
rect 10701 10013 10735 10047
rect 11529 10013 11563 10047
rect 13369 10013 13403 10047
rect 13645 10013 13679 10047
rect 15577 10013 15611 10047
rect 17187 9945 17221 9979
rect 9689 9673 9723 9707
rect 11897 9673 11931 9707
rect 12265 9673 12299 9707
rect 13461 9673 13495 9707
rect 15209 9673 15243 9707
rect 15577 9673 15611 9707
rect 17049 9673 17083 9707
rect 24685 9673 24719 9707
rect 25375 9673 25409 9707
rect 1593 9605 1627 9639
rect 11437 9605 11471 9639
rect 13093 9605 13127 9639
rect 13921 9605 13955 9639
rect 12541 9537 12575 9571
rect 1409 9469 1443 9503
rect 15393 9469 15427 9503
rect 16313 9469 16347 9503
rect 23765 9469 23799 9503
rect 25304 9469 25338 9503
rect 25697 9469 25731 9503
rect 10885 9401 10919 9435
rect 10977 9401 11011 9435
rect 12633 9401 12667 9435
rect 2053 9333 2087 9367
rect 10057 9333 10091 9367
rect 10701 9333 10735 9367
rect 23489 9333 23523 9367
rect 24133 9333 24167 9367
rect 10471 9129 10505 9163
rect 10885 9129 10919 9163
rect 12357 9129 12391 9163
rect 15577 9129 15611 9163
rect 11345 9061 11379 9095
rect 24041 9061 24075 9095
rect 24593 9061 24627 9095
rect 7481 8993 7515 9027
rect 7665 8993 7699 9027
rect 10400 8993 10434 9027
rect 8033 8925 8067 8959
rect 11713 8925 11747 8959
rect 22845 8925 22879 8959
rect 23949 8925 23983 8959
rect 8309 8789 8343 8823
rect 11483 8789 11517 8823
rect 11621 8789 11655 8823
rect 11989 8789 12023 8823
rect 12817 8789 12851 8823
rect 14473 8789 14507 8823
rect 24869 8789 24903 8823
rect 1593 8585 1627 8619
rect 10425 8585 10459 8619
rect 11897 8585 11931 8619
rect 14381 8585 14415 8619
rect 23397 8585 23431 8619
rect 23949 8585 23983 8619
rect 8493 8517 8527 8551
rect 24685 8517 24719 8551
rect 8585 8449 8619 8483
rect 11069 8449 11103 8483
rect 13645 8449 13679 8483
rect 14473 8449 14507 8483
rect 24133 8449 24167 8483
rect 1409 8381 1443 8415
rect 8364 8381 8398 8415
rect 12909 8381 12943 8415
rect 13369 8381 13403 8415
rect 15393 8381 15427 8415
rect 8217 8313 8251 8347
rect 14794 8313 14828 8347
rect 24225 8313 24259 8347
rect 25053 8313 25087 8347
rect 2053 8245 2087 8279
rect 7113 8245 7147 8279
rect 7573 8245 7607 8279
rect 8033 8245 8067 8279
rect 8861 8245 8895 8279
rect 10977 8245 11011 8279
rect 11529 8245 11563 8279
rect 12817 8245 12851 8279
rect 7665 8041 7699 8075
rect 8309 8041 8343 8075
rect 11345 8041 11379 8075
rect 12909 8041 12943 8075
rect 15669 8041 15703 8075
rect 24317 7973 24351 8007
rect 24869 7973 24903 8007
rect 7021 7905 7055 7939
rect 11529 7905 11563 7939
rect 11989 7905 12023 7939
rect 13277 7905 13311 7939
rect 13737 7905 13771 7939
rect 23188 7905 23222 7939
rect 7389 7837 7423 7871
rect 12265 7837 12299 7871
rect 14013 7837 14047 7871
rect 15301 7837 15335 7871
rect 24225 7837 24259 7871
rect 7186 7769 7220 7803
rect 7297 7701 7331 7735
rect 8585 7701 8619 7735
rect 10885 7701 10919 7735
rect 14381 7701 14415 7735
rect 16221 7701 16255 7735
rect 23259 7701 23293 7735
rect 1547 7497 1581 7531
rect 6653 7497 6687 7531
rect 7297 7497 7331 7531
rect 10241 7497 10275 7531
rect 10931 7497 10965 7531
rect 13277 7497 13311 7531
rect 14473 7497 14507 7531
rect 15669 7497 15703 7531
rect 23213 7497 23247 7531
rect 10609 7429 10643 7463
rect 11069 7429 11103 7463
rect 15393 7429 15427 7463
rect 24869 7429 24903 7463
rect 6285 7361 6319 7395
rect 11161 7361 11195 7395
rect 11529 7361 11563 7395
rect 24317 7361 24351 7395
rect 25605 7361 25639 7395
rect 1444 7293 1478 7327
rect 1869 7293 1903 7327
rect 3617 7293 3651 7327
rect 4353 7293 4387 7327
rect 7205 7293 7239 7327
rect 7757 7293 7791 7327
rect 8953 7293 8987 7327
rect 9137 7293 9171 7327
rect 13461 7293 13495 7327
rect 14013 7293 14047 7327
rect 4445 7225 4479 7259
rect 8217 7225 8251 7259
rect 9781 7225 9815 7259
rect 10793 7225 10827 7259
rect 12173 7225 12207 7259
rect 14197 7225 14231 7259
rect 24409 7225 24443 7259
rect 7021 7157 7055 7191
rect 11805 7157 11839 7191
rect 12909 7157 12943 7191
rect 24133 7157 24167 7191
rect 25237 7157 25271 7191
rect 15393 6953 15427 6987
rect 24133 6953 24167 6987
rect 7205 6885 7239 6919
rect 7849 6885 7883 6919
rect 13553 6885 13587 6919
rect 1685 6817 1719 6851
rect 1869 6817 1903 6851
rect 6561 6817 6595 6851
rect 8033 6817 8067 6851
rect 8585 6817 8619 6851
rect 11161 6817 11195 6851
rect 15301 6817 15335 6851
rect 15853 6817 15887 6851
rect 24501 6817 24535 6851
rect 25421 6817 25455 6851
rect 2237 6749 2271 6783
rect 8769 6749 8803 6783
rect 9045 6749 9079 6783
rect 11529 6749 11563 6783
rect 13461 6749 13495 6783
rect 14105 6749 14139 6783
rect 11437 6681 11471 6715
rect 25559 6681 25593 6715
rect 7573 6613 7607 6647
rect 10885 6613 10919 6647
rect 11326 6613 11360 6647
rect 11621 6613 11655 6647
rect 24869 6613 24903 6647
rect 8033 6409 8067 6443
rect 9413 6409 9447 6443
rect 10241 6409 10275 6443
rect 11805 6409 11839 6443
rect 14565 6409 14599 6443
rect 15853 6409 15887 6443
rect 16221 6409 16255 6443
rect 23949 6409 23983 6443
rect 6193 6341 6227 6375
rect 9689 6341 9723 6375
rect 13369 6341 13403 6375
rect 13645 6341 13679 6375
rect 14013 6341 14047 6375
rect 25513 6341 25547 6375
rect 3157 6273 3191 6307
rect 8493 6273 8527 6307
rect 12449 6273 12483 6307
rect 14657 6273 14691 6307
rect 24133 6273 24167 6307
rect 25053 6273 25087 6307
rect 1685 6205 1719 6239
rect 1777 6205 1811 6239
rect 1961 6205 1995 6239
rect 2421 6205 2455 6239
rect 2789 6205 2823 6239
rect 6929 6205 6963 6239
rect 7481 6205 7515 6239
rect 10609 6205 10643 6239
rect 10793 6205 10827 6239
rect 11253 6205 11287 6239
rect 15577 6205 15611 6239
rect 7665 6137 7699 6171
rect 8855 6137 8889 6171
rect 11529 6137 11563 6171
rect 12770 6137 12804 6171
rect 14978 6137 15012 6171
rect 23397 6137 23431 6171
rect 24225 6137 24259 6171
rect 24777 6137 24811 6171
rect 6561 6069 6595 6103
rect 12173 6069 12207 6103
rect 18245 6069 18279 6103
rect 1685 5865 1719 5899
rect 2421 5865 2455 5899
rect 6929 5865 6963 5899
rect 10885 5865 10919 5899
rect 11253 5865 11287 5899
rect 11529 5865 11563 5899
rect 12449 5865 12483 5899
rect 14289 5865 14323 5899
rect 14749 5865 14783 5899
rect 15669 5865 15703 5899
rect 8125 5797 8159 5831
rect 8217 5797 8251 5831
rect 9873 5797 9907 5831
rect 13046 5797 13080 5831
rect 18705 5797 18739 5831
rect 1869 5729 1903 5763
rect 12725 5729 12759 5763
rect 15301 5729 15335 5763
rect 23857 5729 23891 5763
rect 9781 5661 9815 5695
rect 10057 5661 10091 5695
rect 18613 5661 18647 5695
rect 8677 5593 8711 5627
rect 19165 5593 19199 5627
rect 9045 5525 9079 5559
rect 13645 5525 13679 5559
rect 16221 5525 16255 5559
rect 24041 5525 24075 5559
rect 2237 5321 2271 5355
rect 7757 5321 7791 5355
rect 9873 5321 9907 5355
rect 14105 5321 14139 5355
rect 15393 5321 15427 5355
rect 16865 5321 16899 5355
rect 17877 5321 17911 5355
rect 23489 5321 23523 5355
rect 24041 5321 24075 5355
rect 8033 5253 8067 5287
rect 12173 5253 12207 5287
rect 13737 5253 13771 5287
rect 19809 5253 19843 5287
rect 8677 5185 8711 5219
rect 10793 5185 10827 5219
rect 12817 5185 12851 5219
rect 13461 5185 13495 5219
rect 14381 5185 14415 5219
rect 15025 5185 15059 5219
rect 16221 5185 16255 5219
rect 18797 5185 18831 5219
rect 19165 5185 19199 5219
rect 24501 5185 24535 5219
rect 1444 5117 1478 5151
rect 1869 5117 1903 5151
rect 8998 5049 9032 5083
rect 10517 5049 10551 5083
rect 10609 5049 10643 5083
rect 11897 5049 11931 5083
rect 12886 5049 12920 5083
rect 14473 5049 14507 5083
rect 15945 5049 15979 5083
rect 16037 5049 16071 5083
rect 18889 5049 18923 5083
rect 24225 5049 24259 5083
rect 24317 5049 24351 5083
rect 1547 4981 1581 5015
rect 8493 4981 8527 5015
rect 9597 4981 9631 5015
rect 10241 4981 10275 5015
rect 11529 4981 11563 5015
rect 15669 4981 15703 5015
rect 18613 4981 18647 5015
rect 8585 4777 8619 4811
rect 10701 4777 10735 4811
rect 12449 4777 12483 4811
rect 18613 4777 18647 4811
rect 22891 4777 22925 4811
rect 24225 4777 24259 4811
rect 24731 4777 24765 4811
rect 9045 4709 9079 4743
rect 9873 4709 9907 4743
rect 10425 4709 10459 4743
rect 12633 4709 12667 4743
rect 14197 4709 14231 4743
rect 15853 4709 15887 4743
rect 12725 4641 12759 4675
rect 15209 4641 15243 4675
rect 18245 4641 18279 4675
rect 19165 4641 19199 4675
rect 22820 4641 22854 4675
rect 24660 4641 24694 4675
rect 9781 4573 9815 4607
rect 15439 4437 15473 4471
rect 1547 4233 1581 4267
rect 10057 4233 10091 4267
rect 10425 4233 10459 4267
rect 12725 4233 12759 4267
rect 13645 4233 13679 4267
rect 15393 4233 15427 4267
rect 18245 4233 18279 4267
rect 19257 4233 19291 4267
rect 24685 4233 24719 4267
rect 14565 4097 14599 4131
rect 22845 4097 22879 4131
rect 1444 4029 1478 4063
rect 1869 4029 1903 4063
rect 8953 4029 8987 4063
rect 9137 4029 9171 4063
rect 13921 4029 13955 4063
rect 18864 4029 18898 4063
rect 9781 3961 9815 3995
rect 18935 3893 18969 3927
rect 8493 3553 8527 3587
rect 9740 3553 9774 3587
rect 16221 3553 16255 3587
rect 19165 3553 19199 3587
rect 9827 3485 9861 3519
rect 8677 3349 8711 3383
rect 16405 3349 16439 3383
rect 19349 3349 19383 3383
rect 8585 3145 8619 3179
rect 9781 3145 9815 3179
rect 16221 3145 16255 3179
rect 19165 3145 19199 3179
rect 12909 2601 12943 2635
rect 15715 2601 15749 2635
rect 24731 2601 24765 2635
rect 14243 2533 14277 2567
rect 10517 2465 10551 2499
rect 11069 2465 11103 2499
rect 12700 2465 12734 2499
rect 14156 2465 14190 2499
rect 15644 2465 15678 2499
rect 24660 2465 24694 2499
rect 10701 2329 10735 2363
rect 13185 2261 13219 2295
rect 14657 2261 14691 2295
rect 16129 2261 16163 2295
rect 25145 2261 25179 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 10965 24395 11023 24401
rect 10965 24361 10977 24395
rect 11011 24392 11023 24395
rect 13078 24392 13084 24404
rect 11011 24364 13084 24392
rect 11011 24361 11023 24364
rect 10965 24355 11023 24361
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 1464 24259 1522 24265
rect 1464 24225 1476 24259
rect 1510 24256 1522 24259
rect 2222 24256 2228 24268
rect 1510 24228 2228 24256
rect 1510 24225 1522 24228
rect 1464 24219 1522 24225
rect 2222 24216 2228 24228
rect 2280 24216 2286 24268
rect 8640 24259 8698 24265
rect 8640 24225 8652 24259
rect 8686 24256 8698 24259
rect 9398 24256 9404 24268
rect 8686 24228 9404 24256
rect 8686 24225 8698 24228
rect 8640 24219 8698 24225
rect 9398 24216 9404 24228
rect 9456 24216 9462 24268
rect 10778 24256 10784 24268
rect 10739 24228 10784 24256
rect 10778 24216 10784 24228
rect 10836 24216 10842 24268
rect 16482 24265 16488 24268
rect 16460 24259 16488 24265
rect 16460 24256 16472 24259
rect 16395 24228 16472 24256
rect 16460 24225 16472 24228
rect 16540 24256 16546 24268
rect 18322 24256 18328 24268
rect 16540 24228 18328 24256
rect 16460 24219 16488 24225
rect 16482 24216 16488 24219
rect 16540 24216 16546 24228
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 24648 24259 24706 24265
rect 24648 24225 24660 24259
rect 24694 24256 24706 24259
rect 25130 24256 25136 24268
rect 24694 24228 25136 24256
rect 24694 24225 24706 24228
rect 24648 24219 24706 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 1535 24055 1593 24061
rect 1535 24021 1547 24055
rect 1581 24052 1593 24055
rect 3418 24052 3424 24064
rect 1581 24024 3424 24052
rect 1581 24021 1593 24024
rect 1535 24015 1593 24021
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 8386 24052 8392 24064
rect 8347 24024 8392 24052
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 8711 24055 8769 24061
rect 8711 24021 8723 24055
rect 8757 24052 8769 24055
rect 9214 24052 9220 24064
rect 8757 24024 9220 24052
rect 8757 24021 8769 24024
rect 8711 24015 8769 24021
rect 9214 24012 9220 24024
rect 9272 24012 9278 24064
rect 10042 24052 10048 24064
rect 10003 24024 10048 24052
rect 10042 24012 10048 24024
rect 10100 24012 10106 24064
rect 14274 24012 14280 24064
rect 14332 24052 14338 24064
rect 16531 24055 16589 24061
rect 16531 24052 16543 24055
rect 14332 24024 16543 24052
rect 14332 24012 14338 24024
rect 16531 24021 16543 24024
rect 16577 24021 16589 24055
rect 16531 24015 16589 24021
rect 19978 24012 19984 24064
rect 20036 24052 20042 24064
rect 24719 24055 24777 24061
rect 24719 24052 24731 24055
rect 20036 24024 24731 24052
rect 20036 24012 20042 24024
rect 24719 24021 24731 24024
rect 24765 24021 24777 24055
rect 24719 24015 24777 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2222 23848 2228 23860
rect 2183 23820 2228 23848
rect 2222 23808 2228 23820
rect 2280 23808 2286 23860
rect 4246 23848 4252 23860
rect 4207 23820 4252 23848
rect 4246 23808 4252 23820
rect 4304 23808 4310 23860
rect 9398 23848 9404 23860
rect 9359 23820 9404 23848
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 10778 23808 10784 23860
rect 10836 23848 10842 23860
rect 10962 23848 10968 23860
rect 10836 23820 10968 23848
rect 10836 23808 10842 23820
rect 10962 23808 10968 23820
rect 11020 23808 11026 23860
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 14826 23848 14832 23860
rect 14507 23820 14832 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 14826 23808 14832 23820
rect 14884 23808 14890 23860
rect 15933 23851 15991 23857
rect 15933 23817 15945 23851
rect 15979 23848 15991 23851
rect 16574 23848 16580 23860
rect 15979 23820 16580 23848
rect 15979 23817 15991 23820
rect 15933 23811 15991 23817
rect 842 23604 848 23656
rect 900 23644 906 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 900 23616 1444 23644
rect 900 23604 906 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 3764 23647 3822 23653
rect 3764 23613 3776 23647
rect 3810 23644 3822 23647
rect 4246 23644 4252 23656
rect 3810 23616 4252 23644
rect 3810 23613 3822 23616
rect 3764 23607 3822 23613
rect 4246 23604 4252 23616
rect 4304 23604 4310 23656
rect 4617 23647 4675 23653
rect 4617 23613 4629 23647
rect 4663 23644 4675 23647
rect 5353 23647 5411 23653
rect 5353 23644 5365 23647
rect 4663 23616 5365 23644
rect 4663 23613 4675 23616
rect 4617 23607 4675 23613
rect 5353 23613 5365 23616
rect 5399 23644 5411 23647
rect 5442 23644 5448 23656
rect 5399 23616 5448 23644
rect 5399 23613 5411 23616
rect 5353 23607 5411 23613
rect 5442 23604 5448 23616
rect 5500 23604 5506 23656
rect 8297 23647 8355 23653
rect 8297 23644 8309 23647
rect 8128 23616 8309 23644
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 4430 23576 4436 23588
rect 1581 23548 3740 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 3712 23520 3740 23548
rect 4126 23548 4436 23576
rect 3694 23468 3700 23520
rect 3752 23468 3758 23520
rect 3835 23511 3893 23517
rect 3835 23477 3847 23511
rect 3881 23508 3893 23511
rect 4126 23508 4154 23548
rect 4430 23536 4436 23548
rect 4488 23536 4494 23588
rect 4706 23576 4712 23588
rect 4667 23548 4712 23576
rect 4706 23536 4712 23548
rect 4764 23536 4770 23588
rect 3881 23480 4154 23508
rect 3881 23477 3893 23480
rect 3835 23471 3893 23477
rect 6454 23468 6460 23520
rect 6512 23508 6518 23520
rect 8128 23517 8156 23616
rect 8297 23613 8309 23616
rect 8343 23613 8355 23647
rect 8297 23607 8355 23613
rect 8386 23604 8392 23656
rect 8444 23644 8450 23656
rect 8754 23644 8760 23656
rect 8444 23616 8760 23644
rect 8444 23604 8450 23616
rect 8754 23604 8760 23616
rect 8812 23604 8818 23656
rect 9674 23604 9680 23656
rect 9732 23644 9738 23656
rect 9861 23647 9919 23653
rect 9861 23644 9873 23647
rect 9732 23616 9873 23644
rect 9732 23604 9738 23616
rect 9861 23613 9873 23616
rect 9907 23644 9919 23647
rect 9953 23647 10011 23653
rect 9953 23644 9965 23647
rect 9907 23616 9965 23644
rect 9907 23613 9919 23616
rect 9861 23607 9919 23613
rect 9953 23613 9965 23616
rect 9999 23613 10011 23647
rect 9953 23607 10011 23613
rect 10042 23604 10048 23656
rect 10100 23644 10106 23656
rect 10505 23647 10563 23653
rect 10505 23644 10517 23647
rect 10100 23616 10517 23644
rect 10100 23604 10106 23616
rect 10505 23613 10517 23616
rect 10551 23644 10563 23647
rect 11974 23644 11980 23656
rect 10551 23616 11980 23644
rect 10551 23613 10563 23616
rect 10505 23607 10563 23613
rect 11974 23604 11980 23616
rect 12032 23604 12038 23656
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23613 14335 23647
rect 14277 23607 14335 23613
rect 15432 23647 15490 23653
rect 15432 23613 15444 23647
rect 15478 23644 15490 23647
rect 15948 23644 15976 23811
rect 16574 23808 16580 23820
rect 16632 23808 16638 23860
rect 20441 23851 20499 23857
rect 20441 23817 20453 23851
rect 20487 23848 20499 23851
rect 21818 23848 21824 23860
rect 20487 23820 21824 23848
rect 20487 23817 20499 23820
rect 20441 23811 20499 23817
rect 16482 23780 16488 23792
rect 16443 23752 16488 23780
rect 16482 23740 16488 23752
rect 16540 23740 16546 23792
rect 15478 23616 15976 23644
rect 16720 23647 16778 23653
rect 15478 23613 15490 23616
rect 15432 23607 15490 23613
rect 16720 23613 16732 23647
rect 16766 23644 16778 23647
rect 17218 23644 17224 23656
rect 16766 23616 17224 23644
rect 16766 23613 16778 23616
rect 16720 23607 16778 23613
rect 8113 23511 8171 23517
rect 8113 23508 8125 23511
rect 6512 23480 8125 23508
rect 6512 23468 6518 23480
rect 8113 23477 8125 23480
rect 8159 23477 8171 23511
rect 8570 23508 8576 23520
rect 8531 23480 8576 23508
rect 8113 23471 8171 23477
rect 8570 23468 8576 23480
rect 8628 23468 8634 23520
rect 10042 23508 10048 23520
rect 10003 23480 10048 23508
rect 10042 23468 10048 23480
rect 10100 23468 10106 23520
rect 14292 23508 14320 23607
rect 17218 23604 17224 23616
rect 17276 23604 17282 23656
rect 19940 23647 19998 23653
rect 19940 23613 19952 23647
rect 19986 23644 19998 23647
rect 20456 23644 20484 23811
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 25130 23848 25136 23860
rect 25043 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23848 25194 23860
rect 27062 23848 27068 23860
rect 25188 23820 27068 23848
rect 25188 23808 25194 23820
rect 27062 23808 27068 23820
rect 27120 23808 27126 23860
rect 25498 23780 25504 23792
rect 25459 23752 25504 23780
rect 25498 23740 25504 23752
rect 25556 23740 25562 23792
rect 19986 23616 20484 23644
rect 24648 23647 24706 23653
rect 19986 23613 19998 23616
rect 19940 23607 19998 23613
rect 24648 23613 24660 23647
rect 24694 23644 24706 23647
rect 25516 23644 25544 23740
rect 24694 23616 25544 23644
rect 24694 23613 24706 23616
rect 24648 23607 24706 23613
rect 14642 23536 14648 23588
rect 14700 23576 14706 23588
rect 15519 23579 15577 23585
rect 15519 23576 15531 23579
rect 14700 23548 15531 23576
rect 14700 23536 14706 23548
rect 15519 23545 15531 23548
rect 15565 23545 15577 23579
rect 15519 23539 15577 23545
rect 16298 23536 16304 23588
rect 16356 23576 16362 23588
rect 16807 23579 16865 23585
rect 16807 23576 16819 23579
rect 16356 23548 16819 23576
rect 16356 23536 16362 23548
rect 16807 23545 16819 23548
rect 16853 23545 16865 23579
rect 16807 23539 16865 23545
rect 16942 23536 16948 23588
rect 17000 23576 17006 23588
rect 20027 23579 20085 23585
rect 20027 23576 20039 23579
rect 17000 23548 20039 23576
rect 17000 23536 17006 23548
rect 20027 23545 20039 23548
rect 20073 23545 20085 23579
rect 20027 23539 20085 23545
rect 14921 23511 14979 23517
rect 14921 23508 14933 23511
rect 14292 23480 14933 23508
rect 14921 23477 14933 23480
rect 14967 23508 14979 23511
rect 16022 23508 16028 23520
rect 14967 23480 16028 23508
rect 14967 23477 14979 23480
rect 14921 23471 14979 23477
rect 16022 23468 16028 23480
rect 16080 23468 16086 23520
rect 23290 23468 23296 23520
rect 23348 23508 23354 23520
rect 24719 23511 24777 23517
rect 24719 23508 24731 23511
rect 23348 23480 24731 23508
rect 23348 23468 23354 23480
rect 24719 23477 24731 23480
rect 24765 23477 24777 23511
rect 24719 23471 24777 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 9815 23307 9873 23313
rect 9815 23273 9827 23307
rect 9861 23304 9873 23307
rect 10962 23304 10968 23316
rect 9861 23276 10968 23304
rect 9861 23273 9873 23276
rect 9815 23267 9873 23273
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 15930 23264 15936 23316
rect 15988 23304 15994 23316
rect 16301 23307 16359 23313
rect 16301 23304 16313 23307
rect 15988 23276 16313 23304
rect 15988 23264 15994 23276
rect 16301 23273 16313 23276
rect 16347 23304 16359 23307
rect 16942 23304 16948 23316
rect 16347 23276 16948 23304
rect 16347 23273 16359 23276
rect 16301 23267 16359 23273
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 13722 23236 13728 23248
rect 13683 23208 13728 23236
rect 13722 23196 13728 23208
rect 13780 23196 13786 23248
rect 1026 23128 1032 23180
rect 1084 23168 1090 23180
rect 1432 23171 1490 23177
rect 1432 23168 1444 23171
rect 1084 23140 1444 23168
rect 1084 23128 1090 23140
rect 1432 23137 1444 23140
rect 1478 23168 1490 23171
rect 1578 23168 1584 23180
rect 1478 23140 1584 23168
rect 1478 23137 1490 23140
rect 1432 23131 1490 23137
rect 1578 23128 1584 23140
rect 1636 23128 1642 23180
rect 2590 23128 2596 23180
rect 2648 23168 2654 23180
rect 2812 23171 2870 23177
rect 2812 23168 2824 23171
rect 2648 23140 2824 23168
rect 2648 23128 2654 23140
rect 2812 23137 2824 23140
rect 2858 23137 2870 23171
rect 5350 23168 5356 23180
rect 5311 23140 5356 23168
rect 2812 23131 2870 23137
rect 5350 23128 5356 23140
rect 5408 23128 5414 23180
rect 8202 23168 8208 23180
rect 8163 23140 8208 23168
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 9582 23168 9588 23180
rect 9543 23140 9588 23168
rect 9582 23128 9588 23140
rect 9640 23128 9646 23180
rect 11330 23168 11336 23180
rect 11291 23140 11336 23168
rect 11330 23128 11336 23140
rect 11388 23128 11394 23180
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 15470 23168 15476 23180
rect 15335 23140 15476 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 15470 23128 15476 23140
rect 15528 23128 15534 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 13633 23103 13691 23109
rect 13633 23100 13645 23103
rect 13556 23072 13645 23100
rect 13556 22976 13584 23072
rect 13633 23069 13645 23072
rect 13679 23069 13691 23103
rect 14550 23100 14556 23112
rect 14511 23072 14556 23100
rect 13633 23063 13691 23069
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 14185 23035 14243 23041
rect 14185 23001 14197 23035
rect 14231 23032 14243 23035
rect 16206 23032 16212 23044
rect 14231 23004 16212 23032
rect 14231 23001 14243 23004
rect 14185 22995 14243 23001
rect 16206 22992 16212 23004
rect 16264 22992 16270 23044
rect 1535 22967 1593 22973
rect 1535 22933 1547 22967
rect 1581 22964 1593 22967
rect 1854 22964 1860 22976
rect 1581 22936 1860 22964
rect 1581 22933 1593 22936
rect 1535 22927 1593 22933
rect 1854 22924 1860 22936
rect 1912 22924 1918 22976
rect 2041 22967 2099 22973
rect 2041 22933 2053 22967
rect 2087 22964 2099 22967
rect 2314 22964 2320 22976
rect 2087 22936 2320 22964
rect 2087 22933 2099 22936
rect 2041 22927 2099 22933
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 2915 22967 2973 22973
rect 2915 22933 2927 22967
rect 2961 22964 2973 22967
rect 4614 22964 4620 22976
rect 2961 22936 4620 22964
rect 2961 22933 2973 22936
rect 2915 22927 2973 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 5166 22964 5172 22976
rect 5127 22936 5172 22964
rect 5166 22924 5172 22936
rect 5224 22924 5230 22976
rect 8294 22964 8300 22976
rect 8255 22936 8300 22964
rect 8294 22924 8300 22936
rect 8352 22924 8358 22976
rect 11514 22964 11520 22976
rect 11475 22936 11520 22964
rect 11514 22924 11520 22936
rect 11572 22924 11578 22976
rect 13538 22924 13544 22976
rect 13596 22924 13602 22976
rect 15378 22924 15384 22976
rect 15436 22964 15442 22976
rect 15519 22967 15577 22973
rect 15519 22964 15531 22967
rect 15436 22936 15531 22964
rect 15436 22924 15442 22936
rect 15519 22933 15531 22936
rect 15565 22933 15577 22967
rect 15519 22927 15577 22933
rect 15746 22924 15752 22976
rect 15804 22964 15810 22976
rect 15841 22967 15899 22973
rect 15841 22964 15853 22967
rect 15804 22936 15853 22964
rect 15804 22924 15810 22936
rect 15841 22933 15853 22936
rect 15887 22933 15899 22967
rect 15841 22927 15899 22933
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 24719 22967 24777 22973
rect 24719 22964 24731 22967
rect 22152 22936 24731 22964
rect 22152 22924 22158 22936
rect 24719 22933 24731 22936
rect 24765 22933 24777 22967
rect 24719 22927 24777 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 2590 22720 2596 22772
rect 2648 22760 2654 22772
rect 2961 22763 3019 22769
rect 2961 22760 2973 22763
rect 2648 22732 2973 22760
rect 2648 22720 2654 22732
rect 2961 22729 2973 22732
rect 3007 22729 3019 22763
rect 8202 22760 8208 22772
rect 8163 22732 8208 22760
rect 2961 22723 3019 22729
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 11330 22760 11336 22772
rect 11291 22732 11336 22760
rect 11330 22720 11336 22732
rect 11388 22720 11394 22772
rect 15470 22760 15476 22772
rect 15431 22732 15476 22760
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 18693 22763 18751 22769
rect 18693 22729 18705 22763
rect 18739 22760 18751 22763
rect 20070 22760 20076 22772
rect 18739 22732 20076 22760
rect 18739 22729 18751 22732
rect 18693 22723 18751 22729
rect 3651 22695 3709 22701
rect 3651 22661 3663 22695
rect 3697 22692 3709 22695
rect 13906 22692 13912 22704
rect 3697 22664 7420 22692
rect 3697 22661 3709 22664
rect 3651 22655 3709 22661
rect 4614 22624 4620 22636
rect 4575 22596 4620 22624
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 2314 22556 2320 22568
rect 2275 22528 2320 22556
rect 2314 22516 2320 22528
rect 2372 22516 2378 22568
rect 3326 22516 3332 22568
rect 3384 22556 3390 22568
rect 3548 22559 3606 22565
rect 3548 22556 3560 22559
rect 3384 22528 3560 22556
rect 3384 22516 3390 22528
rect 3548 22525 3560 22528
rect 3594 22556 3606 22559
rect 3973 22559 4031 22565
rect 3973 22556 3985 22559
rect 3594 22528 3985 22556
rect 3594 22525 3606 22528
rect 3548 22519 3606 22525
rect 3973 22525 3985 22528
rect 4019 22525 4031 22559
rect 3973 22519 4031 22525
rect 4433 22491 4491 22497
rect 4433 22457 4445 22491
rect 4479 22488 4491 22491
rect 4706 22488 4712 22500
rect 4479 22460 4712 22488
rect 4479 22457 4491 22460
rect 4433 22451 4491 22457
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 5258 22488 5264 22500
rect 5219 22460 5264 22488
rect 5258 22448 5264 22460
rect 5316 22448 5322 22500
rect 7392 22488 7420 22664
rect 13372 22664 13912 22692
rect 8662 22584 8668 22636
rect 8720 22624 8726 22636
rect 9582 22624 9588 22636
rect 8720 22596 9588 22624
rect 8720 22584 8726 22596
rect 9582 22584 9588 22596
rect 9640 22624 9646 22636
rect 9769 22627 9827 22633
rect 9769 22624 9781 22627
rect 9640 22596 9781 22624
rect 9640 22584 9646 22596
rect 9769 22593 9781 22596
rect 9815 22593 9827 22627
rect 9769 22587 9827 22593
rect 10413 22559 10471 22565
rect 10413 22525 10425 22559
rect 10459 22525 10471 22559
rect 10413 22519 10471 22525
rect 8846 22488 8852 22500
rect 7392 22460 8852 22488
rect 8846 22448 8852 22460
rect 8904 22448 8910 22500
rect 8941 22491 8999 22497
rect 8941 22457 8953 22491
rect 8987 22457 8999 22491
rect 8941 22451 8999 22457
rect 9493 22491 9551 22497
rect 9493 22457 9505 22491
rect 9539 22488 9551 22491
rect 9582 22488 9588 22500
rect 9539 22460 9588 22488
rect 9539 22457 9551 22460
rect 9493 22451 9551 22457
rect 2222 22420 2228 22432
rect 2183 22392 2228 22420
rect 2222 22380 2228 22392
rect 2280 22380 2286 22432
rect 5350 22380 5356 22432
rect 5408 22420 5414 22432
rect 5537 22423 5595 22429
rect 5537 22420 5549 22423
rect 5408 22392 5549 22420
rect 5408 22380 5414 22392
rect 5537 22389 5549 22392
rect 5583 22389 5595 22423
rect 5537 22383 5595 22389
rect 7558 22380 7564 22432
rect 7616 22420 7622 22432
rect 7745 22423 7803 22429
rect 7745 22420 7757 22423
rect 7616 22392 7757 22420
rect 7616 22380 7622 22392
rect 7745 22389 7757 22392
rect 7791 22389 7803 22423
rect 7745 22383 7803 22389
rect 8665 22423 8723 22429
rect 8665 22389 8677 22423
rect 8711 22420 8723 22423
rect 8956 22420 8984 22451
rect 9582 22448 9588 22460
rect 9640 22448 9646 22500
rect 10321 22491 10379 22497
rect 10321 22488 10333 22491
rect 9692 22460 10333 22488
rect 9692 22420 9720 22460
rect 10321 22457 10333 22460
rect 10367 22457 10379 22491
rect 10321 22451 10379 22457
rect 10134 22420 10140 22432
rect 8711 22392 9720 22420
rect 10095 22392 10140 22420
rect 8711 22389 8723 22392
rect 8665 22383 8723 22389
rect 10134 22380 10140 22392
rect 10192 22420 10198 22432
rect 10422 22420 10450 22519
rect 12802 22516 12808 22568
rect 12860 22556 12866 22568
rect 13372 22565 13400 22664
rect 13906 22652 13912 22664
rect 13964 22692 13970 22704
rect 13964 22664 15148 22692
rect 13964 22652 13970 22664
rect 13449 22627 13507 22633
rect 13449 22593 13461 22627
rect 13495 22624 13507 22627
rect 13722 22624 13728 22636
rect 13495 22596 13728 22624
rect 13495 22593 13507 22596
rect 13449 22587 13507 22593
rect 13722 22584 13728 22596
rect 13780 22584 13786 22636
rect 14369 22627 14427 22633
rect 14369 22593 14381 22627
rect 14415 22624 14427 22627
rect 14550 22624 14556 22636
rect 14415 22596 14556 22624
rect 14415 22593 14427 22596
rect 14369 22587 14427 22593
rect 14550 22584 14556 22596
rect 14608 22584 14614 22636
rect 13357 22559 13415 22565
rect 13357 22556 13369 22559
rect 12860 22528 13369 22556
rect 12860 22516 12866 22528
rect 13357 22525 13369 22528
rect 13403 22525 13415 22559
rect 13357 22519 13415 22525
rect 14461 22491 14519 22497
rect 14461 22457 14473 22491
rect 14507 22457 14519 22491
rect 15010 22488 15016 22500
rect 14971 22460 15016 22488
rect 14461 22451 14519 22457
rect 14090 22420 14096 22432
rect 10192 22392 10450 22420
rect 14051 22392 14096 22420
rect 10192 22380 10198 22392
rect 14090 22380 14096 22392
rect 14148 22420 14154 22432
rect 14476 22420 14504 22451
rect 15010 22448 15016 22460
rect 15068 22448 15074 22500
rect 15120 22488 15148 22664
rect 15930 22624 15936 22636
rect 15891 22596 15936 22624
rect 15930 22584 15936 22596
rect 15988 22584 15994 22636
rect 16206 22624 16212 22636
rect 16167 22596 16212 22624
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 18208 22559 18266 22565
rect 18208 22525 18220 22559
rect 18254 22556 18266 22559
rect 18708 22556 18736 22723
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 24670 22760 24676 22772
rect 24631 22732 24676 22760
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 18254 22528 18736 22556
rect 18254 22525 18266 22528
rect 18208 22519 18266 22525
rect 15746 22488 15752 22500
rect 15120 22460 15752 22488
rect 15746 22448 15752 22460
rect 15804 22488 15810 22500
rect 16025 22491 16083 22497
rect 16025 22488 16037 22491
rect 15804 22460 16037 22488
rect 15804 22448 15810 22460
rect 16025 22457 16037 22460
rect 16071 22457 16083 22491
rect 16025 22451 16083 22457
rect 14148 22392 14504 22420
rect 14148 22380 14154 22392
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 18279 22423 18337 22429
rect 18279 22420 18291 22423
rect 15896 22392 18291 22420
rect 15896 22380 15902 22392
rect 18279 22389 18291 22392
rect 18325 22389 18337 22423
rect 18279 22383 18337 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 5169 22219 5227 22225
rect 5169 22185 5181 22219
rect 5215 22216 5227 22219
rect 5258 22216 5264 22228
rect 5215 22188 5264 22216
rect 5215 22185 5227 22188
rect 5169 22179 5227 22185
rect 5258 22176 5264 22188
rect 5316 22216 5322 22228
rect 5316 22188 6040 22216
rect 5316 22176 5322 22188
rect 2133 22151 2191 22157
rect 2133 22117 2145 22151
rect 2179 22148 2191 22151
rect 2222 22148 2228 22160
rect 2179 22120 2228 22148
rect 2179 22117 2191 22120
rect 2133 22111 2191 22117
rect 2222 22108 2228 22120
rect 2280 22108 2286 22160
rect 5442 22148 5448 22160
rect 5403 22120 5448 22148
rect 5442 22108 5448 22120
rect 5500 22108 5506 22160
rect 6012 22157 6040 22188
rect 8846 22176 8852 22228
rect 8904 22216 8910 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8904 22188 9045 22216
rect 8904 22176 8910 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 9490 22176 9496 22228
rect 9548 22216 9554 22228
rect 10134 22216 10140 22228
rect 9548 22188 10140 22216
rect 9548 22176 9554 22188
rect 5997 22151 6055 22157
rect 5997 22117 6009 22151
rect 6043 22117 6055 22151
rect 5997 22111 6055 22117
rect 8205 22151 8263 22157
rect 8205 22117 8217 22151
rect 8251 22148 8263 22151
rect 8294 22148 8300 22160
rect 8251 22120 8300 22148
rect 8251 22117 8263 22120
rect 8205 22111 8263 22117
rect 8294 22108 8300 22120
rect 8352 22108 8358 22160
rect 9214 22108 9220 22160
rect 9272 22148 9278 22160
rect 9766 22148 9772 22160
rect 9272 22120 9772 22148
rect 9272 22108 9278 22120
rect 9766 22108 9772 22120
rect 9824 22108 9830 22160
rect 9876 22157 9904 22188
rect 10134 22176 10140 22188
rect 10192 22176 10198 22228
rect 12802 22216 12808 22228
rect 12763 22188 12808 22216
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 13538 22216 13544 22228
rect 13499 22188 13544 22216
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 14090 22216 14096 22228
rect 14051 22188 14096 22216
rect 14090 22176 14096 22188
rect 14148 22176 14154 22228
rect 15010 22176 15016 22228
rect 15068 22216 15074 22228
rect 15746 22216 15752 22228
rect 15068 22188 15752 22216
rect 15068 22176 15074 22188
rect 15746 22176 15752 22188
rect 15804 22216 15810 22228
rect 15804 22188 16068 22216
rect 15804 22176 15810 22188
rect 9861 22151 9919 22157
rect 9861 22117 9873 22151
rect 9907 22117 9919 22151
rect 9861 22111 9919 22117
rect 11514 22108 11520 22160
rect 11572 22148 11578 22160
rect 11609 22151 11667 22157
rect 11609 22148 11621 22151
rect 11572 22120 11621 22148
rect 11572 22108 11578 22120
rect 11609 22117 11621 22120
rect 11655 22117 11667 22151
rect 15378 22148 15384 22160
rect 15339 22120 15384 22148
rect 11609 22111 11667 22117
rect 15378 22108 15384 22120
rect 15436 22108 15442 22160
rect 15470 22108 15476 22160
rect 15528 22148 15534 22160
rect 16040 22157 16068 22188
rect 16025 22151 16083 22157
rect 15528 22120 15573 22148
rect 15528 22108 15534 22120
rect 16025 22117 16037 22151
rect 16071 22117 16083 22151
rect 16025 22111 16083 22117
rect 6984 22083 7042 22089
rect 6984 22049 6996 22083
rect 7030 22080 7042 22083
rect 7098 22080 7104 22092
rect 7030 22052 7104 22080
rect 7030 22049 7042 22052
rect 6984 22043 7042 22049
rect 7098 22040 7104 22052
rect 7156 22040 7162 22092
rect 14277 22083 14335 22089
rect 14277 22049 14289 22083
rect 14323 22049 14335 22083
rect 14277 22043 14335 22049
rect 24581 22083 24639 22089
rect 24581 22049 24593 22083
rect 24627 22080 24639 22083
rect 24670 22080 24676 22092
rect 24627 22052 24676 22080
rect 24627 22049 24639 22052
rect 24581 22043 24639 22049
rect 1210 21972 1216 22024
rect 1268 22012 1274 22024
rect 2041 22015 2099 22021
rect 2041 22012 2053 22015
rect 1268 21984 2053 22012
rect 1268 21972 1274 21984
rect 2041 21981 2053 21984
rect 2087 22012 2099 22015
rect 3510 22012 3516 22024
rect 2087 21984 3516 22012
rect 2087 21981 2099 21984
rect 2041 21975 2099 21981
rect 3510 21972 3516 21984
rect 3568 21972 3574 22024
rect 4246 22012 4252 22024
rect 4207 21984 4252 22012
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 22012 5411 22015
rect 6178 22012 6184 22024
rect 5399 21984 6184 22012
rect 5399 21981 5411 21984
rect 5353 21975 5411 21981
rect 6178 21972 6184 21984
rect 6236 21972 6242 22024
rect 7558 21972 7564 22024
rect 7616 22012 7622 22024
rect 8113 22015 8171 22021
rect 8113 22012 8125 22015
rect 7616 21984 8125 22012
rect 7616 21972 7622 21984
rect 8113 21981 8125 21984
rect 8159 21981 8171 22015
rect 8113 21975 8171 21981
rect 9582 21972 9588 22024
rect 9640 22012 9646 22024
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 9640 21984 10057 22012
rect 9640 21972 9646 21984
rect 10045 21981 10057 21984
rect 10091 21981 10103 22015
rect 10045 21975 10103 21981
rect 11517 22015 11575 22021
rect 11517 21981 11529 22015
rect 11563 22012 11575 22015
rect 11790 22012 11796 22024
rect 11563 21984 11796 22012
rect 11563 21981 11575 21984
rect 11517 21975 11575 21981
rect 11790 21972 11796 21984
rect 11848 22012 11854 22024
rect 11848 21984 12388 22012
rect 11848 21972 11854 21984
rect 2593 21947 2651 21953
rect 2593 21913 2605 21947
rect 2639 21944 2651 21947
rect 2774 21944 2780 21956
rect 2639 21916 2780 21944
rect 2639 21913 2651 21916
rect 2593 21907 2651 21913
rect 2774 21904 2780 21916
rect 2832 21944 2838 21956
rect 7834 21944 7840 21956
rect 2832 21916 7840 21944
rect 2832 21904 2838 21916
rect 7834 21904 7840 21916
rect 7892 21904 7898 21956
rect 8662 21944 8668 21956
rect 8623 21916 8668 21944
rect 8662 21904 8668 21916
rect 8720 21904 8726 21956
rect 12069 21947 12127 21953
rect 12069 21913 12081 21947
rect 12115 21944 12127 21947
rect 12250 21944 12256 21956
rect 12115 21916 12256 21944
rect 12115 21913 12127 21916
rect 12069 21907 12127 21913
rect 12250 21904 12256 21916
rect 12308 21904 12314 21956
rect 12360 21944 12388 21984
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 14292 22012 14320 22043
rect 24670 22040 24676 22052
rect 24728 22040 24734 22092
rect 14458 22012 14464 22024
rect 13780 21984 14464 22012
rect 13780 21972 13786 21984
rect 14458 21972 14464 21984
rect 14516 22012 14522 22024
rect 15470 22012 15476 22024
rect 14516 21984 15476 22012
rect 14516 21972 14522 21984
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 15838 21944 15844 21956
rect 12360 21916 15844 21944
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 4338 21836 4344 21888
rect 4396 21876 4402 21888
rect 5534 21876 5540 21888
rect 4396 21848 5540 21876
rect 4396 21836 4402 21848
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 7055 21879 7113 21885
rect 7055 21876 7067 21879
rect 6880 21848 7067 21876
rect 6880 21836 6886 21848
rect 7055 21845 7067 21848
rect 7101 21845 7113 21879
rect 10870 21876 10876 21888
rect 10831 21848 10876 21876
rect 7055 21839 7113 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 18598 21836 18604 21888
rect 18656 21876 18662 21888
rect 24719 21879 24777 21885
rect 24719 21876 24731 21879
rect 18656 21848 24731 21876
rect 18656 21836 18662 21848
rect 24719 21845 24731 21848
rect 24765 21845 24777 21879
rect 24719 21839 24777 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2041 21675 2099 21681
rect 2041 21641 2053 21675
rect 2087 21672 2099 21675
rect 2222 21672 2228 21684
rect 2087 21644 2228 21672
rect 2087 21641 2099 21644
rect 2041 21635 2099 21641
rect 2222 21632 2228 21644
rect 2280 21632 2286 21684
rect 3510 21672 3516 21684
rect 3471 21644 3516 21672
rect 3510 21632 3516 21644
rect 3568 21632 3574 21684
rect 3878 21672 3884 21684
rect 3839 21644 3884 21672
rect 3878 21632 3884 21644
rect 3936 21632 3942 21684
rect 5442 21632 5448 21684
rect 5500 21672 5506 21684
rect 6089 21675 6147 21681
rect 6089 21672 6101 21675
rect 5500 21644 6101 21672
rect 5500 21632 5506 21644
rect 6089 21641 6101 21644
rect 6135 21641 6147 21675
rect 6089 21635 6147 21641
rect 7009 21675 7067 21681
rect 7009 21641 7021 21675
rect 7055 21672 7067 21675
rect 7650 21672 7656 21684
rect 7055 21644 7656 21672
rect 7055 21641 7067 21644
rect 7009 21635 7067 21641
rect 7650 21632 7656 21644
rect 7708 21632 7714 21684
rect 7929 21675 7987 21681
rect 7929 21641 7941 21675
rect 7975 21672 7987 21675
rect 8294 21672 8300 21684
rect 7975 21644 8300 21672
rect 7975 21641 7987 21644
rect 7929 21635 7987 21641
rect 8294 21632 8300 21644
rect 8352 21632 8358 21684
rect 10321 21675 10379 21681
rect 10321 21641 10333 21675
rect 10367 21672 10379 21675
rect 11054 21672 11060 21684
rect 10367 21644 11060 21672
rect 10367 21641 10379 21644
rect 10321 21635 10379 21641
rect 2774 21604 2780 21616
rect 2735 21576 2780 21604
rect 2774 21564 2780 21576
rect 2832 21564 2838 21616
rect 7558 21604 7564 21616
rect 7519 21576 7564 21604
rect 7558 21564 7564 21576
rect 7616 21564 7622 21616
rect 8662 21604 8668 21616
rect 8623 21576 8668 21604
rect 8662 21564 8668 21576
rect 8720 21564 8726 21616
rect 10336 21604 10364 21635
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11514 21632 11520 21684
rect 11572 21672 11578 21684
rect 11793 21675 11851 21681
rect 11793 21672 11805 21675
rect 11572 21644 11805 21672
rect 11572 21632 11578 21644
rect 11793 21641 11805 21644
rect 11839 21641 11851 21675
rect 13722 21672 13728 21684
rect 13683 21644 13728 21672
rect 11793 21635 11851 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 14461 21675 14519 21681
rect 14461 21641 14473 21675
rect 14507 21672 14519 21675
rect 15378 21672 15384 21684
rect 14507 21644 15384 21672
rect 14507 21641 14519 21644
rect 14461 21635 14519 21641
rect 15378 21632 15384 21644
rect 15436 21632 15442 21684
rect 15470 21632 15476 21684
rect 15528 21672 15534 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 15528 21644 15945 21672
rect 15528 21632 15534 21644
rect 15933 21641 15945 21644
rect 15979 21641 15991 21675
rect 15933 21635 15991 21641
rect 16022 21632 16028 21684
rect 16080 21672 16086 21684
rect 16623 21675 16681 21681
rect 16623 21672 16635 21675
rect 16080 21644 16635 21672
rect 16080 21632 16086 21644
rect 16623 21641 16635 21644
rect 16669 21641 16681 21675
rect 24670 21672 24676 21684
rect 24631 21644 24676 21672
rect 16623 21635 16681 21641
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 9830 21576 10364 21604
rect 1854 21496 1860 21548
rect 1912 21536 1918 21548
rect 2225 21539 2283 21545
rect 2225 21536 2237 21539
rect 1912 21508 2237 21536
rect 1912 21496 1918 21508
rect 2225 21505 2237 21508
rect 2271 21536 2283 21539
rect 3145 21539 3203 21545
rect 3145 21536 3157 21539
rect 2271 21508 3157 21536
rect 2271 21505 2283 21508
rect 2225 21499 2283 21505
rect 3145 21505 3157 21508
rect 3191 21505 3203 21539
rect 3145 21499 3203 21505
rect 5169 21539 5227 21545
rect 5169 21505 5181 21539
rect 5215 21536 5227 21539
rect 5258 21536 5264 21548
rect 5215 21508 5264 21536
rect 5215 21505 5227 21508
rect 5169 21499 5227 21505
rect 5258 21496 5264 21508
rect 5316 21496 5322 21548
rect 5534 21536 5540 21548
rect 5495 21508 5540 21536
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 7834 21496 7840 21548
rect 7892 21536 7898 21548
rect 8113 21539 8171 21545
rect 8113 21536 8125 21539
rect 7892 21508 8125 21536
rect 7892 21496 7898 21508
rect 8113 21505 8125 21508
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 3694 21468 3700 21480
rect 3655 21440 3700 21468
rect 3694 21428 3700 21440
rect 3752 21468 3758 21480
rect 4249 21471 4307 21477
rect 4249 21468 4261 21471
rect 3752 21440 4261 21468
rect 3752 21428 3758 21440
rect 4249 21437 4261 21440
rect 4295 21437 4307 21471
rect 6822 21468 6828 21480
rect 6783 21440 6828 21468
rect 4249 21431 4307 21437
rect 6822 21428 6828 21440
rect 6880 21428 6886 21480
rect 9830 21477 9858 21576
rect 9907 21539 9965 21545
rect 9907 21505 9919 21539
rect 9953 21536 9965 21539
rect 10870 21536 10876 21548
rect 9953 21508 10876 21536
rect 9953 21505 9965 21508
rect 9907 21499 9965 21505
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 9815 21471 9873 21477
rect 9815 21437 9827 21471
rect 9861 21437 9873 21471
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 9815 21431 9873 21437
rect 12360 21440 12449 21468
rect 1673 21403 1731 21409
rect 1673 21369 1685 21403
rect 1719 21400 1731 21403
rect 2314 21400 2320 21412
rect 1719 21372 2320 21400
rect 1719 21369 1731 21372
rect 1673 21363 1731 21369
rect 2314 21360 2320 21372
rect 2372 21400 2378 21412
rect 3326 21400 3332 21412
rect 2372 21372 3332 21400
rect 2372 21360 2378 21372
rect 3326 21360 3332 21372
rect 3384 21360 3390 21412
rect 4985 21403 5043 21409
rect 4985 21369 4997 21403
rect 5031 21400 5043 21403
rect 5258 21400 5264 21412
rect 5031 21372 5264 21400
rect 5031 21369 5043 21372
rect 4985 21363 5043 21369
rect 5258 21360 5264 21372
rect 5316 21360 5322 21412
rect 8202 21400 8208 21412
rect 8163 21372 8208 21400
rect 8202 21360 8208 21372
rect 8260 21400 8266 21412
rect 9033 21403 9091 21409
rect 9033 21400 9045 21403
rect 8260 21372 9045 21400
rect 8260 21360 8266 21372
rect 9033 21369 9045 21372
rect 9079 21369 9091 21403
rect 9033 21363 9091 21369
rect 10689 21403 10747 21409
rect 10689 21369 10701 21403
rect 10735 21400 10747 21403
rect 10965 21403 11023 21409
rect 10965 21400 10977 21403
rect 10735 21372 10977 21400
rect 10735 21369 10747 21372
rect 10689 21363 10747 21369
rect 10965 21369 10977 21372
rect 11011 21400 11023 21403
rect 11330 21400 11336 21412
rect 11011 21372 11336 21400
rect 11011 21369 11023 21372
rect 10965 21363 11023 21369
rect 11330 21360 11336 21372
rect 11388 21360 11394 21412
rect 11517 21403 11575 21409
rect 11517 21369 11529 21403
rect 11563 21400 11575 21403
rect 12250 21400 12256 21412
rect 11563 21372 12256 21400
rect 11563 21369 11575 21372
rect 11517 21363 11575 21369
rect 12250 21360 12256 21372
rect 12308 21360 12314 21412
rect 12360 21344 12388 21440
rect 12437 21437 12449 21440
rect 12483 21437 12495 21471
rect 12894 21468 12900 21480
rect 12855 21440 12900 21468
rect 12437 21431 12495 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 16520 21471 16578 21477
rect 16520 21437 16532 21471
rect 16566 21437 16578 21471
rect 16520 21431 16578 21437
rect 14826 21360 14832 21412
rect 14884 21400 14890 21412
rect 15013 21403 15071 21409
rect 15013 21400 15025 21403
rect 14884 21372 15025 21400
rect 14884 21360 14890 21372
rect 15013 21369 15025 21372
rect 15059 21369 15071 21403
rect 15013 21363 15071 21369
rect 15105 21403 15163 21409
rect 15105 21369 15117 21403
rect 15151 21369 15163 21403
rect 15654 21400 15660 21412
rect 15615 21372 15660 21400
rect 15105 21363 15163 21369
rect 6641 21335 6699 21341
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 7098 21332 7104 21344
rect 6687 21304 7104 21332
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 9490 21292 9496 21344
rect 9548 21332 9554 21344
rect 9585 21335 9643 21341
rect 9585 21332 9597 21335
rect 9548 21304 9597 21332
rect 9548 21292 9554 21304
rect 9585 21301 9597 21304
rect 9631 21301 9643 21335
rect 9585 21295 9643 21301
rect 12161 21335 12219 21341
rect 12161 21301 12173 21335
rect 12207 21332 12219 21335
rect 12342 21332 12348 21344
rect 12207 21304 12348 21332
rect 12207 21301 12219 21304
rect 12161 21295 12219 21301
rect 12342 21292 12348 21304
rect 12400 21292 12406 21344
rect 12526 21332 12532 21344
rect 12487 21304 12532 21332
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 14737 21335 14795 21341
rect 14737 21301 14749 21335
rect 14783 21332 14795 21335
rect 15120 21332 15148 21363
rect 15654 21360 15660 21372
rect 15712 21400 15718 21412
rect 16535 21400 16563 21431
rect 16945 21403 17003 21409
rect 16945 21400 16957 21403
rect 15712 21372 16957 21400
rect 15712 21360 15718 21372
rect 16945 21369 16957 21372
rect 16991 21369 17003 21403
rect 16945 21363 17003 21369
rect 15562 21332 15568 21344
rect 14783 21304 15568 21332
rect 14783 21301 14795 21304
rect 14737 21295 14795 21301
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 5442 21088 5448 21140
rect 5500 21128 5506 21140
rect 5813 21131 5871 21137
rect 5813 21128 5825 21131
rect 5500 21100 5825 21128
rect 5500 21088 5506 21100
rect 5813 21097 5825 21100
rect 5859 21097 5871 21131
rect 5813 21091 5871 21097
rect 6822 21088 6828 21140
rect 6880 21128 6886 21140
rect 7193 21131 7251 21137
rect 7193 21128 7205 21131
rect 6880 21100 7205 21128
rect 6880 21088 6886 21100
rect 7193 21097 7205 21100
rect 7239 21097 7251 21131
rect 7926 21128 7932 21140
rect 7887 21100 7932 21128
rect 7193 21091 7251 21097
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 8202 21088 8208 21140
rect 8260 21128 8266 21140
rect 8481 21131 8539 21137
rect 8481 21128 8493 21131
rect 8260 21100 8493 21128
rect 8260 21088 8266 21100
rect 8481 21097 8493 21100
rect 8527 21097 8539 21131
rect 8481 21091 8539 21097
rect 8570 21088 8576 21140
rect 8628 21128 8634 21140
rect 8757 21131 8815 21137
rect 8757 21128 8769 21131
rect 8628 21100 8769 21128
rect 8628 21088 8634 21100
rect 8757 21097 8769 21100
rect 8803 21097 8815 21131
rect 8757 21091 8815 21097
rect 9766 21088 9772 21140
rect 9824 21128 9830 21140
rect 9861 21131 9919 21137
rect 9861 21128 9873 21131
rect 9824 21100 9873 21128
rect 9824 21088 9830 21100
rect 9861 21097 9873 21100
rect 9907 21097 9919 21131
rect 9861 21091 9919 21097
rect 11330 21088 11336 21140
rect 11388 21128 11394 21140
rect 11425 21131 11483 21137
rect 11425 21128 11437 21131
rect 11388 21100 11437 21128
rect 11388 21088 11394 21100
rect 11425 21097 11437 21100
rect 11471 21097 11483 21131
rect 11790 21128 11796 21140
rect 11751 21100 11796 21128
rect 11425 21091 11483 21097
rect 11790 21088 11796 21100
rect 11848 21088 11854 21140
rect 13906 21128 13912 21140
rect 13867 21100 13912 21128
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 15488 21100 16988 21128
rect 15488 21072 15516 21100
rect 2038 21060 2044 21072
rect 1999 21032 2044 21060
rect 2038 21020 2044 21032
rect 2096 21020 2102 21072
rect 5255 21063 5313 21069
rect 5255 21029 5267 21063
rect 5301 21060 5313 21063
rect 5350 21060 5356 21072
rect 5301 21032 5356 21060
rect 5301 21029 5313 21032
rect 5255 21023 5313 21029
rect 5350 21020 5356 21032
rect 5408 21020 5414 21072
rect 10594 21020 10600 21072
rect 10652 21060 10658 21072
rect 10867 21063 10925 21069
rect 10867 21060 10879 21063
rect 10652 21032 10879 21060
rect 10652 21020 10658 21032
rect 10867 21029 10879 21032
rect 10913 21060 10925 21063
rect 13351 21063 13409 21069
rect 13351 21060 13363 21063
rect 10913 21032 13363 21060
rect 10913 21029 10925 21032
rect 10867 21023 10925 21029
rect 13351 21029 13363 21032
rect 13397 21060 13409 21063
rect 13446 21060 13452 21072
rect 13397 21032 13452 21060
rect 13397 21029 13409 21032
rect 13351 21023 13409 21029
rect 13446 21020 13452 21032
rect 13504 21020 13510 21072
rect 15470 21060 15476 21072
rect 15431 21032 15476 21060
rect 15470 21020 15476 21032
rect 15528 21020 15534 21072
rect 15562 21020 15568 21072
rect 15620 21060 15626 21072
rect 16853 21063 16911 21069
rect 16853 21060 16865 21063
rect 15620 21032 16865 21060
rect 15620 21020 15626 21032
rect 16853 21029 16865 21032
rect 16899 21029 16911 21063
rect 16853 21023 16911 21029
rect 2958 20992 2964 21004
rect 2871 20964 2964 20992
rect 2958 20952 2964 20964
rect 3016 20992 3022 21004
rect 8478 20992 8484 21004
rect 3016 20964 8484 20992
rect 3016 20952 3022 20964
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 10226 20952 10232 21004
rect 10284 20992 10290 21004
rect 10505 20995 10563 21001
rect 10505 20992 10517 20995
rect 10284 20964 10517 20992
rect 10284 20952 10290 20964
rect 10505 20961 10517 20964
rect 10551 20992 10563 20995
rect 12526 20992 12532 21004
rect 10551 20964 12532 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 12526 20952 12532 20964
rect 12584 20952 12590 21004
rect 16960 21001 16988 21100
rect 16945 20995 17003 21001
rect 16945 20961 16957 20995
rect 16991 20992 17003 20995
rect 17218 20992 17224 21004
rect 16991 20964 17224 20992
rect 16991 20961 17003 20964
rect 16945 20955 17003 20961
rect 17218 20952 17224 20964
rect 17276 20952 17282 21004
rect 1946 20924 1952 20936
rect 1907 20896 1952 20924
rect 1946 20884 1952 20896
rect 2004 20884 2010 20936
rect 2590 20924 2596 20936
rect 2551 20896 2596 20924
rect 2590 20884 2596 20896
rect 2648 20884 2654 20936
rect 4890 20924 4896 20936
rect 4851 20896 4896 20924
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 7558 20924 7564 20936
rect 7519 20896 7564 20924
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 12986 20924 12992 20936
rect 12947 20896 12992 20924
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 15378 20924 15384 20936
rect 15339 20896 15384 20924
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 15654 20924 15660 20936
rect 15615 20896 15660 20924
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 1670 20788 1676 20800
rect 1583 20760 1676 20788
rect 1670 20748 1676 20760
rect 1728 20788 1734 20800
rect 5534 20788 5540 20800
rect 1728 20760 5540 20788
rect 1728 20748 1734 20760
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 6178 20788 6184 20800
rect 6139 20760 6184 20788
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 6917 20791 6975 20797
rect 6917 20757 6929 20791
rect 6963 20788 6975 20791
rect 7466 20788 7472 20800
rect 6963 20760 7472 20788
rect 6963 20757 6975 20760
rect 6917 20751 6975 20757
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 11974 20748 11980 20800
rect 12032 20788 12038 20800
rect 12437 20791 12495 20797
rect 12437 20788 12449 20791
rect 12032 20760 12449 20788
rect 12032 20748 12038 20760
rect 12437 20757 12449 20760
rect 12483 20788 12495 20791
rect 12894 20788 12900 20800
rect 12483 20760 12900 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 14182 20748 14188 20800
rect 14240 20788 14246 20800
rect 14826 20788 14832 20800
rect 14240 20760 14832 20788
rect 14240 20748 14246 20760
rect 14826 20748 14832 20760
rect 14884 20788 14890 20800
rect 14921 20791 14979 20797
rect 14921 20788 14933 20791
rect 14884 20760 14933 20788
rect 14884 20748 14890 20760
rect 14921 20757 14933 20760
rect 14967 20757 14979 20791
rect 14921 20751 14979 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 3326 20584 3332 20596
rect 3287 20556 3332 20584
rect 3326 20544 3332 20556
rect 3384 20544 3390 20596
rect 5258 20544 5264 20596
rect 5316 20584 5322 20596
rect 5813 20587 5871 20593
rect 5813 20584 5825 20587
rect 5316 20556 5825 20584
rect 5316 20544 5322 20556
rect 5813 20553 5825 20556
rect 5859 20553 5871 20587
rect 9490 20584 9496 20596
rect 9451 20556 9496 20584
rect 5813 20547 5871 20553
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 10226 20584 10232 20596
rect 10187 20556 10232 20584
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 14458 20584 14464 20596
rect 14419 20556 14464 20584
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 17218 20584 17224 20596
rect 17179 20556 17224 20584
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 4065 20519 4123 20525
rect 4065 20485 4077 20519
rect 4111 20516 4123 20519
rect 4890 20516 4896 20528
rect 4111 20488 4896 20516
rect 4111 20485 4123 20488
rect 4065 20479 4123 20485
rect 4890 20476 4896 20488
rect 4948 20476 4954 20528
rect 7926 20516 7932 20528
rect 7839 20488 7932 20516
rect 7926 20476 7932 20488
rect 7984 20516 7990 20528
rect 8481 20519 8539 20525
rect 8481 20516 8493 20519
rect 7984 20488 8493 20516
rect 7984 20476 7990 20488
rect 8481 20485 8493 20488
rect 8527 20516 8539 20519
rect 10594 20516 10600 20528
rect 8527 20488 10600 20516
rect 8527 20485 8539 20488
rect 8481 20479 8539 20485
rect 2409 20451 2467 20457
rect 2409 20417 2421 20451
rect 2455 20448 2467 20451
rect 2958 20448 2964 20460
rect 2455 20420 2964 20448
rect 2455 20417 2467 20420
rect 2409 20411 2467 20417
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 8570 20448 8576 20460
rect 8531 20420 8576 20448
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 1464 20383 1522 20389
rect 1464 20349 1476 20383
rect 1510 20380 1522 20383
rect 1670 20380 1676 20392
rect 1510 20352 1676 20380
rect 1510 20349 1522 20352
rect 1464 20343 1522 20349
rect 1670 20340 1676 20352
rect 1728 20340 1734 20392
rect 1949 20383 2007 20389
rect 1949 20349 1961 20383
rect 1995 20380 2007 20383
rect 2038 20380 2044 20392
rect 1995 20352 2044 20380
rect 1995 20349 2007 20352
rect 1949 20343 2007 20349
rect 2038 20340 2044 20352
rect 2096 20380 2102 20392
rect 4798 20380 4804 20392
rect 2096 20352 4804 20380
rect 2096 20340 2102 20352
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 4893 20383 4951 20389
rect 4893 20349 4905 20383
rect 4939 20380 4951 20383
rect 6641 20383 6699 20389
rect 4939 20352 6224 20380
rect 4939 20349 4951 20352
rect 4893 20343 4951 20349
rect 2317 20315 2375 20321
rect 2317 20281 2329 20315
rect 2363 20312 2375 20315
rect 2406 20312 2412 20324
rect 2363 20284 2412 20312
rect 2363 20281 2375 20284
rect 2317 20275 2375 20281
rect 2406 20272 2412 20284
rect 2464 20312 2470 20324
rect 2771 20315 2829 20321
rect 2771 20312 2783 20315
rect 2464 20284 2783 20312
rect 2464 20272 2470 20284
rect 2771 20281 2783 20284
rect 2817 20312 2829 20315
rect 4433 20315 4491 20321
rect 4433 20312 4445 20315
rect 2817 20284 3464 20312
rect 2817 20281 2829 20284
rect 2771 20275 2829 20281
rect 1670 20244 1676 20256
rect 1631 20216 1676 20244
rect 1670 20204 1676 20216
rect 1728 20204 1734 20256
rect 3436 20244 3464 20284
rect 4126 20284 4445 20312
rect 4126 20244 4154 20284
rect 4433 20281 4445 20284
rect 4479 20312 4491 20315
rect 4709 20315 4767 20321
rect 4709 20312 4721 20315
rect 4479 20284 4721 20312
rect 4479 20281 4491 20284
rect 4433 20275 4491 20281
rect 4709 20281 4721 20284
rect 4755 20312 4767 20315
rect 5255 20315 5313 20321
rect 5255 20312 5267 20315
rect 4755 20284 5267 20312
rect 4755 20281 4767 20284
rect 4709 20275 4767 20281
rect 5255 20281 5267 20284
rect 5301 20312 5313 20315
rect 5350 20312 5356 20324
rect 5301 20284 5356 20312
rect 5301 20281 5313 20284
rect 5255 20275 5313 20281
rect 5350 20272 5356 20284
rect 5408 20272 5414 20324
rect 6196 20321 6224 20352
rect 6641 20349 6653 20383
rect 6687 20380 6699 20383
rect 7101 20383 7159 20389
rect 7101 20380 7113 20383
rect 6687 20352 7113 20380
rect 6687 20349 6699 20352
rect 6641 20343 6699 20349
rect 7101 20349 7113 20352
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 7377 20383 7435 20389
rect 7377 20349 7389 20383
rect 7423 20380 7435 20383
rect 7466 20380 7472 20392
rect 7423 20352 7472 20380
rect 7423 20349 7435 20352
rect 7377 20343 7435 20349
rect 6181 20315 6239 20321
rect 6181 20281 6193 20315
rect 6227 20312 6239 20315
rect 7116 20312 7144 20343
rect 7466 20340 7472 20352
rect 7524 20340 7530 20392
rect 7926 20312 7932 20324
rect 6227 20284 6684 20312
rect 7116 20284 7932 20312
rect 6227 20281 6239 20284
rect 6181 20275 6239 20281
rect 3436 20216 4154 20244
rect 6656 20244 6684 20284
rect 7926 20272 7932 20284
rect 7984 20272 7990 20324
rect 8909 20321 8937 20488
rect 10594 20476 10600 20488
rect 10652 20476 10658 20528
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 16298 20448 16304 20460
rect 15795 20420 16304 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 9861 20383 9919 20389
rect 9861 20349 9873 20383
rect 9907 20380 9919 20383
rect 10781 20383 10839 20389
rect 10781 20380 10793 20383
rect 9907 20352 10793 20380
rect 9907 20349 9919 20352
rect 9861 20343 9919 20349
rect 10781 20349 10793 20352
rect 10827 20380 10839 20383
rect 11330 20380 11336 20392
rect 10827 20352 11336 20380
rect 10827 20349 10839 20352
rect 10781 20343 10839 20349
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 13354 20340 13360 20392
rect 13412 20380 13418 20392
rect 13541 20383 13599 20389
rect 13541 20380 13553 20383
rect 13412 20352 13553 20380
rect 13412 20340 13418 20352
rect 13541 20349 13553 20352
rect 13587 20349 13599 20383
rect 13541 20343 13599 20349
rect 8894 20315 8952 20321
rect 8894 20281 8906 20315
rect 8940 20281 8952 20315
rect 10594 20312 10600 20324
rect 10555 20284 10600 20312
rect 8894 20275 8952 20281
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 13862 20315 13920 20321
rect 13862 20312 13874 20315
rect 13464 20284 13874 20312
rect 13464 20256 13492 20284
rect 13862 20281 13874 20284
rect 13908 20281 13920 20315
rect 13862 20275 13920 20281
rect 15013 20315 15071 20321
rect 15013 20281 15025 20315
rect 15059 20312 15071 20315
rect 15378 20312 15384 20324
rect 15059 20284 15384 20312
rect 15059 20281 15071 20284
rect 15013 20275 15071 20281
rect 15378 20272 15384 20284
rect 15436 20312 15442 20324
rect 16117 20315 16175 20321
rect 15436 20284 16068 20312
rect 15436 20272 15442 20284
rect 6917 20247 6975 20253
rect 6917 20244 6929 20247
rect 6656 20216 6929 20244
rect 6917 20213 6929 20216
rect 6963 20213 6975 20247
rect 10962 20244 10968 20256
rect 10923 20216 10968 20244
rect 6917 20207 6975 20213
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 12437 20247 12495 20253
rect 12437 20244 12449 20247
rect 11112 20216 12449 20244
rect 11112 20204 11118 20216
rect 12437 20213 12449 20216
rect 12483 20213 12495 20247
rect 12437 20207 12495 20213
rect 13081 20247 13139 20253
rect 13081 20213 13093 20247
rect 13127 20244 13139 20247
rect 13446 20244 13452 20256
rect 13127 20216 13452 20244
rect 13127 20213 13139 20216
rect 13081 20207 13139 20213
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 14884 20216 15301 20244
rect 14884 20204 14890 20216
rect 15289 20213 15301 20216
rect 15335 20244 15347 20247
rect 15470 20244 15476 20256
rect 15335 20216 15476 20244
rect 15335 20213 15347 20216
rect 15289 20207 15347 20213
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 16040 20244 16068 20284
rect 16117 20281 16129 20315
rect 16163 20312 16175 20315
rect 16390 20312 16396 20324
rect 16163 20284 16396 20312
rect 16163 20281 16175 20284
rect 16117 20275 16175 20281
rect 16390 20272 16396 20284
rect 16448 20272 16454 20324
rect 16945 20315 17003 20321
rect 16945 20281 16957 20315
rect 16991 20312 17003 20315
rect 17586 20312 17592 20324
rect 16991 20284 17592 20312
rect 16991 20281 17003 20284
rect 16945 20275 17003 20281
rect 16960 20244 16988 20275
rect 17586 20272 17592 20284
rect 17644 20272 17650 20324
rect 16040 20216 16988 20244
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 4890 20000 4896 20052
rect 4948 20040 4954 20052
rect 6549 20043 6607 20049
rect 6549 20040 6561 20043
rect 4948 20012 6561 20040
rect 4948 20000 4954 20012
rect 6549 20009 6561 20012
rect 6595 20009 6607 20043
rect 7558 20040 7564 20052
rect 7519 20012 7564 20040
rect 6549 20003 6607 20009
rect 7558 20000 7564 20012
rect 7616 20040 7622 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7616 20012 8125 20040
rect 7616 20000 7622 20012
rect 8113 20009 8125 20012
rect 8159 20009 8171 20043
rect 8113 20003 8171 20009
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10229 20043 10287 20049
rect 10229 20040 10241 20043
rect 10100 20012 10241 20040
rect 10100 20000 10106 20012
rect 10229 20009 10241 20012
rect 10275 20009 10287 20043
rect 10229 20003 10287 20009
rect 2409 19975 2467 19981
rect 2409 19941 2421 19975
rect 2455 19972 2467 19975
rect 2498 19972 2504 19984
rect 2455 19944 2504 19972
rect 2455 19941 2467 19944
rect 2409 19935 2467 19941
rect 2498 19932 2504 19944
rect 2556 19932 2562 19984
rect 4246 19932 4252 19984
rect 4304 19972 4310 19984
rect 4982 19972 4988 19984
rect 4304 19944 4988 19972
rect 4304 19932 4310 19944
rect 4982 19932 4988 19944
rect 5040 19932 5046 19984
rect 5077 19975 5135 19981
rect 5077 19941 5089 19975
rect 5123 19972 5135 19975
rect 5166 19972 5172 19984
rect 5123 19944 5172 19972
rect 5123 19941 5135 19944
rect 5077 19935 5135 19941
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 6454 19904 6460 19916
rect 6415 19876 6460 19904
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 7009 19907 7067 19913
rect 7009 19873 7021 19907
rect 7055 19904 7067 19907
rect 7466 19904 7472 19916
rect 7055 19876 7472 19904
rect 7055 19873 7067 19876
rect 7009 19867 7067 19873
rect 7466 19864 7472 19876
rect 7524 19864 7530 19916
rect 8018 19904 8024 19916
rect 7979 19876 8024 19904
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19904 8631 19907
rect 8846 19904 8852 19916
rect 8619 19876 8852 19904
rect 8619 19873 8631 19876
rect 8573 19867 8631 19873
rect 2314 19836 2320 19848
rect 2275 19808 2320 19836
rect 2314 19796 2320 19808
rect 2372 19796 2378 19848
rect 2590 19836 2596 19848
rect 2551 19808 2596 19836
rect 2590 19796 2596 19808
rect 2648 19796 2654 19848
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 8588 19836 8616 19867
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 10244 19904 10272 20003
rect 10686 20000 10692 20052
rect 10744 20040 10750 20052
rect 10781 20043 10839 20049
rect 10781 20040 10793 20043
rect 10744 20012 10793 20040
rect 10744 20000 10750 20012
rect 10781 20009 10793 20012
rect 10827 20009 10839 20043
rect 11330 20040 11336 20052
rect 11291 20012 11336 20040
rect 10781 20003 10839 20009
rect 11330 20000 11336 20012
rect 11388 20040 11394 20052
rect 11388 20012 12388 20040
rect 11388 20000 11394 20012
rect 12360 19981 12388 20012
rect 12986 20000 12992 20052
rect 13044 20040 13050 20052
rect 13173 20043 13231 20049
rect 13173 20040 13185 20043
rect 13044 20012 13185 20040
rect 13044 20000 13050 20012
rect 13173 20009 13185 20012
rect 13219 20009 13231 20043
rect 14182 20040 14188 20052
rect 14143 20012 14188 20040
rect 13173 20003 13231 20009
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 12345 19975 12403 19981
rect 12345 19941 12357 19975
rect 12391 19941 12403 19975
rect 12345 19935 12403 19941
rect 15378 19932 15384 19984
rect 15436 19972 15442 19984
rect 15610 19975 15668 19981
rect 15610 19972 15622 19975
rect 15436 19944 15622 19972
rect 15436 19932 15442 19944
rect 15610 19941 15622 19944
rect 15656 19941 15668 19975
rect 15610 19935 15668 19941
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 17221 19975 17279 19981
rect 17221 19972 17233 19975
rect 17184 19944 17233 19972
rect 17184 19932 17190 19944
rect 17221 19941 17233 19944
rect 17267 19972 17279 19975
rect 18601 19975 18659 19981
rect 18601 19972 18613 19975
rect 17267 19944 18613 19972
rect 17267 19941 17279 19944
rect 17221 19935 17279 19941
rect 18601 19941 18613 19944
rect 18647 19941 18659 19975
rect 18601 19935 18659 19941
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 10244 19876 10425 19904
rect 10413 19873 10425 19876
rect 10459 19873 10471 19907
rect 18690 19904 18696 19916
rect 18651 19876 18696 19904
rect 10413 19867 10471 19873
rect 18690 19864 18696 19876
rect 18748 19864 18754 19916
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19904 24639 19907
rect 24670 19904 24676 19916
rect 24627 19876 24676 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 12250 19836 12256 19848
rect 7975 19808 8616 19836
rect 12211 19808 12256 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 12250 19796 12256 19808
rect 12308 19796 12314 19848
rect 12526 19836 12532 19848
rect 12487 19808 12532 19836
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 15286 19836 15292 19848
rect 15247 19808 15292 19836
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 17129 19839 17187 19845
rect 17129 19805 17141 19839
rect 17175 19836 17187 19839
rect 17494 19836 17500 19848
rect 17175 19808 17500 19836
rect 17175 19805 17187 19808
rect 17129 19799 17187 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 17586 19796 17592 19848
rect 17644 19836 17650 19848
rect 17644 19808 17689 19836
rect 17644 19796 17650 19808
rect 5534 19768 5540 19780
rect 5495 19740 5540 19768
rect 5534 19728 5540 19740
rect 5592 19728 5598 19780
rect 1394 19660 1400 19712
rect 1452 19700 1458 19712
rect 1857 19703 1915 19709
rect 1857 19700 1869 19703
rect 1452 19672 1869 19700
rect 1452 19660 1458 19672
rect 1857 19669 1869 19672
rect 1903 19700 1915 19703
rect 1946 19700 1952 19712
rect 1903 19672 1952 19700
rect 1903 19669 1915 19672
rect 1857 19663 1915 19669
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 3326 19700 3332 19712
rect 3287 19672 3332 19700
rect 3326 19660 3332 19672
rect 3384 19660 3390 19712
rect 4430 19700 4436 19712
rect 4391 19672 4436 19700
rect 4430 19660 4436 19672
rect 4488 19660 4494 19712
rect 13354 19660 13360 19712
rect 13412 19700 13418 19712
rect 13541 19703 13599 19709
rect 13541 19700 13553 19703
rect 13412 19672 13553 19700
rect 13412 19660 13418 19672
rect 13541 19669 13553 19672
rect 13587 19669 13599 19703
rect 13998 19700 14004 19712
rect 13959 19672 14004 19700
rect 13541 19663 13599 19669
rect 13998 19660 14004 19672
rect 14056 19660 14062 19712
rect 16209 19703 16267 19709
rect 16209 19669 16221 19703
rect 16255 19700 16267 19703
rect 16390 19700 16396 19712
rect 16255 19672 16396 19700
rect 16255 19669 16267 19672
rect 16209 19663 16267 19669
rect 16390 19660 16396 19672
rect 16448 19700 16454 19712
rect 18690 19700 18696 19712
rect 16448 19672 18696 19700
rect 16448 19660 16454 19672
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 23382 19660 23388 19712
rect 23440 19700 23446 19712
rect 24719 19703 24777 19709
rect 24719 19700 24731 19703
rect 23440 19672 24731 19700
rect 23440 19660 23446 19672
rect 24719 19669 24731 19672
rect 24765 19669 24777 19703
rect 24719 19663 24777 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 2406 19496 2412 19508
rect 2367 19468 2412 19496
rect 2406 19456 2412 19468
rect 2464 19456 2470 19508
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 5224 19468 5365 19496
rect 5224 19456 5230 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 6454 19496 6460 19508
rect 6415 19468 6460 19496
rect 5353 19459 5411 19465
rect 6454 19456 6460 19468
rect 6512 19496 6518 19508
rect 8205 19499 8263 19505
rect 8205 19496 8217 19499
rect 6512 19468 8217 19496
rect 6512 19456 6518 19468
rect 8205 19465 8217 19468
rect 8251 19465 8263 19499
rect 8205 19459 8263 19465
rect 4982 19388 4988 19440
rect 5040 19428 5046 19440
rect 5721 19431 5779 19437
rect 5721 19428 5733 19431
rect 5040 19400 5733 19428
rect 5040 19388 5046 19400
rect 5721 19397 5733 19400
rect 5767 19397 5779 19431
rect 5721 19391 5779 19397
rect 6181 19431 6239 19437
rect 6181 19397 6193 19431
rect 6227 19428 6239 19431
rect 7466 19428 7472 19440
rect 6227 19400 7472 19428
rect 6227 19397 6239 19400
rect 6181 19391 6239 19397
rect 7466 19388 7472 19400
rect 7524 19388 7530 19440
rect 8220 19428 8248 19459
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10505 19499 10563 19505
rect 10505 19496 10517 19499
rect 10100 19468 10517 19496
rect 10100 19456 10106 19468
rect 10505 19465 10517 19468
rect 10551 19496 10563 19499
rect 10686 19496 10692 19508
rect 10551 19468 10692 19496
rect 10551 19465 10563 19468
rect 10505 19459 10563 19465
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 11330 19456 11336 19508
rect 11388 19496 11394 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11388 19468 11805 19496
rect 11388 19456 11394 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 11793 19459 11851 19465
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14884 19468 14933 19496
rect 14884 19456 14890 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 17126 19496 17132 19508
rect 17087 19468 17132 19496
rect 14921 19459 14979 19465
rect 17126 19456 17132 19468
rect 17184 19456 17190 19508
rect 18690 19496 18696 19508
rect 18651 19468 18696 19496
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 24670 19496 24676 19508
rect 24631 19468 24676 19496
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 12069 19431 12127 19437
rect 12069 19428 12081 19431
rect 8220 19400 12081 19428
rect 2314 19320 2320 19372
rect 2372 19360 2378 19372
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 2372 19332 3801 19360
rect 2372 19320 2378 19332
rect 3789 19329 3801 19332
rect 3835 19360 3847 19363
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 3835 19332 4721 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 6822 19320 6828 19372
rect 6880 19360 6886 19372
rect 6880 19332 6960 19360
rect 6880 19320 6886 19332
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1670 19292 1676 19304
rect 1443 19264 1676 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1670 19252 1676 19264
rect 1728 19292 1734 19304
rect 2222 19292 2228 19304
rect 1728 19264 2228 19292
rect 1728 19252 1734 19264
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 6932 19301 6960 19332
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 6917 19295 6975 19301
rect 2639 19264 3372 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 3344 19236 3372 19264
rect 6917 19261 6929 19295
rect 6963 19261 6975 19295
rect 8220 19292 8248 19400
rect 12069 19397 12081 19400
rect 12115 19428 12127 19431
rect 12161 19431 12219 19437
rect 12161 19428 12173 19431
rect 12115 19400 12173 19428
rect 12115 19397 12127 19400
rect 12069 19391 12127 19397
rect 12161 19397 12173 19400
rect 12207 19397 12219 19431
rect 12161 19391 12219 19397
rect 13446 19388 13452 19440
rect 13504 19428 13510 19440
rect 13906 19428 13912 19440
rect 13504 19400 13912 19428
rect 13504 19388 13510 19400
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19360 10839 19363
rect 11054 19360 11060 19372
rect 10827 19332 11060 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11425 19363 11483 19369
rect 11425 19329 11437 19363
rect 11471 19360 11483 19363
rect 11698 19360 11704 19372
rect 11471 19332 11704 19360
rect 11471 19329 11483 19332
rect 11425 19323 11483 19329
rect 11698 19320 11704 19332
rect 11756 19360 11762 19372
rect 12526 19360 12532 19372
rect 11756 19332 12532 19360
rect 11756 19320 11762 19332
rect 12526 19320 12532 19332
rect 12584 19320 12590 19372
rect 13998 19360 14004 19372
rect 13786 19332 14004 19360
rect 13786 19304 13814 19332
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 15620 19332 15792 19360
rect 15620 19320 15626 19332
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8220 19264 8401 19292
rect 6917 19255 6975 19261
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8846 19292 8852 19304
rect 8807 19264 8852 19292
rect 8389 19255 8447 19261
rect 8846 19252 8852 19264
rect 8904 19292 8910 19304
rect 9401 19295 9459 19301
rect 9401 19292 9413 19295
rect 8904 19264 9413 19292
rect 8904 19252 8910 19264
rect 9401 19261 9413 19264
rect 9447 19261 9459 19295
rect 9401 19255 9459 19261
rect 12069 19295 12127 19301
rect 12069 19261 12081 19295
rect 12115 19292 12127 19295
rect 12342 19292 12348 19304
rect 12115 19264 12348 19292
rect 12115 19261 12127 19264
rect 12069 19255 12127 19261
rect 12342 19252 12348 19264
rect 12400 19292 12406 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12400 19264 12449 19292
rect 12400 19252 12406 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 2133 19227 2191 19233
rect 2133 19193 2145 19227
rect 2179 19224 2191 19227
rect 2498 19224 2504 19236
rect 2179 19196 2504 19224
rect 2179 19193 2191 19196
rect 2133 19187 2191 19193
rect 2498 19184 2504 19196
rect 2556 19224 2562 19236
rect 2955 19227 3013 19233
rect 2556 19196 2855 19224
rect 2556 19184 2562 19196
rect 2827 19156 2855 19196
rect 2955 19193 2967 19227
rect 3001 19224 3013 19227
rect 3050 19224 3056 19236
rect 3001 19196 3056 19224
rect 3001 19193 3013 19196
rect 2955 19187 3013 19193
rect 3050 19184 3056 19196
rect 3108 19184 3114 19236
rect 3326 19184 3332 19236
rect 3384 19224 3390 19236
rect 4246 19224 4252 19236
rect 3384 19196 4252 19224
rect 3384 19184 3390 19196
rect 4246 19184 4252 19196
rect 4304 19184 4310 19236
rect 4430 19224 4436 19236
rect 4391 19196 4436 19224
rect 4430 19184 4436 19196
rect 4488 19184 4494 19236
rect 4525 19227 4583 19233
rect 4525 19193 4537 19227
rect 4571 19193 4583 19227
rect 4525 19187 4583 19193
rect 3510 19156 3516 19168
rect 2827 19128 3516 19156
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4540 19156 4568 19187
rect 4798 19184 4804 19236
rect 4856 19224 4862 19236
rect 6825 19227 6883 19233
rect 6825 19224 6837 19227
rect 4856 19196 6837 19224
rect 4856 19184 4862 19196
rect 6825 19193 6837 19196
rect 6871 19193 6883 19227
rect 6825 19187 6883 19193
rect 10137 19227 10195 19233
rect 10137 19193 10149 19227
rect 10183 19224 10195 19227
rect 10873 19227 10931 19233
rect 10183 19196 10640 19224
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 7926 19156 7932 19168
rect 4212 19128 4568 19156
rect 7887 19128 7932 19156
rect 4212 19116 4218 19128
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8478 19156 8484 19168
rect 8439 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 10612 19156 10640 19196
rect 10873 19193 10885 19227
rect 10919 19224 10931 19227
rect 10962 19224 10968 19236
rect 10919 19196 10968 19224
rect 10919 19193 10931 19196
rect 10873 19187 10931 19193
rect 10888 19156 10916 19187
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 12526 19184 12532 19236
rect 12584 19224 12590 19236
rect 12912 19224 12940 19255
rect 13722 19252 13728 19304
rect 13780 19264 13814 19304
rect 15764 19301 15792 19332
rect 15749 19295 15807 19301
rect 13924 19264 15700 19292
rect 13780 19252 13786 19264
rect 13170 19224 13176 19236
rect 12584 19196 12940 19224
rect 13131 19196 13176 19224
rect 12584 19184 12590 19196
rect 13170 19184 13176 19196
rect 13228 19184 13234 19236
rect 13924 19224 13952 19264
rect 14363 19227 14421 19233
rect 14363 19224 14375 19227
rect 13786 19196 13952 19224
rect 14016 19196 14375 19224
rect 10612 19128 10916 19156
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13786 19156 13814 19196
rect 13044 19128 13814 19156
rect 13044 19116 13050 19128
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 14016 19156 14044 19196
rect 14363 19193 14375 19196
rect 14409 19224 14421 19227
rect 15289 19227 15347 19233
rect 15289 19224 15301 19227
rect 14409 19196 15301 19224
rect 14409 19193 14421 19196
rect 14363 19187 14421 19193
rect 15289 19193 15301 19196
rect 15335 19224 15347 19227
rect 15378 19224 15384 19236
rect 15335 19196 15384 19224
rect 15335 19193 15347 19196
rect 15289 19187 15347 19193
rect 15378 19184 15384 19196
rect 15436 19184 15442 19236
rect 15562 19224 15568 19236
rect 15523 19196 15568 19224
rect 15562 19184 15568 19196
rect 15620 19184 15626 19236
rect 15672 19156 15700 19264
rect 15749 19261 15761 19295
rect 15795 19261 15807 19295
rect 16298 19292 16304 19304
rect 16259 19264 16304 19292
rect 15749 19255 15807 19261
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 13964 19128 14057 19156
rect 15672 19128 15853 19156
rect 13964 19116 13970 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 17494 19156 17500 19168
rect 17455 19128 17500 19156
rect 15841 19119 15899 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 4341 18955 4399 18961
rect 4341 18952 4353 18955
rect 2148 18924 4353 18952
rect 2038 18844 2044 18896
rect 2096 18884 2102 18896
rect 2148 18893 2176 18924
rect 4341 18921 4353 18924
rect 4387 18921 4399 18955
rect 8021 18955 8079 18961
rect 8021 18952 8033 18955
rect 4341 18915 4399 18921
rect 5229 18924 8033 18952
rect 2133 18887 2191 18893
rect 2133 18884 2145 18887
rect 2096 18856 2145 18884
rect 2096 18844 2102 18856
rect 2133 18853 2145 18856
rect 2179 18853 2191 18887
rect 2133 18847 2191 18853
rect 2222 18844 2228 18896
rect 2280 18884 2286 18896
rect 3329 18887 3387 18893
rect 3329 18884 3341 18887
rect 2280 18856 3341 18884
rect 2280 18844 2286 18856
rect 3329 18853 3341 18856
rect 3375 18853 3387 18887
rect 3329 18847 3387 18853
rect 4246 18844 4252 18896
rect 4304 18884 4310 18896
rect 5229 18884 5257 18924
rect 8021 18921 8033 18924
rect 8067 18921 8079 18955
rect 11054 18952 11060 18964
rect 11015 18924 11060 18952
rect 8021 18915 8079 18921
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 12805 18955 12863 18961
rect 12805 18952 12817 18955
rect 12308 18924 12817 18952
rect 12308 18912 12314 18924
rect 12805 18921 12817 18924
rect 12851 18921 12863 18955
rect 12805 18915 12863 18921
rect 13170 18912 13176 18964
rect 13228 18952 13234 18964
rect 15105 18955 15163 18961
rect 15105 18952 15117 18955
rect 13228 18924 15117 18952
rect 13228 18912 13234 18924
rect 15105 18921 15117 18924
rect 15151 18952 15163 18955
rect 15286 18952 15292 18964
rect 15151 18924 15292 18952
rect 15151 18921 15163 18924
rect 15105 18915 15163 18921
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 16114 18952 16120 18964
rect 15580 18924 16120 18952
rect 6546 18884 6552 18896
rect 4304 18856 5257 18884
rect 6507 18856 6552 18884
rect 4304 18844 4310 18856
rect 6546 18844 6552 18856
rect 6604 18844 6610 18896
rect 6822 18844 6828 18896
rect 6880 18884 6886 18896
rect 7377 18887 7435 18893
rect 7377 18884 7389 18887
rect 6880 18856 7389 18884
rect 6880 18844 6886 18856
rect 7377 18853 7389 18856
rect 7423 18853 7435 18887
rect 7377 18847 7435 18853
rect 12526 18844 12532 18896
rect 12584 18884 12590 18896
rect 13722 18884 13728 18896
rect 12584 18856 13492 18884
rect 13683 18856 13728 18884
rect 12584 18844 12590 18856
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 7926 18816 7932 18828
rect 4212 18788 4257 18816
rect 7887 18788 7932 18816
rect 4212 18776 4218 18788
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 8018 18776 8024 18828
rect 8076 18816 8082 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 8076 18788 8401 18816
rect 8076 18776 8082 18788
rect 8389 18785 8401 18788
rect 8435 18785 8447 18819
rect 10226 18816 10232 18828
rect 10187 18788 10232 18816
rect 8389 18779 8447 18785
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 11698 18816 11704 18828
rect 11655 18788 11704 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13464 18825 13492 18856
rect 13722 18844 13728 18856
rect 13780 18844 13786 18896
rect 15580 18893 15608 18924
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 15565 18887 15623 18893
rect 15565 18853 15577 18887
rect 15611 18853 15623 18887
rect 15565 18847 15623 18853
rect 15930 18844 15936 18896
rect 15988 18884 15994 18896
rect 16945 18887 17003 18893
rect 16945 18884 16957 18887
rect 15988 18856 16957 18884
rect 15988 18844 15994 18856
rect 16945 18853 16957 18856
rect 16991 18853 17003 18887
rect 16945 18847 17003 18853
rect 12989 18819 13047 18825
rect 12989 18816 13001 18819
rect 12768 18788 13001 18816
rect 12768 18776 12774 18788
rect 12989 18785 13001 18788
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18785 13507 18819
rect 13449 18779 13507 18785
rect 1854 18708 1860 18760
rect 1912 18748 1918 18760
rect 2041 18751 2099 18757
rect 2041 18748 2053 18751
rect 1912 18720 2053 18748
rect 1912 18708 1918 18720
rect 2041 18717 2053 18720
rect 2087 18717 2099 18751
rect 2314 18748 2320 18760
rect 2275 18720 2320 18748
rect 2041 18711 2099 18717
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 5169 18751 5227 18757
rect 5169 18748 5181 18751
rect 3476 18720 5181 18748
rect 3476 18708 3482 18720
rect 5169 18717 5181 18720
rect 5215 18748 5227 18751
rect 5258 18748 5264 18760
rect 5215 18720 5264 18748
rect 5215 18717 5227 18720
rect 5169 18711 5227 18717
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18717 6515 18751
rect 7098 18748 7104 18760
rect 7059 18720 7104 18748
rect 6457 18711 6515 18717
rect 1670 18680 1676 18692
rect 1583 18652 1676 18680
rect 1670 18640 1676 18652
rect 1728 18680 1734 18692
rect 2590 18680 2596 18692
rect 1728 18652 2596 18680
rect 1728 18640 1734 18652
rect 2590 18640 2596 18652
rect 2648 18640 2654 18692
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 5994 18572 6000 18624
rect 6052 18612 6058 18624
rect 6181 18615 6239 18621
rect 6181 18612 6193 18615
rect 6052 18584 6193 18612
rect 6052 18572 6058 18584
rect 6181 18581 6193 18584
rect 6227 18612 6239 18615
rect 6472 18612 6500 18711
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 15470 18748 15476 18760
rect 15383 18720 15476 18748
rect 15470 18708 15476 18720
rect 15528 18748 15534 18760
rect 15746 18748 15752 18760
rect 15528 18720 15752 18748
rect 15528 18708 15534 18720
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16206 18748 16212 18760
rect 16163 18720 16212 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 9858 18640 9864 18692
rect 9916 18680 9922 18692
rect 11747 18683 11805 18689
rect 11747 18680 11759 18683
rect 9916 18652 11759 18680
rect 9916 18640 9922 18652
rect 11747 18649 11759 18652
rect 11793 18649 11805 18683
rect 11747 18643 11805 18649
rect 6227 18584 6500 18612
rect 6227 18581 6239 18584
rect 6181 18575 6239 18581
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10321 18615 10379 18621
rect 10321 18612 10333 18615
rect 10192 18584 10333 18612
rect 10192 18572 10198 18584
rect 10321 18581 10333 18584
rect 10367 18581 10379 18615
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 10321 18575 10379 18581
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 14090 18612 14096 18624
rect 14051 18584 14096 18612
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14826 18572 14832 18624
rect 14884 18612 14890 18624
rect 16298 18612 16304 18624
rect 14884 18584 16304 18612
rect 14884 18572 14890 18584
rect 16298 18572 16304 18584
rect 16356 18612 16362 18624
rect 16393 18615 16451 18621
rect 16393 18612 16405 18615
rect 16356 18584 16405 18612
rect 16356 18572 16362 18584
rect 16393 18581 16405 18584
rect 16439 18581 16451 18615
rect 16393 18575 16451 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2038 18408 2044 18420
rect 1999 18380 2044 18408
rect 2038 18368 2044 18380
rect 2096 18368 2102 18420
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 4154 18408 4160 18420
rect 4120 18380 4160 18408
rect 4120 18368 4126 18380
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 6086 18368 6092 18420
rect 6144 18408 6150 18420
rect 7926 18408 7932 18420
rect 6144 18380 7932 18408
rect 6144 18368 6150 18380
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 11698 18408 11704 18420
rect 11659 18380 11704 18408
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 1627 18343 1685 18349
rect 1627 18309 1639 18343
rect 1673 18340 1685 18343
rect 3694 18340 3700 18352
rect 1673 18312 3700 18340
rect 1673 18309 1685 18312
rect 1627 18303 1685 18309
rect 3694 18300 3700 18312
rect 3752 18300 3758 18352
rect 7098 18300 7104 18352
rect 7156 18340 7162 18352
rect 7469 18343 7527 18349
rect 7469 18340 7481 18343
rect 7156 18312 7481 18340
rect 7156 18300 7162 18312
rect 7469 18309 7481 18312
rect 7515 18309 7527 18343
rect 7944 18340 7972 18368
rect 9674 18340 9680 18352
rect 7944 18312 9680 18340
rect 7469 18303 7527 18309
rect 9674 18300 9680 18312
rect 9732 18340 9738 18352
rect 12161 18343 12219 18349
rect 12161 18340 12173 18343
rect 9732 18312 12173 18340
rect 9732 18300 9738 18312
rect 12161 18309 12173 18312
rect 12207 18309 12219 18343
rect 12161 18303 12219 18309
rect 15013 18343 15071 18349
rect 15013 18309 15025 18343
rect 15059 18340 15071 18343
rect 16114 18340 16120 18352
rect 15059 18312 16120 18340
rect 15059 18309 15071 18312
rect 15013 18303 15071 18309
rect 5258 18272 5264 18284
rect 5219 18244 5264 18272
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 6273 18275 6331 18281
rect 6273 18241 6285 18275
rect 6319 18272 6331 18275
rect 6917 18275 6975 18281
rect 6917 18272 6929 18275
rect 6319 18244 6929 18272
rect 6319 18241 6331 18244
rect 6273 18235 6331 18241
rect 6917 18241 6929 18244
rect 6963 18272 6975 18275
rect 8386 18272 8392 18284
rect 6963 18244 8392 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 9640 18244 10149 18272
rect 9640 18232 9646 18244
rect 10137 18241 10149 18244
rect 10183 18272 10195 18275
rect 10870 18272 10876 18284
rect 10183 18244 10876 18272
rect 10183 18241 10195 18244
rect 10137 18235 10195 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 1556 18207 1614 18213
rect 1556 18173 1568 18207
rect 1602 18204 1614 18207
rect 1670 18204 1676 18216
rect 1602 18176 1676 18204
rect 1602 18173 1614 18176
rect 1556 18167 1614 18173
rect 1670 18164 1676 18176
rect 1728 18164 1734 18216
rect 2777 18207 2835 18213
rect 2777 18173 2789 18207
rect 2823 18204 2835 18207
rect 2958 18204 2964 18216
rect 2823 18176 2964 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 2958 18164 2964 18176
rect 3016 18204 3022 18216
rect 4798 18204 4804 18216
rect 3016 18176 4804 18204
rect 3016 18164 3022 18176
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 7650 18164 7656 18216
rect 7708 18204 7714 18216
rect 9033 18207 9091 18213
rect 9033 18204 9045 18207
rect 7708 18176 9045 18204
rect 7708 18164 7714 18176
rect 9033 18173 9045 18176
rect 9079 18204 9091 18207
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 9079 18176 9413 18204
rect 9079 18173 9091 18176
rect 9033 18167 9091 18173
rect 9401 18173 9413 18176
rect 9447 18173 9459 18207
rect 12176 18204 12204 18303
rect 16114 18300 16120 18312
rect 16172 18300 16178 18352
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18272 13323 18275
rect 14090 18272 14096 18284
rect 13311 18244 14096 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 14090 18232 14096 18244
rect 14148 18232 14154 18284
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18272 15439 18275
rect 15930 18272 15936 18284
rect 15427 18244 15936 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16206 18272 16212 18284
rect 16167 18244 16212 18272
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 12529 18207 12587 18213
rect 12529 18204 12541 18207
rect 12176 18176 12541 18204
rect 9401 18167 9459 18173
rect 12529 18173 12541 18176
rect 12575 18204 12587 18207
rect 12710 18204 12716 18216
rect 12575 18176 12716 18204
rect 12575 18173 12587 18176
rect 12529 18167 12587 18173
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 12986 18204 12992 18216
rect 12947 18176 12992 18204
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 5258 18136 5264 18148
rect 3160 18108 5264 18136
rect 2685 18071 2743 18077
rect 2685 18037 2697 18071
rect 2731 18068 2743 18071
rect 3050 18068 3056 18080
rect 2731 18040 3056 18068
rect 2731 18037 2743 18040
rect 2685 18031 2743 18037
rect 3050 18028 3056 18040
rect 3108 18068 3114 18080
rect 3160 18077 3188 18108
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 5353 18139 5411 18145
rect 5353 18105 5365 18139
rect 5399 18105 5411 18139
rect 5353 18099 5411 18105
rect 5905 18139 5963 18145
rect 5905 18105 5917 18139
rect 5951 18136 5963 18139
rect 5994 18136 6000 18148
rect 5951 18108 6000 18136
rect 5951 18105 5963 18108
rect 5905 18099 5963 18105
rect 3145 18071 3203 18077
rect 3145 18068 3157 18071
rect 3108 18040 3157 18068
rect 3108 18028 3114 18040
rect 3145 18037 3157 18040
rect 3191 18037 3203 18071
rect 3145 18031 3203 18037
rect 3697 18071 3755 18077
rect 3697 18037 3709 18071
rect 3743 18068 3755 18071
rect 4062 18068 4068 18080
rect 3743 18040 4068 18068
rect 3743 18037 3755 18040
rect 3697 18031 3755 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 5077 18071 5135 18077
rect 5077 18037 5089 18071
rect 5123 18068 5135 18071
rect 5368 18068 5396 18099
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 8389 18139 8447 18145
rect 8389 18136 8401 18139
rect 7055 18108 8401 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 8389 18105 8401 18108
rect 8435 18105 8447 18139
rect 8389 18099 8447 18105
rect 6362 18068 6368 18080
rect 5123 18040 6368 18068
rect 5123 18037 5135 18040
rect 5077 18031 5135 18037
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 6641 18071 6699 18077
rect 6641 18037 6653 18071
rect 6687 18068 6699 18071
rect 7024 18068 7052 18099
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 10778 18136 10784 18148
rect 10284 18108 10377 18136
rect 10739 18108 10784 18136
rect 10284 18096 10290 18108
rect 10778 18096 10784 18108
rect 10836 18096 10842 18148
rect 13446 18096 13452 18148
rect 13504 18136 13510 18148
rect 14414 18139 14472 18145
rect 14414 18136 14426 18139
rect 13504 18108 14426 18136
rect 13504 18096 13510 18108
rect 6687 18040 7052 18068
rect 9953 18071 10011 18077
rect 6687 18037 6699 18040
rect 6641 18031 6699 18037
rect 9953 18037 9965 18071
rect 9999 18068 10011 18071
rect 10244 18068 10272 18096
rect 11054 18068 11060 18080
rect 9999 18040 11060 18068
rect 9999 18037 10011 18040
rect 9953 18031 10011 18037
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13541 18071 13599 18077
rect 13541 18068 13553 18071
rect 12768 18040 13553 18068
rect 12768 18028 12774 18040
rect 13541 18037 13553 18040
rect 13587 18068 13599 18071
rect 13814 18068 13820 18080
rect 13587 18040 13820 18068
rect 13587 18037 13599 18040
rect 13541 18031 13599 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14016 18077 14044 18108
rect 14414 18105 14426 18108
rect 14460 18105 14472 18139
rect 14414 18099 14472 18105
rect 16025 18139 16083 18145
rect 16025 18105 16037 18139
rect 16071 18105 16083 18139
rect 16025 18099 16083 18105
rect 14001 18071 14059 18077
rect 14001 18037 14013 18071
rect 14047 18037 14059 18071
rect 15746 18068 15752 18080
rect 15707 18040 15752 18068
rect 14001 18031 14059 18037
rect 15746 18028 15752 18040
rect 15804 18068 15810 18080
rect 16040 18068 16068 18099
rect 15804 18040 16068 18068
rect 15804 18028 15810 18040
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 16172 18040 16865 18068
rect 16172 18028 16178 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1394 17864 1400 17876
rect 1355 17836 1400 17864
rect 1394 17824 1400 17836
rect 1452 17824 1458 17876
rect 6457 17867 6515 17873
rect 6457 17833 6469 17867
rect 6503 17864 6515 17867
rect 6546 17864 6552 17876
rect 6503 17836 6552 17864
rect 6503 17833 6515 17836
rect 6457 17827 6515 17833
rect 6546 17824 6552 17836
rect 6604 17864 6610 17876
rect 7561 17867 7619 17873
rect 7561 17864 7573 17867
rect 6604 17836 7573 17864
rect 6604 17824 6610 17836
rect 7561 17833 7573 17836
rect 7607 17864 7619 17867
rect 7650 17864 7656 17876
rect 7607 17836 7656 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 8018 17864 8024 17876
rect 7979 17836 8024 17864
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 8386 17864 8392 17876
rect 8347 17836 8392 17864
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 10042 17864 10048 17876
rect 10003 17836 10048 17864
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 10597 17867 10655 17873
rect 10597 17833 10609 17867
rect 10643 17864 10655 17867
rect 11054 17864 11060 17876
rect 10643 17836 11060 17864
rect 10643 17833 10655 17836
rect 10597 17827 10655 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 13354 17864 13360 17876
rect 13315 17836 13360 17864
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 15105 17867 15163 17873
rect 15105 17833 15117 17867
rect 15151 17864 15163 17867
rect 15470 17864 15476 17876
rect 15151 17836 15476 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 15746 17864 15752 17876
rect 15707 17836 15752 17864
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 2222 17756 2228 17808
rect 2280 17796 2286 17808
rect 2593 17799 2651 17805
rect 2593 17796 2605 17799
rect 2280 17768 2605 17796
rect 2280 17756 2286 17768
rect 2593 17765 2605 17768
rect 2639 17765 2651 17799
rect 2593 17759 2651 17765
rect 5255 17799 5313 17805
rect 5255 17765 5267 17799
rect 5301 17796 5313 17799
rect 5350 17796 5356 17808
rect 5301 17768 5356 17796
rect 5301 17765 5313 17768
rect 5255 17759 5313 17765
rect 5350 17756 5356 17768
rect 5408 17796 5414 17808
rect 6638 17796 6644 17808
rect 5408 17768 6644 17796
rect 5408 17756 5414 17768
rect 6638 17756 6644 17768
rect 6696 17796 6702 17808
rect 7003 17799 7061 17805
rect 7003 17796 7015 17799
rect 6696 17768 7015 17796
rect 6696 17756 6702 17768
rect 7003 17765 7015 17768
rect 7049 17796 7061 17799
rect 10060 17796 10088 17824
rect 10870 17796 10876 17808
rect 7049 17768 10088 17796
rect 10831 17768 10876 17796
rect 7049 17765 7061 17768
rect 7003 17759 7061 17765
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 12253 17799 12311 17805
rect 12253 17765 12265 17799
rect 12299 17796 12311 17799
rect 12526 17796 12532 17808
rect 12299 17768 12532 17796
rect 12299 17765 12311 17768
rect 12253 17759 12311 17765
rect 12526 17756 12532 17768
rect 12584 17796 12590 17808
rect 12897 17799 12955 17805
rect 12897 17796 12909 17799
rect 12584 17768 12909 17796
rect 12584 17756 12590 17768
rect 12897 17765 12909 17768
rect 12943 17765 12955 17799
rect 12897 17759 12955 17765
rect 12986 17756 12992 17808
rect 13044 17796 13050 17808
rect 13044 17768 13584 17796
rect 13044 17756 13050 17768
rect 8938 17728 8944 17740
rect 4126 17700 8944 17728
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 2501 17663 2559 17669
rect 2501 17660 2513 17663
rect 2363 17632 2513 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 2501 17629 2513 17632
rect 2547 17660 2559 17663
rect 4126 17660 4154 17700
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 11238 17688 11244 17740
rect 11296 17728 11302 17740
rect 11517 17731 11575 17737
rect 11517 17728 11529 17731
rect 11296 17700 11529 17728
rect 11296 17688 11302 17700
rect 11517 17697 11529 17700
rect 11563 17697 11575 17731
rect 11517 17691 11575 17697
rect 12342 17688 12348 17740
rect 12400 17728 12406 17740
rect 13556 17737 13584 17768
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 13872 17768 16896 17796
rect 13872 17756 13878 17768
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12400 17700 13093 17728
rect 12400 17688 12406 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 16114 17728 16120 17740
rect 15979 17700 16120 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 2547 17632 4154 17660
rect 4893 17663 4951 17669
rect 2547 17629 2559 17632
rect 2501 17623 2559 17629
rect 4893 17629 4905 17663
rect 4939 17660 4951 17663
rect 5166 17660 5172 17672
rect 4939 17632 5172 17660
rect 4939 17629 4951 17632
rect 4893 17623 4951 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 6236 17632 6653 17660
rect 6236 17620 6242 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 11882 17660 11888 17672
rect 11843 17632 11888 17660
rect 9677 17623 9735 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 3053 17595 3111 17601
rect 3053 17592 3065 17595
rect 2740 17564 3065 17592
rect 2740 17552 2746 17564
rect 3053 17561 3065 17564
rect 3099 17561 3111 17595
rect 3053 17555 3111 17561
rect 5813 17595 5871 17601
rect 5813 17561 5825 17595
rect 5859 17592 5871 17595
rect 7006 17592 7012 17604
rect 5859 17564 7012 17592
rect 5859 17561 5871 17564
rect 5813 17555 5871 17561
rect 7006 17552 7012 17564
rect 7064 17552 7070 17604
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 9692 17592 9720 17623
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 13556 17660 13584 17691
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 16868 17737 16896 17768
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17218 17728 17224 17740
rect 16899 17700 17224 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 17586 17728 17592 17740
rect 17359 17700 17592 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 13906 17660 13912 17672
rect 13556 17632 13912 17660
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 14016 17632 17417 17660
rect 14016 17592 14044 17632
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 9548 17564 14044 17592
rect 9548 17552 9554 17564
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 1854 17524 1860 17536
rect 1452 17496 1860 17524
rect 1452 17484 1458 17496
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4522 17524 4528 17536
rect 4387 17496 4528 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4522 17484 4528 17496
rect 4580 17484 4586 17536
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 8849 17527 8907 17533
rect 8849 17524 8861 17527
rect 8628 17496 8861 17524
rect 8628 17484 8634 17496
rect 8849 17493 8861 17496
rect 8895 17493 8907 17527
rect 11330 17524 11336 17536
rect 11291 17496 11336 17524
rect 8849 17487 8907 17493
rect 11330 17484 11336 17496
rect 11388 17524 11394 17536
rect 11655 17527 11713 17533
rect 11655 17524 11667 17527
rect 11388 17496 11667 17524
rect 11388 17484 11394 17496
rect 11655 17493 11667 17496
rect 11701 17493 11713 17527
rect 11790 17524 11796 17536
rect 11751 17496 11796 17524
rect 11655 17487 11713 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 12158 17484 12164 17536
rect 12216 17524 12222 17536
rect 12529 17527 12587 17533
rect 12529 17524 12541 17527
rect 12216 17496 12541 17524
rect 12216 17484 12222 17496
rect 12529 17493 12541 17496
rect 12575 17524 12587 17527
rect 12986 17524 12992 17536
rect 12575 17496 12992 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 14090 17524 14096 17536
rect 14051 17496 14096 17524
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 8018 17320 8024 17332
rect 5408 17292 8024 17320
rect 5408 17280 5414 17292
rect 8018 17280 8024 17292
rect 8076 17320 8082 17332
rect 8849 17323 8907 17329
rect 8849 17320 8861 17323
rect 8076 17292 8861 17320
rect 8076 17280 8082 17292
rect 8849 17289 8861 17292
rect 8895 17289 8907 17323
rect 10134 17320 10140 17332
rect 10095 17292 10140 17320
rect 8849 17283 8907 17289
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 12342 17280 12348 17332
rect 12400 17320 12406 17332
rect 13081 17323 13139 17329
rect 13081 17320 13093 17323
rect 12400 17292 13093 17320
rect 12400 17280 12406 17292
rect 13081 17289 13093 17292
rect 13127 17289 13139 17323
rect 13081 17283 13139 17289
rect 13906 17280 13912 17332
rect 13964 17320 13970 17332
rect 14645 17323 14703 17329
rect 14645 17320 14657 17323
rect 13964 17292 14657 17320
rect 13964 17280 13970 17292
rect 14645 17289 14657 17292
rect 14691 17289 14703 17323
rect 14645 17283 14703 17289
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16577 17323 16635 17329
rect 16577 17320 16589 17323
rect 16264 17292 16589 17320
rect 16264 17280 16270 17292
rect 16577 17289 16589 17292
rect 16623 17289 16635 17323
rect 17218 17320 17224 17332
rect 17179 17292 17224 17320
rect 16577 17283 16635 17289
rect 5721 17255 5779 17261
rect 5721 17221 5733 17255
rect 5767 17252 5779 17255
rect 6638 17252 6644 17264
rect 5767 17224 6644 17252
rect 5767 17221 5779 17224
rect 5721 17215 5779 17221
rect 6638 17212 6644 17224
rect 6696 17212 6702 17264
rect 8386 17212 8392 17264
rect 8444 17252 8450 17264
rect 8527 17255 8585 17261
rect 8527 17252 8539 17255
rect 8444 17224 8539 17252
rect 8444 17212 8450 17224
rect 8527 17221 8539 17224
rect 8573 17221 8585 17255
rect 8527 17215 8585 17221
rect 8665 17255 8723 17261
rect 8665 17221 8677 17255
rect 8711 17252 8723 17255
rect 9214 17252 9220 17264
rect 8711 17224 9220 17252
rect 8711 17221 8723 17224
rect 8665 17215 8723 17221
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 2498 17184 2504 17196
rect 1903 17156 2504 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 2682 17184 2688 17196
rect 2643 17156 2688 17184
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4614 17184 4620 17196
rect 4203 17156 4620 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 4614 17144 4620 17156
rect 4672 17184 4678 17196
rect 4672 17156 5396 17184
rect 4672 17144 4678 17156
rect 4522 17116 4528 17128
rect 4483 17088 4528 17116
rect 4522 17076 4528 17088
rect 4580 17076 4586 17128
rect 5092 17125 5120 17156
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 5261 17119 5319 17125
rect 5261 17085 5273 17119
rect 5307 17085 5319 17119
rect 5368 17116 5396 17156
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6052 17156 7205 17184
rect 6052 17144 6058 17156
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17184 7987 17187
rect 8680 17184 8708 17215
rect 9214 17212 9220 17224
rect 9272 17252 9278 17264
rect 11790 17252 11796 17264
rect 9272 17224 11796 17252
rect 9272 17212 9278 17224
rect 11790 17212 11796 17224
rect 11848 17252 11854 17264
rect 11885 17255 11943 17261
rect 11885 17252 11897 17255
rect 11848 17224 11897 17252
rect 11848 17212 11854 17224
rect 11885 17221 11897 17224
rect 11931 17221 11943 17255
rect 11885 17215 11943 17221
rect 7975 17156 8708 17184
rect 8757 17187 8815 17193
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 9306 17184 9312 17196
rect 8803 17156 9312 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 6454 17116 6460 17128
rect 5368 17088 6460 17116
rect 5261 17079 5319 17085
rect 2130 17008 2136 17060
rect 2188 17048 2194 17060
rect 2409 17051 2467 17057
rect 2409 17048 2421 17051
rect 2188 17020 2421 17048
rect 2188 17008 2194 17020
rect 2409 17017 2421 17020
rect 2455 17017 2467 17051
rect 2409 17011 2467 17017
rect 2222 16980 2228 16992
rect 2183 16952 2228 16980
rect 2222 16940 2228 16952
rect 2280 16940 2286 16992
rect 2424 16980 2452 17011
rect 2498 17008 2504 17060
rect 2556 17048 2562 17060
rect 2556 17020 2601 17048
rect 2556 17008 2562 17020
rect 3510 17008 3516 17060
rect 3568 17048 3574 17060
rect 3789 17051 3847 17057
rect 3789 17048 3801 17051
rect 3568 17020 3801 17048
rect 3568 17008 3574 17020
rect 3789 17017 3801 17020
rect 3835 17048 3847 17051
rect 5276 17048 5304 17079
rect 6454 17076 6460 17088
rect 6512 17076 6518 17128
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 8772 17116 8800 17147
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 9769 17187 9827 17193
rect 9769 17153 9781 17187
rect 9815 17184 9827 17187
rect 10042 17184 10048 17196
rect 9815 17156 10048 17184
rect 9815 17153 9827 17156
rect 9769 17147 9827 17153
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 10686 17184 10692 17196
rect 10459 17156 10692 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 16172 17156 16221 17184
rect 16172 17144 16178 17156
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 13446 17116 13452 17128
rect 8343 17088 8800 17116
rect 13407 17088 13452 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 13446 17076 13452 17088
rect 13504 17116 13510 17128
rect 14090 17116 14096 17128
rect 13504 17088 14096 17116
rect 13504 17076 13510 17088
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 15105 17119 15163 17125
rect 15105 17116 15117 17119
rect 14415 17088 15117 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 15105 17085 15117 17088
rect 15151 17116 15163 17119
rect 15746 17116 15752 17128
rect 15151 17088 15752 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15746 17076 15752 17088
rect 15804 17076 15810 17128
rect 16592 17116 16620 17283
rect 17218 17280 17224 17292
rect 17276 17280 17282 17332
rect 24762 17252 24768 17264
rect 24723 17224 24768 17252
rect 24762 17212 24768 17224
rect 24820 17212 24826 17264
rect 24486 17184 24492 17196
rect 24447 17156 24492 17184
rect 24486 17144 24492 17156
rect 24544 17184 24550 17196
rect 25133 17187 25191 17193
rect 25133 17184 25145 17187
rect 24544 17156 25145 17184
rect 24544 17144 24550 17156
rect 25133 17153 25145 17156
rect 25179 17153 25191 17187
rect 25133 17147 25191 17153
rect 16796 17119 16854 17125
rect 16796 17116 16808 17119
rect 16592 17088 16808 17116
rect 16796 17085 16808 17088
rect 16842 17085 16854 17119
rect 16796 17079 16854 17085
rect 16899 17119 16957 17125
rect 16899 17085 16911 17119
rect 16945 17116 16957 17119
rect 17218 17116 17224 17128
rect 16945 17088 17224 17116
rect 16945 17085 16957 17088
rect 16899 17079 16957 17085
rect 17218 17076 17224 17088
rect 17276 17076 17282 17128
rect 5534 17048 5540 17060
rect 3835 17020 5540 17048
rect 3835 17017 3847 17020
rect 3789 17011 3847 17017
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 6917 17051 6975 17057
rect 6917 17017 6929 17051
rect 6963 17017 6975 17051
rect 6917 17011 6975 17017
rect 3329 16983 3387 16989
rect 3329 16980 3341 16983
rect 2424 16952 3341 16980
rect 3329 16949 3341 16952
rect 3375 16949 3387 16983
rect 5166 16980 5172 16992
rect 5127 16952 5172 16980
rect 3329 16943 3387 16949
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 6178 16980 6184 16992
rect 6139 16952 6184 16980
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6932 16980 6960 17011
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 8389 17051 8447 17057
rect 7064 17020 7109 17048
rect 7064 17008 7070 17020
rect 8389 17017 8401 17051
rect 8435 17048 8447 17051
rect 8570 17048 8576 17060
rect 8435 17020 8576 17048
rect 8435 17017 8447 17020
rect 8389 17011 8447 17017
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17017 10563 17051
rect 10505 17011 10563 17017
rect 7558 16980 7564 16992
rect 6932 16952 7564 16980
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10520 16980 10548 17011
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 11057 17051 11115 17057
rect 11057 17048 11069 17051
rect 10836 17020 11069 17048
rect 10836 17008 10842 17020
rect 11057 17017 11069 17020
rect 11103 17048 11115 17051
rect 12066 17048 12072 17060
rect 11103 17020 12072 17048
rect 11103 17017 11115 17020
rect 11057 17011 11115 17017
rect 12066 17008 12072 17020
rect 12124 17008 12130 17060
rect 13811 17051 13869 17057
rect 13811 17017 13823 17051
rect 13857 17048 13869 17051
rect 13998 17048 14004 17060
rect 13857 17020 14004 17048
rect 13857 17017 13869 17020
rect 13811 17011 13869 17017
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 10192 16952 10548 16980
rect 10192 16940 10198 16952
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 11204 16952 11529 16980
rect 11204 16940 11210 16952
rect 11517 16949 11529 16952
rect 11563 16949 11575 16983
rect 12434 16980 12440 16992
rect 12395 16952 12440 16980
rect 11517 16943 11575 16949
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 15470 16980 15476 16992
rect 15431 16952 15476 16980
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 17586 16980 17592 16992
rect 17547 16952 17592 16980
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 4338 16776 4344 16788
rect 4299 16748 4344 16776
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 5166 16776 5172 16788
rect 5127 16748 5172 16776
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 6178 16776 6184 16788
rect 6139 16748 6184 16776
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 6917 16779 6975 16785
rect 6917 16745 6929 16779
rect 6963 16776 6975 16779
rect 7006 16776 7012 16788
rect 6963 16748 7012 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 9490 16776 9496 16788
rect 9451 16748 9496 16776
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10744 16748 10977 16776
rect 10744 16736 10750 16748
rect 10965 16745 10977 16748
rect 11011 16776 11023 16779
rect 12434 16776 12440 16788
rect 11011 16748 12440 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 13265 16779 13323 16785
rect 13265 16745 13277 16779
rect 13311 16776 13323 16779
rect 13446 16776 13452 16788
rect 13311 16748 13452 16776
rect 13311 16745 13323 16748
rect 13265 16739 13323 16745
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 13998 16776 14004 16788
rect 13959 16748 14004 16776
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 16022 16776 16028 16788
rect 15396 16748 16028 16776
rect 2406 16668 2412 16720
rect 2464 16708 2470 16720
rect 2587 16711 2645 16717
rect 2587 16708 2599 16711
rect 2464 16680 2599 16708
rect 2464 16668 2470 16680
rect 2587 16677 2599 16680
rect 2633 16708 2645 16711
rect 3050 16708 3056 16720
rect 2633 16680 3056 16708
rect 2633 16677 2645 16680
rect 2587 16671 2645 16677
rect 3050 16668 3056 16680
rect 3108 16668 3114 16720
rect 4801 16711 4859 16717
rect 4801 16677 4813 16711
rect 4847 16708 4859 16711
rect 5350 16708 5356 16720
rect 4847 16680 5356 16708
rect 4847 16677 4859 16680
rect 4801 16671 4859 16677
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4246 16640 4252 16652
rect 4203 16612 4252 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 4522 16600 4528 16652
rect 4580 16640 4586 16652
rect 5445 16643 5503 16649
rect 5445 16640 5457 16643
rect 4580 16612 5457 16640
rect 4580 16600 4586 16612
rect 5445 16609 5457 16612
rect 5491 16609 5503 16643
rect 5445 16603 5503 16609
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2314 16572 2320 16584
rect 2271 16544 2320 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 5460 16572 5488 16603
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 5592 16612 5733 16640
rect 5592 16600 5598 16612
rect 5721 16609 5733 16612
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 5994 16600 6000 16652
rect 6052 16640 6058 16652
rect 6089 16643 6147 16649
rect 6089 16640 6101 16643
rect 6052 16612 6101 16640
rect 6052 16600 6058 16612
rect 6089 16609 6101 16612
rect 6135 16609 6147 16643
rect 7024 16640 7052 16736
rect 10597 16711 10655 16717
rect 10597 16677 10609 16711
rect 10643 16708 10655 16711
rect 11974 16708 11980 16720
rect 10643 16680 11980 16708
rect 10643 16677 10655 16680
rect 10597 16671 10655 16677
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 12158 16708 12164 16720
rect 12119 16680 12164 16708
rect 12158 16668 12164 16680
rect 12216 16668 12222 16720
rect 12710 16668 12716 16720
rect 12768 16708 12774 16720
rect 15396 16717 15424 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 15381 16711 15439 16717
rect 12768 16680 13032 16708
rect 12768 16668 12774 16680
rect 7190 16640 7196 16652
rect 7024 16612 7196 16640
rect 6089 16603 6147 16609
rect 7190 16600 7196 16612
rect 7248 16640 7254 16652
rect 7285 16643 7343 16649
rect 7285 16640 7297 16643
rect 7248 16612 7297 16640
rect 7248 16600 7254 16612
rect 7285 16609 7297 16612
rect 7331 16609 7343 16643
rect 7285 16603 7343 16609
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9824 16612 9873 16640
rect 9824 16600 9830 16612
rect 9861 16609 9873 16612
rect 9907 16640 9919 16643
rect 11238 16640 11244 16652
rect 9907 16612 11244 16640
rect 9907 16609 9919 16612
rect 9861 16603 9919 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11422 16640 11428 16652
rect 11383 16612 11428 16640
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11882 16640 11888 16652
rect 11532 16612 11888 16640
rect 6178 16572 6184 16584
rect 5460 16544 6184 16572
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 10008 16575 10066 16581
rect 10008 16541 10020 16575
rect 10054 16572 10066 16575
rect 10134 16572 10140 16584
rect 10054 16544 10140 16572
rect 10054 16541 10066 16544
rect 10008 16535 10066 16541
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 11146 16572 11152 16584
rect 10284 16544 11152 16572
rect 10284 16532 10290 16544
rect 11146 16532 11152 16544
rect 11204 16572 11210 16584
rect 11532 16572 11560 16612
rect 11882 16600 11888 16612
rect 11940 16640 11946 16652
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 11940 16612 12449 16640
rect 11940 16600 11946 16612
rect 12437 16609 12449 16612
rect 12483 16640 12495 16643
rect 12802 16640 12808 16652
rect 12483 16612 12808 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13004 16649 13032 16680
rect 15381 16677 15393 16711
rect 15427 16677 15439 16711
rect 15381 16671 15439 16677
rect 15473 16711 15531 16717
rect 15473 16677 15485 16711
rect 15519 16708 15531 16711
rect 15746 16708 15752 16720
rect 15519 16680 15752 16708
rect 15519 16677 15531 16680
rect 15473 16671 15531 16677
rect 15746 16668 15752 16680
rect 15804 16668 15810 16720
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16609 13047 16643
rect 12989 16603 13047 16609
rect 11204 16544 11560 16572
rect 11204 16532 11210 16544
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11756 16544 11805 16572
rect 11756 16532 11762 16544
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 13004 16572 13032 16603
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13136 16612 13553 16640
rect 13136 16600 13142 16612
rect 13541 16609 13553 16612
rect 13587 16640 13599 16643
rect 14826 16640 14832 16652
rect 13587 16612 14832 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 24670 16649 24676 16652
rect 24648 16643 24676 16649
rect 24648 16640 24660 16643
rect 24583 16612 24660 16640
rect 24648 16609 24660 16612
rect 24728 16640 24734 16652
rect 25038 16640 25044 16652
rect 24728 16612 25044 16640
rect 24648 16603 24676 16609
rect 24670 16600 24676 16603
rect 24728 16600 24734 16612
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 13262 16572 13268 16584
rect 13004 16544 13268 16572
rect 11793 16535 11851 16541
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 15654 16572 15660 16584
rect 15615 16544 15660 16572
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 2498 16464 2504 16516
rect 2556 16504 2562 16516
rect 3145 16507 3203 16513
rect 3145 16504 3157 16507
rect 2556 16476 3157 16504
rect 2556 16464 2562 16476
rect 3145 16473 3157 16476
rect 3191 16473 3203 16507
rect 3145 16467 3203 16473
rect 6362 16464 6368 16516
rect 6420 16504 6426 16516
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 6420 16476 7481 16504
rect 6420 16464 6426 16476
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 7469 16467 7527 16473
rect 8386 16464 8392 16516
rect 8444 16504 8450 16516
rect 8757 16507 8815 16513
rect 8757 16504 8769 16507
rect 8444 16476 8769 16504
rect 8444 16464 8450 16476
rect 8757 16473 8769 16476
rect 8803 16504 8815 16507
rect 11330 16504 11336 16516
rect 8803 16476 11336 16504
rect 8803 16473 8815 16476
rect 8757 16467 8815 16473
rect 11330 16464 11336 16476
rect 11388 16504 11394 16516
rect 11563 16507 11621 16513
rect 11563 16504 11575 16507
rect 11388 16476 11575 16504
rect 11388 16464 11394 16476
rect 11563 16473 11575 16476
rect 11609 16504 11621 16507
rect 11882 16504 11888 16516
rect 11609 16476 11888 16504
rect 11609 16473 11621 16476
rect 11563 16467 11621 16473
rect 11882 16464 11888 16476
rect 11940 16504 11946 16516
rect 12805 16507 12863 16513
rect 12805 16504 12817 16507
rect 11940 16476 12817 16504
rect 11940 16464 11946 16476
rect 12805 16473 12817 16476
rect 12851 16473 12863 16507
rect 12805 16467 12863 16473
rect 8481 16439 8539 16445
rect 8481 16405 8493 16439
rect 8527 16436 8539 16439
rect 8662 16436 8668 16448
rect 8527 16408 8668 16436
rect 8527 16405 8539 16408
rect 8481 16399 8539 16405
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 10042 16396 10048 16448
rect 10100 16436 10106 16448
rect 10137 16439 10195 16445
rect 10137 16436 10149 16439
rect 10100 16408 10149 16436
rect 10100 16396 10106 16408
rect 10137 16405 10149 16408
rect 10183 16405 10195 16439
rect 10137 16399 10195 16405
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11790 16436 11796 16448
rect 11747 16408 11796 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 18414 16396 18420 16448
rect 18472 16436 18478 16448
rect 24719 16439 24777 16445
rect 24719 16436 24731 16439
rect 18472 16408 24731 16436
rect 18472 16396 18478 16408
rect 24719 16405 24731 16408
rect 24765 16405 24777 16439
rect 24719 16399 24777 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2317 16235 2375 16241
rect 2317 16201 2329 16235
rect 2363 16232 2375 16235
rect 2406 16232 2412 16244
rect 2363 16204 2412 16232
rect 2363 16201 2375 16204
rect 2317 16195 2375 16201
rect 2406 16192 2412 16204
rect 2464 16192 2470 16244
rect 4614 16232 4620 16244
rect 4575 16204 4620 16232
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 4706 16192 4712 16244
rect 4764 16232 4770 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 4764 16204 8217 16232
rect 4764 16192 4770 16204
rect 8205 16201 8217 16204
rect 8251 16232 8263 16235
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 8251 16204 8677 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 8665 16201 8677 16204
rect 8711 16201 8723 16235
rect 8846 16232 8852 16244
rect 8807 16204 8852 16232
rect 8665 16195 8723 16201
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 4632 16096 4660 16192
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 8386 16164 8392 16176
rect 7984 16136 8392 16164
rect 7984 16124 7990 16136
rect 8386 16124 8392 16136
rect 8444 16164 8450 16176
rect 8527 16167 8585 16173
rect 8527 16164 8539 16167
rect 8444 16136 8539 16164
rect 8444 16124 8450 16136
rect 8527 16133 8539 16136
rect 8573 16133 8585 16167
rect 8680 16164 8708 16195
rect 8846 16192 8852 16204
rect 8904 16192 8910 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9140 16204 9873 16232
rect 9140 16164 9168 16204
rect 9861 16201 9873 16204
rect 9907 16232 9919 16235
rect 10042 16232 10048 16244
rect 9907 16204 10048 16232
rect 9907 16201 9919 16204
rect 9861 16195 9919 16201
rect 10042 16192 10048 16204
rect 10100 16232 10106 16244
rect 10870 16232 10876 16244
rect 10100 16204 10876 16232
rect 10100 16192 10106 16204
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11790 16232 11796 16244
rect 11751 16204 11796 16232
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 13078 16232 13084 16244
rect 13039 16204 13084 16232
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 13320 16204 13461 16232
rect 13320 16192 13326 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 15746 16232 15752 16244
rect 15707 16204 15752 16232
rect 13449 16195 13507 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 16117 16235 16175 16241
rect 16117 16232 16129 16235
rect 16080 16204 16129 16232
rect 16080 16192 16086 16204
rect 16117 16201 16129 16204
rect 16163 16201 16175 16235
rect 24670 16232 24676 16244
rect 24631 16204 24676 16232
rect 16117 16195 16175 16201
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 10226 16164 10232 16176
rect 8680 16136 9168 16164
rect 9508 16136 10232 16164
rect 8527 16127 8585 16133
rect 9508 16108 9536 16136
rect 10226 16124 10232 16136
rect 10284 16124 10290 16176
rect 2731 16068 4752 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 1448 16031 1506 16037
rect 1448 15997 1460 16031
rect 1494 16028 1506 16031
rect 1854 16028 1860 16040
rect 1494 16000 1860 16028
rect 1494 15997 1506 16000
rect 1448 15991 1506 15997
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 3050 16028 3056 16040
rect 3011 16000 3056 16028
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 3421 16031 3479 16037
rect 3421 15997 3433 16031
rect 3467 16028 3479 16031
rect 3510 16028 3516 16040
rect 3467 16000 3516 16028
rect 3467 15997 3479 16000
rect 3421 15991 3479 15997
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 3620 16037 3648 16068
rect 4724 16037 4752 16068
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 7156 16068 7205 16096
rect 7156 16056 7162 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 8754 16096 8760 16108
rect 8667 16068 8760 16096
rect 7193 16059 7251 16065
rect 8754 16056 8760 16068
rect 8812 16096 8818 16108
rect 9490 16096 9496 16108
rect 8812 16068 9496 16096
rect 8812 16056 8818 16068
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 10888 16096 10916 16192
rect 11882 16124 11888 16176
rect 11940 16164 11946 16176
rect 12575 16167 12633 16173
rect 12575 16164 12587 16167
rect 11940 16136 12587 16164
rect 11940 16124 11946 16136
rect 12575 16133 12587 16136
rect 12621 16133 12633 16167
rect 12575 16127 12633 16133
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 10888 16068 12173 16096
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12802 16096 12808 16108
rect 12763 16068 12808 16096
rect 12161 16059 12219 16065
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 4709 16031 4767 16037
rect 4709 15997 4721 16031
rect 4755 15997 4767 16031
rect 4709 15991 4767 15997
rect 5261 16031 5319 16037
rect 5261 15997 5273 16031
rect 5307 16028 5319 16031
rect 5350 16028 5356 16040
rect 5307 16000 5356 16028
rect 5307 15997 5319 16000
rect 5261 15991 5319 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 12176 16028 12204 16059
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 15654 16096 15660 16108
rect 15519 16068 15660 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 12667 16031 12725 16037
rect 12667 16028 12679 16031
rect 12176 16000 12679 16028
rect 12667 15997 12679 16000
rect 12713 15997 12725 16031
rect 12667 15991 12725 15997
rect 1535 15963 1593 15969
rect 1535 15929 1547 15963
rect 1581 15960 1593 15963
rect 6546 15960 6552 15972
rect 1581 15932 6552 15960
rect 1581 15929 1593 15932
rect 1535 15923 1593 15929
rect 6546 15920 6552 15932
rect 6604 15920 6610 15972
rect 6914 15960 6920 15972
rect 6875 15932 6920 15960
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7006 15920 7012 15972
rect 7064 15960 7070 15972
rect 8389 15963 8447 15969
rect 7064 15932 7109 15960
rect 7064 15920 7070 15932
rect 8389 15929 8401 15963
rect 8435 15960 8447 15963
rect 8570 15960 8576 15972
rect 8435 15932 8576 15960
rect 8435 15929 8447 15932
rect 8389 15923 8447 15929
rect 8570 15920 8576 15932
rect 8628 15960 8634 15972
rect 8846 15960 8852 15972
rect 8628 15932 8852 15960
rect 8628 15920 8634 15932
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 9398 15920 9404 15972
rect 9456 15960 9462 15972
rect 10321 15963 10379 15969
rect 10321 15960 10333 15963
rect 9456 15932 10333 15960
rect 9456 15920 9462 15932
rect 10321 15929 10333 15932
rect 10367 15929 10379 15963
rect 10321 15923 10379 15929
rect 10413 15963 10471 15969
rect 10413 15929 10425 15963
rect 10459 15960 10471 15963
rect 10686 15960 10692 15972
rect 10459 15932 10692 15960
rect 10459 15929 10471 15932
rect 10413 15923 10471 15929
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 10965 15963 11023 15969
rect 10965 15929 10977 15963
rect 11011 15960 11023 15963
rect 11330 15960 11336 15972
rect 11011 15932 11336 15960
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 11330 15920 11336 15932
rect 11388 15920 11394 15972
rect 12434 15960 12440 15972
rect 12395 15932 12440 15960
rect 12434 15920 12440 15932
rect 12492 15960 12498 15972
rect 13817 15963 13875 15969
rect 13817 15960 13829 15963
rect 12492 15932 13829 15960
rect 12492 15920 12498 15932
rect 13817 15929 13829 15932
rect 13863 15929 13875 15963
rect 14826 15960 14832 15972
rect 14787 15932 14832 15960
rect 13817 15923 13875 15929
rect 14826 15920 14832 15932
rect 14884 15920 14890 15972
rect 14921 15963 14979 15969
rect 14921 15929 14933 15963
rect 14967 15960 14979 15963
rect 15470 15960 15476 15972
rect 14967 15932 15476 15960
rect 14967 15929 14979 15932
rect 14921 15923 14979 15929
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 2869 15895 2927 15901
rect 2869 15892 2881 15895
rect 2372 15864 2881 15892
rect 2372 15852 2378 15864
rect 2869 15861 2881 15864
rect 2915 15861 2927 15895
rect 4246 15892 4252 15904
rect 4207 15864 4252 15892
rect 2869 15855 2927 15861
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5721 15895 5779 15901
rect 5721 15892 5733 15895
rect 5224 15864 5733 15892
rect 5224 15852 5230 15864
rect 5721 15861 5733 15864
rect 5767 15892 5779 15895
rect 5994 15892 6000 15904
rect 5767 15864 6000 15892
rect 5767 15861 5779 15864
rect 5721 15855 5779 15861
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6178 15892 6184 15904
rect 6139 15864 6184 15892
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7024 15892 7052 15920
rect 7926 15892 7932 15904
rect 6687 15864 7052 15892
rect 7887 15864 7932 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 9490 15892 9496 15904
rect 9451 15864 9496 15892
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 11425 15895 11483 15901
rect 11425 15892 11437 15895
rect 9732 15864 11437 15892
rect 9732 15852 9738 15864
rect 11425 15861 11437 15864
rect 11471 15892 11483 15895
rect 11698 15892 11704 15904
rect 11471 15864 11704 15892
rect 11471 15861 11483 15864
rect 11425 15855 11483 15861
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 14645 15895 14703 15901
rect 14645 15861 14657 15895
rect 14691 15892 14703 15895
rect 14936 15892 14964 15923
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 14691 15864 14964 15892
rect 14691 15861 14703 15864
rect 14645 15855 14703 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1535 15691 1593 15697
rect 1535 15657 1547 15691
rect 1581 15688 1593 15691
rect 2130 15688 2136 15700
rect 1581 15660 2136 15688
rect 1581 15657 1593 15660
rect 1535 15651 1593 15657
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3108 15660 3433 15688
rect 3108 15648 3114 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 3421 15651 3479 15657
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 5445 15691 5503 15697
rect 5445 15657 5457 15691
rect 5491 15688 5503 15691
rect 7190 15688 7196 15700
rect 5491 15660 7046 15688
rect 7151 15660 7196 15688
rect 5491 15657 5503 15660
rect 5445 15651 5503 15657
rect 2222 15580 2228 15632
rect 2280 15620 2286 15632
rect 2409 15623 2467 15629
rect 2409 15620 2421 15623
rect 2280 15592 2421 15620
rect 2280 15580 2286 15592
rect 2409 15589 2421 15592
rect 2455 15589 2467 15623
rect 2409 15583 2467 15589
rect 4617 15623 4675 15629
rect 4617 15589 4629 15623
rect 4663 15620 4675 15623
rect 6086 15620 6092 15632
rect 4663 15592 6092 15620
rect 4663 15589 4675 15592
rect 4617 15583 4675 15589
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 6270 15620 6276 15632
rect 6231 15592 6276 15620
rect 6270 15580 6276 15592
rect 6328 15580 6334 15632
rect 6365 15623 6423 15629
rect 6365 15589 6377 15623
rect 6411 15620 6423 15623
rect 7018 15620 7046 15660
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 10192 15660 10241 15688
rect 10192 15648 10198 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 11882 15688 11888 15700
rect 11843 15660 11888 15688
rect 10229 15651 10287 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 13136 15660 13461 15688
rect 13136 15648 13142 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 14826 15688 14832 15700
rect 14787 15660 14832 15688
rect 13449 15651 13507 15657
rect 14826 15648 14832 15660
rect 14884 15688 14890 15700
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 14884 15660 15301 15688
rect 14884 15648 14890 15660
rect 15289 15657 15301 15660
rect 15335 15657 15347 15691
rect 15289 15651 15347 15657
rect 9306 15620 9312 15632
rect 6411 15592 6960 15620
rect 7018 15592 9312 15620
rect 6411 15589 6423 15592
rect 6365 15583 6423 15589
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 1432 15555 1490 15561
rect 1432 15552 1444 15555
rect 1360 15524 1444 15552
rect 1360 15512 1366 15524
rect 1432 15521 1444 15524
rect 1478 15521 1490 15555
rect 2498 15552 2504 15564
rect 2459 15524 2504 15552
rect 1432 15515 1490 15521
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 4522 15512 4528 15564
rect 4580 15552 4586 15564
rect 4764 15555 4822 15561
rect 4764 15552 4776 15555
rect 4580 15524 4776 15552
rect 4580 15512 4586 15524
rect 4764 15521 4776 15524
rect 4810 15521 4822 15555
rect 6932 15552 6960 15592
rect 9306 15580 9312 15592
rect 9364 15580 9370 15632
rect 11057 15623 11115 15629
rect 11057 15589 11069 15623
rect 11103 15620 11115 15623
rect 11146 15620 11152 15632
rect 11103 15592 11152 15620
rect 11103 15589 11115 15592
rect 11057 15583 11115 15589
rect 11146 15580 11152 15592
rect 11204 15620 11210 15632
rect 12437 15623 12495 15629
rect 12437 15620 12449 15623
rect 11204 15592 12449 15620
rect 11204 15580 11210 15592
rect 12437 15589 12449 15592
rect 12483 15589 12495 15623
rect 12437 15583 12495 15589
rect 8018 15552 8024 15564
rect 6932 15524 8024 15552
rect 4764 15515 4822 15521
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 12802 15552 12808 15564
rect 12763 15524 12808 15552
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 16298 15552 16304 15564
rect 16356 15561 16362 15564
rect 16356 15555 16394 15561
rect 15712 15524 16304 15552
rect 15712 15512 15718 15524
rect 16298 15512 16304 15524
rect 16382 15521 16394 15555
rect 16356 15515 16394 15521
rect 16356 15512 16362 15515
rect 4338 15444 4344 15496
rect 4396 15484 4402 15496
rect 4985 15487 5043 15493
rect 4985 15484 4997 15487
rect 4396 15456 4997 15484
rect 4396 15444 4402 15456
rect 4985 15453 4997 15456
rect 5031 15484 5043 15487
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5031 15456 5457 15484
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 5445 15447 5503 15453
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7064 15456 7757 15484
rect 7064 15444 7070 15456
rect 7745 15453 7757 15456
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15484 11023 15487
rect 11238 15484 11244 15496
rect 11011 15456 11244 15484
rect 11011 15453 11023 15456
rect 10965 15447 11023 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 11388 15456 11433 15484
rect 11388 15444 11394 15456
rect 6546 15376 6552 15428
rect 6604 15416 6610 15428
rect 9398 15416 9404 15428
rect 6604 15388 9404 15416
rect 6604 15376 6610 15388
rect 9398 15376 9404 15388
rect 9456 15376 9462 15428
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 11422 15416 11428 15428
rect 11112 15388 11428 15416
rect 11112 15376 11118 15388
rect 11422 15376 11428 15388
rect 11480 15416 11486 15428
rect 12253 15419 12311 15425
rect 12253 15416 12265 15419
rect 11480 15388 12265 15416
rect 11480 15376 11486 15388
rect 12253 15385 12265 15388
rect 12299 15416 12311 15419
rect 12434 15416 12440 15428
rect 12299 15388 12440 15416
rect 12299 15385 12311 15388
rect 12253 15379 12311 15385
rect 12434 15376 12440 15388
rect 12492 15376 12498 15428
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 4893 15351 4951 15357
rect 4893 15348 4905 15351
rect 4764 15320 4905 15348
rect 4764 15308 4770 15320
rect 4893 15317 4905 15320
rect 4939 15317 4951 15351
rect 4893 15311 4951 15317
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 5592 15320 5641 15348
rect 5592 15308 5598 15320
rect 5629 15317 5641 15320
rect 5675 15317 5687 15351
rect 5994 15348 6000 15360
rect 5955 15320 6000 15348
rect 5629 15311 5687 15317
rect 5994 15308 6000 15320
rect 6052 15348 6058 15360
rect 6270 15348 6276 15360
rect 6052 15320 6276 15348
rect 6052 15308 6058 15320
rect 6270 15308 6276 15320
rect 6328 15308 6334 15360
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 6972 15320 7021 15348
rect 6972 15308 6978 15320
rect 7009 15317 7021 15320
rect 7055 15348 7067 15351
rect 7098 15348 7104 15360
rect 7055 15320 7104 15348
rect 7055 15317 7067 15320
rect 7009 15311 7067 15317
rect 7098 15308 7104 15320
rect 7156 15308 7162 15360
rect 7558 15348 7564 15360
rect 7519 15320 7564 15348
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 8846 15348 8852 15360
rect 8807 15320 8852 15348
rect 8846 15308 8852 15320
rect 8904 15348 8910 15360
rect 9766 15348 9772 15360
rect 8904 15320 9772 15348
rect 8904 15308 8910 15320
rect 9766 15308 9772 15320
rect 9824 15348 9830 15360
rect 9861 15351 9919 15357
rect 9861 15348 9873 15351
rect 9824 15320 9873 15348
rect 9824 15308 9830 15320
rect 9861 15317 9873 15320
rect 9907 15317 9919 15351
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 9861 15311 9919 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 16439 15351 16497 15357
rect 16439 15317 16451 15351
rect 16485 15348 16497 15351
rect 16666 15348 16672 15360
rect 16485 15320 16672 15348
rect 16485 15317 16497 15320
rect 16439 15311 16497 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1302 15104 1308 15156
rect 1360 15144 1366 15156
rect 1581 15147 1639 15153
rect 1581 15144 1593 15147
rect 1360 15116 1593 15144
rect 1360 15104 1366 15116
rect 1581 15113 1593 15116
rect 1627 15113 1639 15147
rect 1581 15107 1639 15113
rect 2409 15147 2467 15153
rect 2409 15113 2421 15147
rect 2455 15144 2467 15147
rect 2498 15144 2504 15156
rect 2455 15116 2504 15144
rect 2455 15113 2467 15116
rect 2409 15107 2467 15113
rect 2498 15104 2504 15116
rect 2556 15104 2562 15156
rect 4338 15144 4344 15156
rect 4299 15116 4344 15144
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 4706 15144 4712 15156
rect 4667 15116 4712 15144
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 6638 15144 6644 15156
rect 6599 15116 6644 15144
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 8018 15144 8024 15156
rect 7979 15116 8024 15144
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 8478 15144 8484 15156
rect 8439 15116 8484 15144
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 9306 15104 9312 15156
rect 9364 15144 9370 15156
rect 9674 15144 9680 15156
rect 9364 15116 9680 15144
rect 9364 15104 9370 15116
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 9950 15144 9956 15156
rect 9815 15116 9956 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 11146 15144 11152 15156
rect 11107 15116 11152 15144
rect 11146 15104 11152 15116
rect 11204 15104 11210 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11296 15116 11529 15144
rect 11296 15104 11302 15116
rect 11517 15113 11529 15116
rect 11563 15144 11575 15147
rect 14642 15144 14648 15156
rect 11563 15116 14648 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 14642 15104 14648 15116
rect 14700 15104 14706 15156
rect 16298 15144 16304 15156
rect 16259 15116 16304 15144
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 10686 15036 10692 15088
rect 10744 15076 10750 15088
rect 10781 15079 10839 15085
rect 10781 15076 10793 15079
rect 10744 15048 10793 15076
rect 10744 15036 10750 15048
rect 10781 15045 10793 15048
rect 10827 15076 10839 15079
rect 12802 15076 12808 15088
rect 10827 15048 12808 15076
rect 10827 15045 10839 15048
rect 10781 15039 10839 15045
rect 12802 15036 12808 15048
rect 12860 15036 12866 15088
rect 5261 15011 5319 15017
rect 5261 14977 5273 15011
rect 5307 15008 5319 15011
rect 5718 15008 5724 15020
rect 5307 14980 5724 15008
rect 5307 14977 5319 14980
rect 5261 14971 5319 14977
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 11885 15011 11943 15017
rect 11885 15008 11897 15011
rect 9732 14980 11897 15008
rect 9732 14968 9738 14980
rect 11885 14977 11897 14980
rect 11931 15008 11943 15011
rect 11931 14980 12848 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2869 14943 2927 14949
rect 2869 14940 2881 14943
rect 2087 14912 2881 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 2869 14909 2881 14912
rect 2915 14940 2927 14943
rect 2958 14940 2964 14952
rect 2915 14912 2964 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 7374 14940 7380 14952
rect 6871 14912 7380 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 9861 14943 9919 14949
rect 9861 14909 9873 14943
rect 9907 14940 9919 14943
rect 9950 14940 9956 14952
rect 9907 14912 9956 14940
rect 9907 14909 9919 14912
rect 9861 14903 9919 14909
rect 9950 14900 9956 14912
rect 10008 14940 10014 14952
rect 12253 14943 12311 14949
rect 10008 14912 10818 14940
rect 10008 14900 10014 14912
rect 2777 14875 2835 14881
rect 2777 14841 2789 14875
rect 2823 14872 2835 14875
rect 3231 14875 3289 14881
rect 3231 14872 3243 14875
rect 2823 14844 3243 14872
rect 2823 14841 2835 14844
rect 2777 14835 2835 14841
rect 3231 14841 3243 14844
rect 3277 14872 3289 14875
rect 3878 14872 3884 14884
rect 3277 14844 3884 14872
rect 3277 14841 3289 14844
rect 3231 14835 3289 14841
rect 3878 14832 3884 14844
rect 3936 14832 3942 14884
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 5905 14875 5963 14881
rect 5408 14844 5453 14872
rect 5408 14832 5414 14844
rect 5905 14841 5917 14875
rect 5951 14872 5963 14875
rect 6086 14872 6092 14884
rect 5951 14844 6092 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 6178 14832 6184 14884
rect 6236 14872 6242 14884
rect 6273 14875 6331 14881
rect 6273 14872 6285 14875
rect 6236 14844 6285 14872
rect 6236 14832 6242 14844
rect 6273 14841 6285 14844
rect 6319 14872 6331 14875
rect 7006 14872 7012 14884
rect 6319 14844 7012 14872
rect 6319 14841 6331 14844
rect 6273 14835 6331 14841
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 7187 14875 7245 14881
rect 7187 14841 7199 14875
rect 7233 14841 7245 14875
rect 7187 14835 7245 14841
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5368 14804 5396 14832
rect 5123 14776 5396 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 6638 14804 6644 14816
rect 6420 14776 6644 14804
rect 6420 14764 6426 14776
rect 6638 14764 6644 14776
rect 6696 14804 6702 14816
rect 7202 14804 7230 14835
rect 7282 14832 7288 14884
rect 7340 14872 7346 14884
rect 8573 14875 8631 14881
rect 8573 14872 8585 14875
rect 7340 14844 8585 14872
rect 7340 14832 7346 14844
rect 8573 14841 8585 14844
rect 8619 14841 8631 14875
rect 8573 14835 8631 14841
rect 10042 14832 10048 14884
rect 10100 14872 10106 14884
rect 10182 14875 10240 14881
rect 10182 14872 10194 14875
rect 10100 14844 10194 14872
rect 10100 14832 10106 14844
rect 10182 14841 10194 14844
rect 10228 14841 10240 14875
rect 10790 14872 10818 14912
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12342 14940 12348 14952
rect 12299 14912 12348 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12342 14900 12348 14912
rect 12400 14940 12406 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12400 14912 12449 14940
rect 12400 14900 12406 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12820 14940 12848 14980
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12820 14912 12909 14940
rect 12437 14903 12495 14909
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 10790 14844 12480 14872
rect 10182 14835 10240 14841
rect 7742 14804 7748 14816
rect 6696 14776 7230 14804
rect 7703 14776 7748 14804
rect 6696 14764 6702 14776
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 12452 14804 12480 14844
rect 12529 14807 12587 14813
rect 12529 14804 12541 14807
rect 12452 14776 12541 14804
rect 12529 14773 12541 14776
rect 12575 14773 12587 14807
rect 12529 14767 12587 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 4522 14600 4528 14612
rect 4483 14572 4528 14600
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 5350 14560 5356 14612
rect 5408 14600 5414 14612
rect 7101 14603 7159 14609
rect 5408 14572 6684 14600
rect 5408 14560 5414 14572
rect 2593 14535 2651 14541
rect 2593 14501 2605 14535
rect 2639 14532 2651 14535
rect 2866 14532 2872 14544
rect 2639 14504 2872 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 2866 14492 2872 14504
rect 2924 14532 2930 14544
rect 3786 14532 3792 14544
rect 2924 14504 3792 14532
rect 2924 14492 2930 14504
rect 3786 14492 3792 14504
rect 3844 14492 3850 14544
rect 3878 14492 3884 14544
rect 3936 14532 3942 14544
rect 6362 14532 6368 14544
rect 3936 14504 6368 14532
rect 3936 14492 3942 14504
rect 6362 14492 6368 14504
rect 6420 14532 6426 14544
rect 6502 14535 6560 14541
rect 6502 14532 6514 14535
rect 6420 14504 6514 14532
rect 6420 14492 6426 14504
rect 6502 14501 6514 14504
rect 6548 14501 6560 14535
rect 6656 14532 6684 14572
rect 7101 14569 7113 14603
rect 7147 14600 7159 14603
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 7147 14572 7205 14600
rect 7147 14569 7159 14572
rect 7101 14563 7159 14569
rect 7193 14569 7205 14572
rect 7239 14600 7251 14603
rect 8018 14600 8024 14612
rect 7239 14572 8024 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 12802 14600 12808 14612
rect 12763 14572 12808 14600
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 16850 14600 16856 14612
rect 16811 14572 16856 14600
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 7929 14535 7987 14541
rect 7929 14532 7941 14535
rect 6656 14504 7941 14532
rect 6502 14495 6560 14501
rect 7929 14501 7941 14504
rect 7975 14501 7987 14535
rect 7929 14495 7987 14501
rect 10042 14492 10048 14544
rect 10100 14532 10106 14544
rect 10226 14532 10232 14544
rect 10100 14504 10232 14532
rect 10100 14492 10106 14504
rect 10226 14492 10232 14504
rect 10284 14532 10290 14544
rect 10366 14535 10424 14541
rect 10366 14532 10378 14535
rect 10284 14504 10378 14532
rect 10284 14492 10290 14504
rect 10366 14501 10378 14504
rect 10412 14501 10424 14535
rect 11974 14532 11980 14544
rect 11935 14504 11980 14532
rect 10366 14495 10424 14501
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 4614 14464 4620 14476
rect 4575 14436 4620 14464
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14464 5227 14467
rect 5258 14464 5264 14476
rect 5215 14436 5264 14464
rect 5215 14433 5227 14436
rect 5169 14427 5227 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5718 14464 5724 14476
rect 5631 14436 5724 14464
rect 5718 14424 5724 14436
rect 5776 14464 5782 14476
rect 7282 14464 7288 14476
rect 5776 14436 7288 14464
rect 5776 14424 5782 14436
rect 7282 14424 7288 14436
rect 7340 14424 7346 14476
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7800 14436 8033 14464
rect 7800 14424 7806 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 16666 14464 16672 14476
rect 16627 14436 16672 14464
rect 8021 14427 8079 14433
rect 16666 14424 16672 14436
rect 16724 14424 16730 14476
rect 2222 14356 2228 14408
rect 2280 14396 2286 14408
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 2280 14368 2513 14396
rect 2280 14356 2286 14368
rect 2501 14365 2513 14368
rect 2547 14396 2559 14399
rect 2682 14396 2688 14408
rect 2547 14368 2688 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3142 14396 3148 14408
rect 3103 14368 3148 14396
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 5399 14368 6193 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 6181 14365 6193 14368
rect 6227 14396 6239 14399
rect 6546 14396 6552 14408
rect 6227 14368 6552 14396
rect 6227 14365 6239 14368
rect 6181 14359 6239 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 10042 14396 10048 14408
rect 10003 14368 10048 14396
rect 10042 14356 10048 14368
rect 10100 14356 10106 14408
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11882 14396 11888 14408
rect 11388 14368 11888 14396
rect 11388 14356 11394 14368
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12158 14396 12164 14408
rect 12119 14368 12164 14396
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 6089 14331 6147 14337
rect 6089 14297 6101 14331
rect 6135 14328 6147 14331
rect 7193 14331 7251 14337
rect 7193 14328 7205 14331
rect 6135 14300 7205 14328
rect 6135 14297 6147 14300
rect 6089 14291 6147 14297
rect 7193 14297 7205 14300
rect 7239 14297 7251 14331
rect 7193 14291 7251 14297
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8938 14260 8944 14272
rect 8899 14232 8944 14260
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 10965 14263 11023 14269
rect 10965 14260 10977 14263
rect 10744 14232 10977 14260
rect 10744 14220 10750 14232
rect 10965 14229 10977 14232
rect 11011 14229 11023 14263
rect 11330 14260 11336 14272
rect 11291 14232 11336 14260
rect 10965 14223 11023 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 2866 14056 2872 14068
rect 1811 14028 2872 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 5534 14056 5540 14068
rect 4126 14028 5540 14056
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 3568 13960 3832 13988
rect 3568 13948 3574 13960
rect 3804 13929 3832 13960
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 3789 13923 3847 13929
rect 2823 13892 3740 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 3050 13852 3056 13864
rect 2884 13824 3056 13852
rect 2884 13784 2912 13824
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3712 13861 3740 13892
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 4126 13920 4154 14028
rect 5534 14016 5540 14028
rect 5592 14056 5598 14068
rect 6178 14056 6184 14068
rect 5592 14028 6184 14056
rect 5592 14016 5598 14028
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6273 14059 6331 14065
rect 6273 14025 6285 14059
rect 6319 14056 6331 14059
rect 6362 14056 6368 14068
rect 6319 14028 6368 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7800 14028 7941 14056
rect 7800 14016 7806 14028
rect 7929 14025 7941 14028
rect 7975 14056 7987 14059
rect 8018 14056 8024 14068
rect 7975 14028 8024 14056
rect 7975 14025 7987 14028
rect 7929 14019 7987 14025
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 10134 14056 10140 14068
rect 9646 14028 10140 14056
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 7469 13991 7527 13997
rect 7469 13988 7481 13991
rect 6144 13960 7481 13988
rect 6144 13948 6150 13960
rect 7469 13957 7481 13960
rect 7515 13957 7527 13991
rect 9646 13988 9674 14028
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 10744 14028 11897 14056
rect 10744 14016 10750 14028
rect 11885 14025 11897 14028
rect 11931 14056 11943 14059
rect 11974 14056 11980 14068
rect 11931 14028 11980 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 16666 14056 16672 14068
rect 16627 14028 16672 14056
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 7469 13951 7527 13957
rect 8680 13960 9674 13988
rect 11149 13991 11207 13997
rect 3835 13892 4154 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 4522 13880 4528 13932
rect 4580 13920 4586 13932
rect 5905 13923 5963 13929
rect 4580 13892 5856 13920
rect 4580 13880 4586 13892
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13852 3755 13855
rect 4985 13855 5043 13861
rect 4985 13852 4997 13855
rect 3743 13824 4997 13852
rect 3743 13821 3755 13824
rect 3697 13815 3755 13821
rect 4985 13821 4997 13824
rect 5031 13852 5043 13855
rect 5166 13852 5172 13864
rect 5031 13824 5172 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5258 13812 5264 13864
rect 5316 13852 5322 13864
rect 5534 13852 5540 13864
rect 5316 13824 5540 13852
rect 5316 13812 5322 13824
rect 5534 13812 5540 13824
rect 5592 13852 5598 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5592 13824 5641 13852
rect 5592 13812 5598 13824
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 2424 13756 2912 13784
rect 4341 13787 4399 13793
rect 2424 13728 2452 13756
rect 4341 13753 4353 13787
rect 4387 13784 4399 13787
rect 5276 13784 5304 13812
rect 4387 13756 5304 13784
rect 4387 13753 4399 13756
rect 4341 13747 4399 13753
rect 1854 13716 1860 13728
rect 1815 13688 1860 13716
rect 1854 13676 1860 13688
rect 1912 13676 1918 13728
rect 2406 13716 2412 13728
rect 2367 13688 2412 13716
rect 2406 13676 2412 13688
rect 2464 13676 2470 13728
rect 2958 13716 2964 13728
rect 2919 13688 2964 13716
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 4706 13716 4712 13728
rect 4619 13688 4712 13716
rect 4706 13676 4712 13688
rect 4764 13716 4770 13728
rect 4982 13716 4988 13728
rect 4764 13688 4988 13716
rect 4764 13676 4770 13688
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 5828 13716 5856 13892
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 7374 13920 7380 13932
rect 5951 13892 7380 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 8680 13852 8708 13960
rect 11149 13957 11161 13991
rect 11195 13988 11207 13991
rect 11606 13988 11612 14000
rect 11195 13960 11612 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 11606 13948 11612 13960
rect 11664 13988 11670 14000
rect 12158 13988 12164 14000
rect 11664 13960 12164 13988
rect 11664 13948 11670 13960
rect 12158 13948 12164 13960
rect 12216 13948 12222 14000
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 9306 13920 9312 13932
rect 8812 13892 9312 13920
rect 8812 13880 8818 13892
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 9674 13920 9680 13932
rect 9635 13892 9680 13920
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 10226 13920 10232 13932
rect 10183 13892 10232 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 11330 13920 11336 13932
rect 10643 13892 11336 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 11330 13880 11336 13892
rect 11388 13920 11394 13932
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 11388 13892 12449 13920
rect 11388 13880 11394 13892
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 9088 13855 9146 13861
rect 9088 13852 9100 13855
rect 8404 13824 9100 13852
rect 6914 13784 6920 13796
rect 6875 13756 6920 13784
rect 6914 13744 6920 13756
rect 6972 13744 6978 13796
rect 7006 13744 7012 13796
rect 7064 13784 7070 13796
rect 8018 13784 8024 13796
rect 7064 13756 8024 13784
rect 7064 13744 7070 13756
rect 8018 13744 8024 13756
rect 8076 13744 8082 13796
rect 7190 13716 7196 13728
rect 5828 13688 7196 13716
rect 7190 13676 7196 13688
rect 7248 13716 7254 13728
rect 8404 13725 8432 13824
rect 9088 13821 9100 13824
rect 9134 13821 9146 13855
rect 9088 13815 9146 13821
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9950 13852 9956 13864
rect 9272 13824 9956 13852
rect 9272 13812 9278 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 8938 13784 8944 13796
rect 8899 13756 8944 13784
rect 8938 13744 8944 13756
rect 8996 13744 9002 13796
rect 10689 13787 10747 13793
rect 10689 13753 10701 13787
rect 10735 13784 10747 13787
rect 11330 13784 11336 13796
rect 10735 13756 11336 13784
rect 10735 13753 10747 13756
rect 10689 13747 10747 13753
rect 11330 13744 11336 13756
rect 11388 13784 11394 13796
rect 11517 13787 11575 13793
rect 11517 13784 11529 13787
rect 11388 13756 11529 13784
rect 11388 13744 11394 13756
rect 11517 13753 11529 13756
rect 11563 13753 11575 13787
rect 11517 13747 11575 13753
rect 8389 13719 8447 13725
rect 8389 13716 8401 13719
rect 7248 13688 8401 13716
rect 7248 13676 7254 13688
rect 8389 13685 8401 13688
rect 8435 13685 8447 13719
rect 8754 13716 8760 13728
rect 8715 13688 8760 13716
rect 8389 13679 8447 13685
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2222 13512 2228 13524
rect 2183 13484 2228 13512
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 3510 13512 3516 13524
rect 2332 13484 3188 13512
rect 3471 13484 3516 13512
rect 1464 13379 1522 13385
rect 1464 13345 1476 13379
rect 1510 13376 1522 13379
rect 1670 13376 1676 13388
rect 1510 13348 1676 13376
rect 1510 13345 1522 13348
rect 1464 13339 1522 13345
rect 1670 13336 1676 13348
rect 1728 13376 1734 13388
rect 2332 13376 2360 13484
rect 3160 13456 3188 13484
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 5123 13515 5181 13521
rect 5123 13481 5135 13515
rect 5169 13512 5181 13515
rect 5994 13512 6000 13524
rect 5169 13484 6000 13512
rect 5169 13481 5181 13484
rect 5123 13475 5181 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 6914 13512 6920 13524
rect 6595 13484 6920 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 8113 13515 8171 13521
rect 8113 13512 8125 13515
rect 7524 13484 8125 13512
rect 7524 13472 7530 13484
rect 8113 13481 8125 13484
rect 8159 13481 8171 13515
rect 8113 13475 8171 13481
rect 8849 13515 8907 13521
rect 8849 13481 8861 13515
rect 8895 13512 8907 13515
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8895 13484 9045 13512
rect 8895 13481 8907 13484
rect 8849 13475 8907 13481
rect 9033 13481 9045 13484
rect 9079 13512 9091 13515
rect 9214 13512 9220 13524
rect 9079 13484 9220 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 11882 13512 11888 13524
rect 11843 13484 11888 13512
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 2590 13444 2596 13456
rect 2551 13416 2596 13444
rect 2590 13404 2596 13416
rect 2648 13404 2654 13456
rect 3142 13444 3148 13456
rect 3103 13416 3148 13444
rect 3142 13404 3148 13416
rect 3200 13404 3206 13456
rect 11330 13444 11336 13456
rect 11291 13416 11336 13444
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 1728 13348 2360 13376
rect 1728 13336 1734 13348
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 5020 13379 5078 13385
rect 5020 13376 5032 13379
rect 4948 13348 5032 13376
rect 4948 13336 4954 13348
rect 5020 13345 5032 13348
rect 5066 13345 5078 13379
rect 5020 13339 5078 13345
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6086 13376 6092 13388
rect 6043 13348 6092 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7006 13376 7012 13388
rect 6963 13348 7012 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7156 13348 7481 13376
rect 7156 13336 7162 13348
rect 7469 13345 7481 13348
rect 7515 13376 7527 13379
rect 8294 13376 8300 13388
rect 7515 13348 8300 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 8294 13336 8300 13348
rect 8352 13376 8358 13388
rect 8938 13376 8944 13388
rect 8352 13348 8944 13376
rect 8352 13336 8358 13348
rect 8938 13336 8944 13348
rect 8996 13336 9002 13388
rect 10686 13376 10692 13388
rect 10647 13348 10692 13376
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12196 13379 12254 13385
rect 12196 13376 12208 13379
rect 12124 13348 12208 13376
rect 12124 13336 12130 13348
rect 12196 13345 12208 13348
rect 12242 13345 12254 13379
rect 12196 13339 12254 13345
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 1912 13280 2513 13308
rect 1912 13268 1918 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 7834 13308 7840 13320
rect 7795 13280 7840 13308
rect 2501 13271 2559 13277
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 4246 13200 4252 13252
rect 4304 13240 4310 13252
rect 6135 13243 6193 13249
rect 6135 13240 6147 13243
rect 4304 13212 6147 13240
rect 4304 13200 4310 13212
rect 6135 13209 6147 13212
rect 6181 13209 6193 13243
rect 6135 13203 6193 13209
rect 7634 13243 7692 13249
rect 7634 13209 7646 13243
rect 7680 13240 7692 13243
rect 7926 13240 7932 13252
rect 7680 13212 7932 13240
rect 7680 13209 7692 13212
rect 7634 13203 7692 13209
rect 7926 13200 7932 13212
rect 7984 13240 7990 13252
rect 8386 13240 8392 13252
rect 7984 13212 8392 13240
rect 7984 13200 7990 13212
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 5534 13172 5540 13184
rect 5447 13144 5540 13172
rect 5534 13132 5540 13144
rect 5592 13172 5598 13184
rect 6270 13172 6276 13184
rect 5592 13144 6276 13172
rect 5592 13132 5598 13144
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 7374 13172 7380 13184
rect 7335 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 7742 13172 7748 13184
rect 7655 13144 7748 13172
rect 7742 13132 7748 13144
rect 7800 13172 7806 13184
rect 8849 13175 8907 13181
rect 8849 13172 8861 13175
rect 7800 13144 8861 13172
rect 7800 13132 7806 13144
rect 8849 13141 8861 13144
rect 8895 13141 8907 13175
rect 10042 13172 10048 13184
rect 10003 13144 10048 13172
rect 8849 13135 8907 13141
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 12299 13175 12357 13181
rect 12299 13141 12311 13175
rect 12345 13172 12357 13175
rect 18598 13172 18604 13184
rect 12345 13144 18604 13172
rect 12345 13141 12357 13144
rect 12299 13135 12357 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1670 12968 1676 12980
rect 1631 12940 1676 12968
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 2041 12971 2099 12977
rect 2041 12968 2053 12971
rect 1912 12940 2053 12968
rect 1912 12928 1918 12940
rect 2041 12937 2053 12940
rect 2087 12937 2099 12971
rect 2041 12931 2099 12937
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4948 12940 4997 12968
rect 4948 12928 4954 12940
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 6086 12968 6092 12980
rect 6047 12940 6092 12968
rect 4985 12931 5043 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 6328 12940 7941 12968
rect 6328 12928 6334 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 10686 12968 10692 12980
rect 10647 12940 10692 12968
rect 7929 12931 7987 12937
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 11606 12968 11612 12980
rect 11567 12940 11612 12968
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 12124 12940 12173 12968
rect 12124 12928 12130 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 7190 12860 7196 12912
rect 7248 12900 7254 12912
rect 7607 12903 7665 12909
rect 7607 12900 7619 12903
rect 7248 12872 7619 12900
rect 7248 12860 7254 12872
rect 7607 12869 7619 12872
rect 7653 12869 7665 12903
rect 7742 12900 7748 12912
rect 7703 12872 7748 12900
rect 7607 12863 7665 12869
rect 7742 12860 7748 12872
rect 7800 12900 7806 12912
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 7800 12872 8493 12900
rect 7800 12860 7806 12872
rect 8481 12869 8493 12872
rect 8527 12869 8539 12903
rect 8481 12863 8539 12869
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2590 12832 2596 12844
rect 2547 12804 2596 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 2590 12792 2596 12804
rect 2648 12832 2654 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2648 12804 2789 12832
rect 2648 12792 2654 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 7834 12832 7840 12844
rect 7340 12804 7840 12832
rect 7340 12792 7346 12804
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 10042 12832 10048 12844
rect 10003 12804 10048 12832
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 2866 12764 2872 12776
rect 2827 12736 2872 12764
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 7742 12764 7748 12776
rect 6687 12736 7748 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 9582 12764 9588 12776
rect 9543 12736 9588 12764
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 9732 12736 9965 12764
rect 9732 12724 9738 12736
rect 9953 12733 9965 12736
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 11124 12767 11182 12773
rect 11124 12733 11136 12767
rect 11170 12764 11182 12767
rect 11606 12764 11612 12776
rect 11170 12736 11612 12764
rect 11170 12733 11182 12736
rect 11124 12727 11182 12733
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12764 13415 12767
rect 13814 12764 13820 12776
rect 13403 12736 13820 12764
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 7374 12656 7380 12708
rect 7432 12696 7438 12708
rect 7469 12699 7527 12705
rect 7469 12696 7481 12699
rect 7432 12668 7481 12696
rect 7432 12656 7438 12668
rect 7469 12665 7481 12668
rect 7515 12696 7527 12699
rect 8202 12696 8208 12708
rect 7515 12668 8208 12696
rect 7515 12665 7527 12668
rect 7469 12659 7527 12665
rect 8202 12656 8208 12668
rect 8260 12656 8266 12708
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8941 12699 8999 12705
rect 8941 12696 8953 12699
rect 8352 12668 8953 12696
rect 8352 12656 8358 12668
rect 8941 12665 8953 12668
rect 8987 12696 8999 12699
rect 10962 12696 10968 12708
rect 8987 12668 10968 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 9582 12628 9588 12640
rect 9447 12600 9588 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 11195 12631 11253 12637
rect 11195 12628 11207 12631
rect 10100 12600 11207 12628
rect 10100 12588 10106 12600
rect 11195 12597 11207 12600
rect 11241 12597 11253 12631
rect 11195 12591 11253 12597
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12492 12600 12633 12628
rect 12492 12588 12498 12600
rect 12621 12597 12633 12600
rect 12667 12628 12679 12631
rect 12820 12628 12848 12727
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 13538 12696 13544 12708
rect 13499 12668 13544 12696
rect 13538 12656 13544 12668
rect 13596 12656 13602 12708
rect 12667 12600 12848 12628
rect 12667 12597 12679 12600
rect 12621 12591 12679 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2866 12424 2872 12436
rect 2827 12396 2872 12424
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 9732 12396 9873 12424
rect 9732 12384 9738 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 9861 12387 9919 12393
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 10137 12359 10195 12365
rect 10137 12356 10149 12359
rect 10008 12328 10149 12356
rect 10008 12316 10014 12328
rect 10137 12325 10149 12328
rect 10183 12325 10195 12359
rect 10137 12319 10195 12325
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1578 12288 1584 12300
rect 1443 12260 1584 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1578 12248 1584 12260
rect 1636 12288 1642 12300
rect 2222 12288 2228 12300
rect 1636 12260 2228 12288
rect 1636 12248 1642 12260
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 5074 12248 5080 12300
rect 5132 12288 5138 12300
rect 7742 12288 7748 12300
rect 7800 12297 7806 12300
rect 7800 12291 7838 12297
rect 5132 12260 7748 12288
rect 5132 12248 5138 12260
rect 7742 12248 7748 12260
rect 7826 12257 7838 12291
rect 10226 12288 10232 12300
rect 10187 12260 10232 12288
rect 7800 12251 7838 12257
rect 7800 12248 7806 12251
rect 10226 12248 10232 12260
rect 10284 12288 10290 12300
rect 10870 12288 10876 12300
rect 10284 12260 10876 12288
rect 10284 12248 10290 12260
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11020 12260 11713 12288
rect 11020 12248 11026 12260
rect 11701 12257 11713 12260
rect 11747 12288 11759 12291
rect 12158 12288 12164 12300
rect 11747 12260 12164 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 13262 12288 13268 12300
rect 13223 12260 13268 12288
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 13814 12288 13820 12300
rect 13786 12248 13820 12288
rect 13872 12288 13878 12300
rect 13872 12260 13917 12288
rect 13872 12248 13878 12260
rect 12066 12220 12072 12232
rect 12027 12192 12072 12220
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 12483 12192 12909 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 12897 12189 12909 12192
rect 12943 12220 12955 12223
rect 13786 12220 13814 12248
rect 13998 12220 14004 12232
rect 12943 12192 13814 12220
rect 13959 12192 14004 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 7282 12112 7288 12164
rect 7340 12152 7346 12164
rect 7561 12155 7619 12161
rect 7561 12152 7573 12155
rect 7340 12124 7573 12152
rect 7340 12112 7346 12124
rect 7561 12121 7573 12124
rect 7607 12152 7619 12155
rect 8478 12152 8484 12164
rect 7607 12124 8484 12152
rect 7607 12121 7619 12124
rect 7561 12115 7619 12121
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 106 12044 112 12096
rect 164 12084 170 12096
rect 1581 12087 1639 12093
rect 1581 12084 1593 12087
rect 164 12056 1593 12084
rect 164 12044 170 12056
rect 1581 12053 1593 12056
rect 1627 12053 1639 12087
rect 1581 12047 1639 12053
rect 7883 12087 7941 12093
rect 7883 12053 7895 12087
rect 7929 12084 7941 12087
rect 8110 12084 8116 12096
rect 7929 12056 8116 12084
rect 7929 12053 7941 12056
rect 7883 12047 7941 12053
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 8297 12087 8355 12093
rect 8297 12053 8309 12087
rect 8343 12084 8355 12087
rect 8386 12084 8392 12096
rect 8343 12056 8392 12084
rect 8343 12053 8355 12056
rect 8297 12047 8355 12053
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 10778 12084 10784 12096
rect 10192 12056 10784 12084
rect 10192 12044 10198 12056
rect 10778 12044 10784 12056
rect 10836 12084 10842 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10836 12056 11161 12084
rect 10836 12044 10842 12056
rect 11149 12053 11161 12056
rect 11195 12084 11207 12087
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 11195 12056 11529 12084
rect 11195 12053 11207 12056
rect 11149 12047 11207 12053
rect 11517 12053 11529 12056
rect 11563 12084 11575 12087
rect 11839 12087 11897 12093
rect 11839 12084 11851 12087
rect 11563 12056 11851 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 11839 12053 11851 12056
rect 11885 12053 11897 12087
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11839 12047 11897 12053
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 14366 12084 14372 12096
rect 14327 12056 14372 12084
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 15838 12084 15844 12096
rect 15799 12056 15844 12084
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2222 11880 2228 11892
rect 2183 11852 2228 11880
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 9861 11883 9919 11889
rect 9861 11849 9873 11883
rect 9907 11880 9919 11883
rect 9950 11880 9956 11892
rect 9907 11852 9956 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 9950 11840 9956 11852
rect 10008 11880 10014 11892
rect 10781 11883 10839 11889
rect 10781 11880 10793 11883
rect 10008 11852 10793 11880
rect 10008 11840 10014 11852
rect 10781 11849 10793 11852
rect 10827 11880 10839 11883
rect 11974 11880 11980 11892
rect 10827 11852 11980 11880
rect 10827 11849 10839 11852
rect 10781 11843 10839 11849
rect 11974 11840 11980 11852
rect 12032 11880 12038 11892
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 12032 11852 12081 11880
rect 12032 11840 12038 11852
rect 12069 11849 12081 11852
rect 12115 11849 12127 11883
rect 12069 11843 12127 11849
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 24765 11883 24823 11889
rect 13872 11852 13917 11880
rect 13872 11840 13878 11852
rect 24765 11849 24777 11883
rect 24811 11880 24823 11883
rect 27614 11880 27620 11892
rect 24811 11852 27620 11880
rect 24811 11849 24823 11852
rect 24765 11843 24823 11849
rect 27614 11840 27620 11852
rect 27672 11840 27678 11892
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 10686 11812 10692 11824
rect 8812 11784 10692 11812
rect 8812 11772 8818 11784
rect 10686 11772 10692 11784
rect 10744 11812 10750 11824
rect 10744 11784 11002 11812
rect 10744 11772 10750 11784
rect 1535 11747 1593 11753
rect 1535 11713 1547 11747
rect 1581 11744 1593 11747
rect 8938 11744 8944 11756
rect 1581 11716 8944 11744
rect 1581 11713 1593 11716
rect 1535 11707 1593 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 10873 11747 10931 11753
rect 9324 11716 9674 11744
rect 1118 11636 1124 11688
rect 1176 11676 1182 11688
rect 9324 11685 9352 11716
rect 1432 11679 1490 11685
rect 1432 11676 1444 11679
rect 1176 11648 1444 11676
rect 1176 11636 1182 11648
rect 1432 11645 1444 11648
rect 1478 11676 1490 11679
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1478 11648 1869 11676
rect 1478 11645 1490 11648
rect 1432 11639 1490 11645
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 1857 11639 1915 11645
rect 8496 11648 9321 11676
rect 8496 11552 8524 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9646 11676 9674 11716
rect 10873 11713 10885 11747
rect 10919 11744 10931 11747
rect 10974 11744 11002 11784
rect 15838 11744 15844 11756
rect 10919 11716 11002 11744
rect 15799 11716 15844 11744
rect 10919 11713 10931 11716
rect 10873 11707 10931 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16206 11744 16212 11756
rect 16167 11716 16212 11744
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 10652 11679 10710 11685
rect 9646 11648 10456 11676
rect 9309 11639 9367 11645
rect 8665 11611 8723 11617
rect 8665 11577 8677 11611
rect 8711 11608 8723 11611
rect 8754 11608 8760 11620
rect 8711 11580 8760 11608
rect 8711 11577 8723 11580
rect 8665 11571 8723 11577
rect 8754 11568 8760 11580
rect 8812 11568 8818 11620
rect 10226 11568 10232 11620
rect 10284 11568 10290 11620
rect 8478 11540 8484 11552
rect 8439 11512 8484 11540
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10137 11543 10195 11549
rect 10137 11540 10149 11543
rect 10008 11512 10149 11540
rect 10008 11500 10014 11512
rect 10137 11509 10149 11512
rect 10183 11540 10195 11543
rect 10244 11540 10272 11568
rect 10183 11512 10272 11540
rect 10428 11540 10456 11648
rect 10652 11645 10664 11679
rect 10698 11676 10710 11679
rect 10778 11676 10784 11688
rect 10698 11648 10784 11676
rect 10698 11645 10710 11648
rect 10652 11639 10710 11645
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11020 11648 11713 11676
rect 11020 11636 11026 11648
rect 11701 11645 11713 11648
rect 11747 11676 11759 11679
rect 12066 11676 12072 11688
rect 11747 11648 12072 11676
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12618 11676 12624 11688
rect 12579 11648 12624 11676
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 14366 11676 14372 11688
rect 14327 11648 14372 11676
rect 14366 11636 14372 11648
rect 14424 11636 14430 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 15654 11676 15660 11688
rect 14967 11648 15660 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 24210 11636 24216 11688
rect 24268 11676 24274 11688
rect 24581 11679 24639 11685
rect 24581 11676 24593 11679
rect 24268 11648 24593 11676
rect 24268 11636 24274 11648
rect 24581 11645 24593 11648
rect 24627 11676 24639 11679
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 24627 11648 25145 11676
rect 24627 11645 24639 11648
rect 24581 11639 24639 11645
rect 25133 11645 25145 11648
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 10505 11611 10563 11617
rect 10505 11577 10517 11611
rect 10551 11608 10563 11611
rect 11330 11608 11336 11620
rect 10551 11580 11336 11608
rect 10551 11577 10563 11580
rect 10505 11571 10563 11577
rect 11330 11568 11336 11580
rect 11388 11568 11394 11620
rect 13170 11608 13176 11620
rect 13131 11580 13176 11608
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 15580 11580 15945 11608
rect 15580 11552 15608 11580
rect 15933 11577 15945 11580
rect 15979 11577 15991 11611
rect 15933 11571 15991 11577
rect 10962 11540 10968 11552
rect 10428 11512 10968 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11146 11540 11152 11552
rect 11107 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 13262 11540 13268 11552
rect 12952 11512 13268 11540
rect 12952 11500 12958 11512
rect 13262 11500 13268 11512
rect 13320 11540 13326 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13320 11512 13461 11540
rect 13320 11500 13326 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 15562 11540 15568 11552
rect 15523 11512 15568 11540
rect 13449 11503 13507 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 10686 11336 10692 11348
rect 10647 11308 10692 11336
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 12618 11336 12624 11348
rect 12579 11308 12624 11336
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 14366 11336 14372 11348
rect 14327 11308 14372 11336
rect 14366 11296 14372 11308
rect 14424 11336 14430 11348
rect 14424 11308 15516 11336
rect 14424 11296 14430 11308
rect 15488 11280 15516 11308
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 16853 11339 16911 11345
rect 16853 11336 16865 11339
rect 15896 11308 16865 11336
rect 15896 11296 15902 11308
rect 16853 11305 16865 11308
rect 16899 11305 16911 11339
rect 16853 11299 16911 11305
rect 13811 11271 13869 11277
rect 13811 11237 13823 11271
rect 13857 11268 13869 11271
rect 13906 11268 13912 11280
rect 13857 11240 13912 11268
rect 13857 11237 13869 11240
rect 13811 11231 13869 11237
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 15470 11268 15476 11280
rect 15383 11240 15476 11268
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10229 11203 10287 11209
rect 10229 11200 10241 11203
rect 10192 11172 10241 11200
rect 10192 11160 10198 11172
rect 10229 11169 10241 11172
rect 10275 11200 10287 11203
rect 11146 11200 11152 11212
rect 10275 11172 11152 11200
rect 10275 11169 10287 11172
rect 10229 11163 10287 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11514 11200 11520 11212
rect 11475 11172 11520 11200
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11200 13507 11203
rect 13538 11200 13544 11212
rect 13495 11172 13544 11200
rect 13495 11169 13507 11172
rect 13449 11163 13507 11169
rect 13538 11160 13544 11172
rect 13596 11200 13602 11212
rect 14274 11200 14280 11212
rect 13596 11172 14280 11200
rect 13596 11160 13602 11172
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 10410 11132 10416 11144
rect 10371 11104 10416 11132
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 11238 11132 11244 11144
rect 11199 11104 11244 11132
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 15378 11132 15384 11144
rect 15339 11104 15384 11132
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15396 11064 15424 11092
rect 16942 11064 16948 11076
rect 15396 11036 16948 11064
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 11149 10999 11207 11005
rect 11149 10965 11161 10999
rect 11195 10996 11207 10999
rect 11330 10996 11336 11008
rect 11195 10968 11336 10996
rect 11195 10965 11207 10968
rect 11149 10959 11207 10965
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 12158 10956 12164 11008
rect 12216 10996 12222 11008
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 12216 10968 12265 10996
rect 12216 10956 12222 10968
rect 12253 10965 12265 10968
rect 12299 10965 12311 10999
rect 16298 10996 16304 11008
rect 16259 10968 16304 10996
rect 12253 10959 12311 10965
rect 16298 10956 16304 10968
rect 16356 10956 16362 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 10134 10792 10140 10804
rect 10095 10764 10140 10792
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11514 10792 11520 10804
rect 11475 10764 11520 10792
rect 11514 10752 11520 10764
rect 11572 10792 11578 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11572 10764 11805 10792
rect 11572 10752 11578 10764
rect 11793 10761 11805 10764
rect 11839 10792 11851 10795
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11839 10764 12173 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 12161 10761 12173 10764
rect 12207 10792 12219 10795
rect 12618 10792 12624 10804
rect 12207 10764 12624 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 13906 10792 13912 10804
rect 13587 10764 13912 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 11882 10684 11888 10736
rect 11940 10724 11946 10736
rect 13556 10724 13584 10755
rect 13906 10752 13912 10764
rect 13964 10792 13970 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13964 10764 14013 10792
rect 13964 10752 13970 10764
rect 14001 10761 14013 10764
rect 14047 10792 14059 10795
rect 15470 10792 15476 10804
rect 14047 10764 14596 10792
rect 15431 10764 15476 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 11940 10696 13584 10724
rect 11940 10684 11946 10696
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10468 10628 10609 10656
rect 10468 10616 10474 10628
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 10962 10656 10968 10668
rect 10643 10628 10968 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12710 10656 12716 10668
rect 12575 10628 12716 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 12802 10616 12808 10668
rect 12860 10656 12866 10668
rect 12860 10628 12905 10656
rect 12860 10616 12866 10628
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 14056 10628 14197 10656
rect 14056 10616 14062 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 14568 10588 14596 10764
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 15712 10764 15761 10792
rect 15712 10752 15718 10764
rect 15749 10761 15761 10764
rect 15795 10761 15807 10795
rect 16942 10792 16948 10804
rect 16903 10764 16948 10792
rect 15749 10755 15807 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 24946 10792 24952 10804
rect 24811 10764 24952 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 16577 10727 16635 10733
rect 16577 10724 16589 10727
rect 15896 10696 16589 10724
rect 15896 10684 15902 10696
rect 16577 10693 16589 10696
rect 16623 10693 16635 10727
rect 16577 10687 16635 10693
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16298 10656 16304 10668
rect 16071 10628 16304 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 14424 10560 14596 10588
rect 14424 10548 14430 10560
rect 10505 10523 10563 10529
rect 10505 10489 10517 10523
rect 10551 10520 10563 10523
rect 10959 10523 11017 10529
rect 10959 10520 10971 10523
rect 10551 10492 10971 10520
rect 10551 10489 10563 10492
rect 10505 10483 10563 10489
rect 10959 10489 10971 10492
rect 11005 10520 11017 10523
rect 11882 10520 11888 10532
rect 11005 10492 11888 10520
rect 11005 10489 11017 10492
rect 10959 10483 11017 10489
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 14568 10529 14596 10560
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10588 24639 10591
rect 24627 10560 25268 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 14547 10523 14605 10529
rect 12676 10492 12721 10520
rect 12676 10480 12682 10492
rect 14547 10489 14559 10523
rect 14593 10489 14605 10523
rect 14547 10483 14605 10489
rect 16117 10523 16175 10529
rect 16117 10489 16129 10523
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 9674 10452 9680 10464
rect 9635 10424 9680 10452
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 15105 10455 15163 10461
rect 15105 10421 15117 10455
rect 15151 10452 15163 10455
rect 15286 10452 15292 10464
rect 15151 10424 15292 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15654 10412 15660 10464
rect 15712 10452 15718 10464
rect 16132 10452 16160 10483
rect 25240 10464 25268 10560
rect 25222 10452 25228 10464
rect 15712 10424 16160 10452
rect 25183 10424 25228 10452
rect 15712 10412 15718 10424
rect 25222 10412 25228 10424
rect 25280 10412 25286 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 10962 10248 10968 10260
rect 10923 10220 10968 10248
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11882 10248 11888 10260
rect 11843 10220 11888 10248
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12526 10248 12532 10260
rect 12483 10220 12532 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 14274 10248 14280 10260
rect 14235 10220 14280 10248
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 24765 10251 24823 10257
rect 24765 10217 24777 10251
rect 24811 10248 24823 10251
rect 27614 10248 27620 10260
rect 24811 10220 27620 10248
rect 24811 10217 24823 10220
rect 24765 10211 24823 10217
rect 27614 10208 27620 10220
rect 27672 10208 27678 10260
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13449 10183 13507 10189
rect 13449 10180 13461 10183
rect 13228 10152 13461 10180
rect 13228 10140 13234 10152
rect 13449 10149 13461 10152
rect 13495 10149 13507 10183
rect 13449 10143 13507 10149
rect 13998 10140 14004 10192
rect 14056 10180 14062 10192
rect 14645 10183 14703 10189
rect 14645 10180 14657 10183
rect 14056 10152 14657 10180
rect 14056 10140 14062 10152
rect 14645 10149 14657 10152
rect 14691 10149 14703 10183
rect 14645 10143 14703 10149
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15657 10183 15715 10189
rect 15657 10180 15669 10183
rect 15344 10152 15669 10180
rect 15344 10140 15350 10152
rect 15657 10149 15669 10152
rect 15703 10149 15715 10183
rect 16206 10180 16212 10192
rect 16167 10152 16212 10180
rect 15657 10143 15715 10149
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10060 10044 10088 10075
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 10413 10115 10471 10121
rect 10413 10112 10425 10115
rect 10192 10084 10425 10112
rect 10192 10072 10198 10084
rect 10413 10081 10425 10084
rect 10459 10081 10471 10115
rect 16224 10112 16252 10140
rect 17034 10112 17040 10124
rect 17092 10121 17098 10124
rect 17092 10115 17130 10121
rect 16224 10084 17040 10112
rect 10413 10075 10471 10081
rect 17034 10072 17040 10084
rect 17118 10081 17130 10115
rect 24578 10112 24584 10124
rect 24539 10084 24584 10112
rect 17092 10075 17130 10081
rect 17092 10072 17098 10075
rect 24578 10072 24584 10084
rect 24636 10072 24642 10124
rect 10226 10044 10232 10056
rect 10060 10016 10232 10044
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 10735 10016 11529 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 11517 10013 11529 10016
rect 11563 10044 11575 10047
rect 12342 10044 12348 10056
rect 11563 10016 12348 10044
rect 11563 10013 11575 10016
rect 11517 10007 11575 10013
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10044 15623 10047
rect 15654 10044 15660 10056
rect 15611 10016 15660 10044
rect 15611 10013 15623 10016
rect 15565 10007 15623 10013
rect 12710 9936 12716 9988
rect 12768 9976 12774 9988
rect 13648 9976 13676 10007
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 12768 9948 13676 9976
rect 17175 9979 17233 9985
rect 12768 9936 12774 9948
rect 17175 9945 17187 9979
rect 17221 9976 17233 9979
rect 18874 9976 18880 9988
rect 17221 9948 18880 9976
rect 17221 9945 17233 9948
rect 17175 9939 17233 9945
rect 18874 9936 18880 9948
rect 18932 9936 18938 9988
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 10134 9704 10140 9716
rect 9723 9676 10140 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 11882 9704 11888 9716
rect 11843 9676 11888 9704
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 12253 9707 12311 9713
rect 12253 9673 12265 9707
rect 12299 9704 12311 9707
rect 12526 9704 12532 9716
rect 12299 9676 12532 9704
rect 12299 9673 12311 9676
rect 12253 9667 12311 9673
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 12802 9704 12808 9716
rect 12636 9676 12808 9704
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 10686 9596 10692 9648
rect 10744 9636 10750 9648
rect 11425 9639 11483 9645
rect 11425 9636 11437 9639
rect 10744 9608 11437 9636
rect 10744 9596 10750 9608
rect 11425 9605 11437 9608
rect 11471 9636 11483 9639
rect 12636 9636 12664 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13228 9676 13461 9704
rect 13228 9664 13234 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 15197 9707 15255 9713
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 15286 9704 15292 9716
rect 15243 9676 15292 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 15562 9704 15568 9716
rect 15523 9676 15568 9704
rect 15562 9664 15568 9676
rect 15620 9664 15626 9716
rect 17034 9704 17040 9716
rect 16995 9676 17040 9704
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 24670 9704 24676 9716
rect 24631 9676 24676 9704
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 25222 9664 25228 9716
rect 25280 9704 25286 9716
rect 25363 9707 25421 9713
rect 25363 9704 25375 9707
rect 25280 9676 25375 9704
rect 25280 9664 25286 9676
rect 25363 9673 25375 9676
rect 25409 9673 25421 9707
rect 25363 9667 25421 9673
rect 11471 9608 12664 9636
rect 11471 9605 11483 9608
rect 11425 9599 11483 9605
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 13081 9639 13139 9645
rect 13081 9636 13093 9639
rect 12768 9608 13093 9636
rect 12768 9596 12774 9608
rect 13081 9605 13093 9608
rect 13127 9605 13139 9639
rect 13081 9599 13139 9605
rect 13354 9596 13360 9648
rect 13412 9636 13418 9648
rect 13909 9639 13967 9645
rect 13909 9636 13921 9639
rect 13412 9608 13921 9636
rect 13412 9596 13418 9608
rect 13909 9605 13921 9608
rect 13955 9636 13967 9639
rect 23382 9636 23388 9648
rect 13955 9608 23388 9636
rect 13955 9605 13967 9608
rect 13909 9599 13967 9605
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12802 9568 12808 9580
rect 12575 9540 12808 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1443 9472 2084 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 2056 9373 2084 9472
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15344 9472 15393 9500
rect 15344 9460 15350 9472
rect 15381 9469 15393 9472
rect 15427 9500 15439 9503
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 15427 9472 16313 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 16301 9469 16313 9472
rect 16347 9469 16359 9503
rect 23753 9503 23811 9509
rect 23753 9500 23765 9503
rect 16301 9463 16359 9469
rect 23492 9472 23765 9500
rect 10870 9432 10876 9444
rect 10831 9404 10876 9432
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10965 9435 11023 9441
rect 10965 9401 10977 9435
rect 11011 9432 11023 9435
rect 11238 9432 11244 9444
rect 11011 9404 11244 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 9490 9364 9496 9376
rect 2087 9336 9496 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10045 9367 10103 9373
rect 10045 9333 10057 9367
rect 10091 9364 10103 9367
rect 10134 9364 10140 9376
rect 10091 9336 10140 9364
rect 10091 9333 10103 9336
rect 10045 9327 10103 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10689 9367 10747 9373
rect 10689 9333 10701 9367
rect 10735 9364 10747 9367
rect 10980 9364 11008 9395
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 12618 9392 12624 9444
rect 12676 9432 12682 9444
rect 12676 9404 12721 9432
rect 12676 9392 12682 9404
rect 23492 9376 23520 9472
rect 23753 9469 23765 9472
rect 23799 9469 23811 9503
rect 23753 9463 23811 9469
rect 24578 9460 24584 9512
rect 24636 9500 24642 9512
rect 25292 9503 25350 9509
rect 25292 9500 25304 9503
rect 24636 9472 25304 9500
rect 24636 9460 24642 9472
rect 25292 9469 25304 9472
rect 25338 9500 25350 9503
rect 25685 9503 25743 9509
rect 25685 9500 25697 9503
rect 25338 9472 25697 9500
rect 25338 9469 25350 9472
rect 25292 9463 25350 9469
rect 25685 9469 25697 9472
rect 25731 9469 25743 9503
rect 25685 9463 25743 9469
rect 23474 9364 23480 9376
rect 10735 9336 11008 9364
rect 23435 9336 23480 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 23474 9324 23480 9336
rect 23532 9324 23538 9376
rect 24118 9364 24124 9376
rect 24079 9336 24124 9364
rect 24118 9324 24124 9336
rect 24176 9324 24182 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 10459 9163 10517 9169
rect 10459 9160 10471 9163
rect 9548 9132 10471 9160
rect 9548 9120 9554 9132
rect 10459 9129 10471 9132
rect 10505 9129 10517 9163
rect 10870 9160 10876 9172
rect 10831 9132 10876 9160
rect 10459 9123 10517 9129
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 12342 9160 12348 9172
rect 12303 9132 12348 9160
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 15654 9160 15660 9172
rect 15611 9132 15660 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 8202 9052 8208 9104
rect 8260 9092 8266 9104
rect 11330 9092 11336 9104
rect 8260 9064 11336 9092
rect 8260 9052 8266 9064
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 24029 9095 24087 9101
rect 24029 9061 24041 9095
rect 24075 9092 24087 9095
rect 24118 9092 24124 9104
rect 24075 9064 24124 9092
rect 24075 9061 24087 9064
rect 24029 9055 24087 9061
rect 24118 9052 24124 9064
rect 24176 9052 24182 9104
rect 24578 9092 24584 9104
rect 24539 9064 24584 9092
rect 24578 9052 24584 9064
rect 24636 9052 24642 9104
rect 7374 8984 7380 9036
rect 7432 9024 7438 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 7432 8996 7481 9024
rect 7432 8984 7438 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 7558 8984 7564 9036
rect 7616 9024 7622 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 7616 8996 7665 9024
rect 7616 8984 7622 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 10388 9027 10446 9033
rect 10388 8993 10400 9027
rect 10434 9024 10446 9027
rect 10686 9024 10692 9036
rect 10434 8996 10692 9024
rect 10434 8993 10446 8996
rect 10388 8987 10446 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8036 8888 8064 8919
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 11701 8959 11759 8965
rect 11701 8956 11713 8959
rect 8812 8928 11713 8956
rect 8812 8916 8818 8928
rect 11701 8925 11713 8928
rect 11747 8956 11759 8959
rect 11882 8956 11888 8968
rect 11747 8928 11888 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8956 22891 8959
rect 23382 8956 23388 8968
rect 22879 8928 23388 8956
rect 22879 8925 22891 8928
rect 22833 8919 22891 8925
rect 23382 8916 23388 8928
rect 23440 8956 23446 8968
rect 23937 8959 23995 8965
rect 23937 8956 23949 8959
rect 23440 8928 23949 8956
rect 23440 8916 23446 8928
rect 23937 8925 23949 8928
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 8386 8888 8392 8900
rect 8036 8860 8392 8888
rect 8386 8848 8392 8860
rect 8444 8888 8450 8900
rect 8444 8860 11284 8888
rect 8444 8848 8450 8860
rect 11256 8832 11284 8860
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8297 8823 8355 8829
rect 8297 8820 8309 8823
rect 8260 8792 8309 8820
rect 8260 8780 8266 8792
rect 8297 8789 8309 8792
rect 8343 8789 8355 8823
rect 8297 8783 8355 8789
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 11471 8823 11529 8829
rect 11471 8820 11483 8823
rect 11296 8792 11483 8820
rect 11296 8780 11302 8792
rect 11471 8789 11483 8792
rect 11517 8789 11529 8823
rect 11606 8820 11612 8832
rect 11567 8792 11612 8820
rect 11471 8783 11529 8789
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 11974 8820 11980 8832
rect 11935 8792 11980 8820
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 14458 8820 14464 8832
rect 14419 8792 14464 8820
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 24854 8820 24860 8832
rect 24815 8792 24860 8820
rect 24854 8780 24860 8792
rect 24912 8780 24918 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10686 8616 10692 8628
rect 10459 8588 10692 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11882 8616 11888 8628
rect 11843 8588 11888 8616
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 14366 8616 14372 8628
rect 14327 8588 14372 8616
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 23382 8616 23388 8628
rect 23343 8588 23388 8616
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 23937 8619 23995 8625
rect 23937 8585 23949 8619
rect 23983 8616 23995 8619
rect 24118 8616 24124 8628
rect 23983 8588 24124 8616
rect 23983 8585 23995 8588
rect 23937 8579 23995 8585
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 8018 8508 8024 8560
rect 8076 8548 8082 8560
rect 8481 8551 8539 8557
rect 8481 8548 8493 8551
rect 8076 8520 8493 8548
rect 8076 8508 8082 8520
rect 8481 8517 8493 8520
rect 8527 8517 8539 8551
rect 24670 8548 24676 8560
rect 24631 8520 24676 8548
rect 8481 8511 8539 8517
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 8754 8480 8760 8492
rect 8619 8452 8760 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10928 8452 11069 8480
rect 10928 8440 10934 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 14458 8480 14464 8492
rect 13679 8452 14464 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 24121 8483 24179 8489
rect 24121 8449 24133 8483
rect 24167 8480 24179 8483
rect 24854 8480 24860 8492
rect 24167 8452 24860 8480
rect 24167 8449 24179 8452
rect 24121 8443 24179 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2038 8412 2044 8424
rect 1443 8384 2044 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 8352 8415 8410 8421
rect 8352 8381 8364 8415
rect 8398 8381 8410 8415
rect 8352 8375 8410 8381
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8381 12955 8415
rect 13354 8412 13360 8424
rect 13315 8384 13360 8412
rect 12897 8375 12955 8381
rect 1762 8304 1768 8356
rect 1820 8344 1826 8356
rect 2406 8344 2412 8356
rect 1820 8316 2412 8344
rect 1820 8304 1826 8316
rect 2406 8304 2412 8316
rect 2464 8344 2470 8356
rect 8202 8344 8208 8356
rect 2464 8316 8208 8344
rect 2464 8304 2470 8316
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8367 8344 8395 8375
rect 8570 8344 8576 8356
rect 8367 8316 8576 8344
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 12912 8288 12940 8375
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 15381 8415 15439 8421
rect 15381 8381 15393 8415
rect 15427 8412 15439 8415
rect 15427 8384 19334 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 14366 8304 14372 8356
rect 14424 8344 14430 8356
rect 14782 8347 14840 8353
rect 14782 8344 14794 8347
rect 14424 8316 14794 8344
rect 14424 8304 14430 8316
rect 14782 8313 14794 8316
rect 14828 8344 14840 8347
rect 15654 8344 15660 8356
rect 14828 8316 15660 8344
rect 14828 8313 14840 8316
rect 14782 8307 14840 8313
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 19306 8344 19334 8384
rect 23474 8344 23480 8356
rect 19306 8316 23480 8344
rect 23474 8304 23480 8316
rect 23532 8344 23538 8356
rect 24213 8347 24271 8353
rect 24213 8344 24225 8347
rect 23532 8316 24225 8344
rect 23532 8304 23538 8316
rect 24213 8313 24225 8316
rect 24259 8344 24271 8347
rect 25041 8347 25099 8353
rect 25041 8344 25053 8347
rect 24259 8316 25053 8344
rect 24259 8313 24271 8316
rect 24213 8307 24271 8313
rect 25041 8313 25053 8316
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 2038 8276 2044 8288
rect 1999 8248 2044 8276
rect 2038 8236 2044 8248
rect 2096 8236 2102 8288
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 7101 8279 7159 8285
rect 7101 8276 7113 8279
rect 6604 8248 7113 8276
rect 6604 8236 6610 8248
rect 7101 8245 7113 8248
rect 7147 8276 7159 8279
rect 7374 8276 7380 8288
rect 7147 8248 7380 8276
rect 7147 8245 7159 8248
rect 7101 8239 7159 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7558 8276 7564 8288
rect 7519 8248 7564 8276
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 8018 8276 8024 8288
rect 7979 8248 8024 8276
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 8846 8276 8852 8288
rect 8807 8248 8852 8276
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 10965 8279 11023 8285
rect 10965 8245 10977 8279
rect 11011 8276 11023 8279
rect 11238 8276 11244 8288
rect 11011 8248 11244 8276
rect 11011 8245 11023 8248
rect 10965 8239 11023 8245
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 11480 8248 11529 8276
rect 11480 8236 11486 8248
rect 11517 8245 11529 8248
rect 11563 8276 11575 8279
rect 11606 8276 11612 8288
rect 11563 8248 11612 8276
rect 11563 8245 11575 8248
rect 11517 8239 11575 8245
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12805 8279 12863 8285
rect 12805 8245 12817 8279
rect 12851 8276 12863 8279
rect 12894 8276 12900 8288
rect 12851 8248 12900 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 6236 8044 7665 8072
rect 6236 8032 6242 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8754 8072 8760 8084
rect 8343 8044 8760 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 11330 8072 11336 8084
rect 11291 8044 11336 8072
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12032 8044 12909 8072
rect 12032 8032 12038 8044
rect 12897 8041 12909 8044
rect 12943 8072 12955 8075
rect 13354 8072 13360 8084
rect 12943 8044 13360 8072
rect 12943 8041 12955 8044
rect 12897 8035 12955 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 15654 8072 15660 8084
rect 15615 8044 15660 8072
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 27614 8072 27620 8084
rect 23446 8044 27620 8072
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 7190 7936 7196 7948
rect 7055 7908 7196 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 11514 7936 11520 7948
rect 11475 7908 11520 7936
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 11974 7936 11980 7948
rect 11935 7908 11980 7936
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 13262 7936 13268 7948
rect 13223 7908 13268 7936
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 13372 7936 13400 8032
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13372 7908 13737 7936
rect 13725 7905 13737 7908
rect 13771 7936 13783 7939
rect 14458 7936 14464 7948
rect 13771 7908 14464 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 23198 7945 23204 7948
rect 23176 7939 23204 7945
rect 23176 7936 23188 7939
rect 23111 7908 23188 7936
rect 23176 7905 23188 7908
rect 23256 7936 23262 7948
rect 23446 7936 23474 8044
rect 27614 8032 27620 8044
rect 27672 8032 27678 8084
rect 24305 8007 24363 8013
rect 24305 7973 24317 8007
rect 24351 8004 24363 8007
rect 24670 8004 24676 8016
rect 24351 7976 24676 8004
rect 24351 7973 24363 7976
rect 24305 7967 24363 7973
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 24854 8004 24860 8016
rect 24815 7976 24860 8004
rect 24854 7964 24860 7976
rect 24912 7964 24918 8016
rect 23256 7908 23474 7936
rect 23176 7899 23204 7905
rect 23198 7896 23204 7899
rect 23256 7896 23262 7908
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 6696 7840 7389 7868
rect 6696 7828 6702 7840
rect 7377 7837 7389 7840
rect 7423 7868 7435 7871
rect 8478 7868 8484 7880
rect 7423 7840 8484 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 8478 7828 8484 7840
rect 8536 7868 8542 7880
rect 10962 7868 10968 7880
rect 8536 7840 10968 7868
rect 8536 7828 8542 7840
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 12250 7868 12256 7880
rect 12211 7840 12256 7868
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 14001 7871 14059 7877
rect 14001 7837 14013 7871
rect 14047 7868 14059 7871
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 14047 7840 15301 7868
rect 14047 7837 14059 7840
rect 14001 7831 14059 7837
rect 15289 7837 15301 7840
rect 15335 7868 15347 7871
rect 15654 7868 15660 7880
rect 15335 7840 15660 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15654 7828 15660 7840
rect 15712 7828 15718 7880
rect 24213 7871 24271 7877
rect 24213 7837 24225 7871
rect 24259 7837 24271 7871
rect 24213 7831 24271 7837
rect 7174 7803 7232 7809
rect 7174 7769 7186 7803
rect 7220 7800 7232 7803
rect 7558 7800 7564 7812
rect 7220 7772 7564 7800
rect 7220 7769 7232 7772
rect 7174 7763 7232 7769
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 24228 7800 24256 7831
rect 24762 7800 24768 7812
rect 24228 7772 24768 7800
rect 24762 7760 24768 7772
rect 24820 7760 24826 7812
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7064 7704 7297 7732
rect 7064 7692 7070 7704
rect 7285 7701 7297 7704
rect 7331 7732 7343 7735
rect 8018 7732 8024 7744
rect 7331 7704 8024 7732
rect 7331 7701 7343 7704
rect 7285 7695 7343 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 8570 7732 8576 7744
rect 8531 7704 8576 7732
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 10870 7732 10876 7744
rect 10831 7704 10876 7732
rect 10870 7692 10876 7704
rect 10928 7732 10934 7744
rect 12158 7732 12164 7744
rect 10928 7704 12164 7732
rect 10928 7692 10934 7704
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 14366 7732 14372 7744
rect 14327 7704 14372 7732
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 16206 7732 16212 7744
rect 16167 7704 16212 7732
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 23247 7735 23305 7741
rect 23247 7701 23259 7735
rect 23293 7732 23305 7735
rect 24118 7732 24124 7744
rect 23293 7704 24124 7732
rect 23293 7701 23305 7704
rect 23247 7695 23305 7701
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 1535 7531 1593 7537
rect 1535 7528 1547 7531
rect 1452 7500 1547 7528
rect 1452 7488 1458 7500
rect 1535 7497 1547 7500
rect 1581 7497 1593 7531
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 1535 7491 1593 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 8570 7528 8576 7540
rect 7331 7500 8576 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 8570 7488 8576 7500
rect 8628 7528 8634 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 8628 7500 10241 7528
rect 8628 7488 8634 7500
rect 10229 7497 10241 7500
rect 10275 7528 10287 7531
rect 10778 7528 10784 7540
rect 10275 7500 10784 7528
rect 10275 7497 10287 7500
rect 10229 7491 10287 7497
rect 10778 7488 10784 7500
rect 10836 7528 10842 7540
rect 10919 7531 10977 7537
rect 10919 7528 10931 7531
rect 10836 7500 10931 7528
rect 10836 7488 10842 7500
rect 10919 7497 10931 7500
rect 10965 7497 10977 7531
rect 10919 7491 10977 7497
rect 11514 7488 11520 7540
rect 11572 7528 11578 7540
rect 13262 7528 13268 7540
rect 11572 7500 13268 7528
rect 11572 7488 11578 7500
rect 13262 7488 13268 7500
rect 13320 7528 13326 7540
rect 14274 7528 14280 7540
rect 13320 7500 14280 7528
rect 13320 7488 13326 7500
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 14458 7528 14464 7540
rect 14419 7500 14464 7528
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 15654 7528 15660 7540
rect 15615 7500 15660 7528
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 23198 7528 23204 7540
rect 23159 7500 23204 7528
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 9950 7460 9956 7472
rect 8076 7432 9956 7460
rect 8076 7420 8082 7432
rect 9950 7420 9956 7432
rect 10008 7460 10014 7472
rect 10597 7463 10655 7469
rect 10597 7460 10609 7463
rect 10008 7432 10609 7460
rect 10008 7420 10014 7432
rect 10597 7429 10609 7432
rect 10643 7460 10655 7463
rect 11057 7463 11115 7469
rect 11057 7460 11069 7463
rect 10643 7432 11069 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 11057 7429 11069 7432
rect 11103 7460 11115 7463
rect 11422 7460 11428 7472
rect 11103 7432 11428 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 11422 7420 11428 7432
rect 11480 7420 11486 7472
rect 15381 7463 15439 7469
rect 15381 7429 15393 7463
rect 15427 7460 15439 7463
rect 15562 7460 15568 7472
rect 15427 7432 15568 7460
rect 15427 7429 15439 7432
rect 15381 7423 15439 7429
rect 15562 7420 15568 7432
rect 15620 7420 15626 7472
rect 24854 7460 24860 7472
rect 24815 7432 24860 7460
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 6273 7395 6331 7401
rect 6273 7361 6285 7395
rect 6319 7392 6331 7395
rect 6319 7364 7696 7392
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 7668 7336 7696 7364
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 11020 7364 11161 7392
rect 11020 7352 11026 7364
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 11563 7364 13814 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 198 7284 204 7336
rect 256 7324 262 7336
rect 1432 7327 1490 7333
rect 1432 7324 1444 7327
rect 256 7296 1444 7324
rect 256 7284 262 7296
rect 1432 7293 1444 7296
rect 1478 7324 1490 7327
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1478 7296 1869 7324
rect 1478 7293 1490 7296
rect 1432 7287 1490 7293
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 1857 7287 1915 7293
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 3651 7296 4353 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 4341 7293 4353 7296
rect 4387 7324 4399 7327
rect 4982 7324 4988 7336
rect 4387 7296 4988 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 7190 7324 7196 7336
rect 7151 7296 7196 7324
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7708 7296 7757 7324
rect 7708 7284 7714 7296
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 8987 7296 9137 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 9125 7293 9137 7296
rect 9171 7324 9183 7327
rect 9398 7324 9404 7336
rect 9171 7296 9404 7324
rect 9171 7293 9183 7296
rect 9125 7287 9183 7293
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 12894 7324 12900 7336
rect 12807 7296 12900 7324
rect 12894 7284 12900 7296
rect 12952 7324 12958 7336
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 12952 7296 13461 7324
rect 12952 7284 12958 7296
rect 13449 7293 13461 7296
rect 13495 7293 13507 7327
rect 13786 7324 13814 7364
rect 24118 7352 24124 7404
rect 24176 7392 24182 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 24176 7364 24317 7392
rect 24176 7352 24182 7364
rect 24305 7361 24317 7364
rect 24351 7392 24363 7395
rect 25593 7395 25651 7401
rect 25593 7392 25605 7395
rect 24351 7364 25605 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 25593 7361 25605 7364
rect 25639 7361 25651 7395
rect 25593 7355 25651 7361
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13786 7296 14013 7324
rect 13449 7287 13507 7293
rect 14001 7293 14013 7296
rect 14047 7324 14059 7327
rect 14366 7324 14372 7336
rect 14047 7296 14372 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 14366 7284 14372 7296
rect 14424 7324 14430 7336
rect 15930 7324 15936 7336
rect 14424 7296 15936 7324
rect 14424 7284 14430 7296
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 4433 7259 4491 7265
rect 4433 7225 4445 7259
rect 4479 7256 4491 7259
rect 6914 7256 6920 7268
rect 4479 7228 6920 7256
rect 4479 7225 4491 7228
rect 4433 7219 4491 7225
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7208 7256 7236 7284
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 7208 7228 8217 7256
rect 8205 7225 8217 7228
rect 8251 7225 8263 7259
rect 9766 7256 9772 7268
rect 9727 7228 9772 7256
rect 8205 7219 8263 7225
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 10778 7256 10784 7268
rect 10739 7228 10784 7256
rect 10778 7216 10784 7228
rect 10836 7216 10842 7268
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 11974 7256 11980 7268
rect 11664 7228 11980 7256
rect 11664 7216 11670 7228
rect 11974 7216 11980 7228
rect 12032 7256 12038 7268
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 12032 7228 12173 7256
rect 12032 7216 12038 7228
rect 12161 7225 12173 7228
rect 12207 7225 12219 7259
rect 12161 7219 12219 7225
rect 7006 7188 7012 7200
rect 6967 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 10134 7188 10140 7200
rect 8076 7160 10140 7188
rect 8076 7148 8082 7160
rect 10134 7148 10140 7160
rect 10192 7188 10198 7200
rect 11514 7188 11520 7200
rect 10192 7160 11520 7188
rect 10192 7148 10198 7160
rect 11514 7148 11520 7160
rect 11572 7188 11578 7200
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11572 7160 11805 7188
rect 11572 7148 11578 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 11793 7151 11851 7157
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12912 7197 12940 7284
rect 14182 7256 14188 7268
rect 14143 7228 14188 7256
rect 14182 7216 14188 7228
rect 14240 7216 14246 7268
rect 24397 7259 24455 7265
rect 24397 7225 24409 7259
rect 24443 7225 24455 7259
rect 24397 7219 24455 7225
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12124 7160 12909 7188
rect 12124 7148 12130 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 24118 7188 24124 7200
rect 24031 7160 24124 7188
rect 12897 7151 12955 7157
rect 24118 7148 24124 7160
rect 24176 7188 24182 7200
rect 24412 7188 24440 7219
rect 24176 7160 24440 7188
rect 24176 7148 24182 7160
rect 24486 7148 24492 7200
rect 24544 7188 24550 7200
rect 24670 7188 24676 7200
rect 24544 7160 24676 7188
rect 24544 7148 24550 7160
rect 24670 7148 24676 7160
rect 24728 7188 24734 7200
rect 25225 7191 25283 7197
rect 25225 7188 25237 7191
rect 24728 7160 25237 7188
rect 24728 7148 24734 7160
rect 25225 7157 25237 7160
rect 25271 7157 25283 7191
rect 25225 7151 25283 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 15378 6984 15384 6996
rect 15339 6956 15384 6984
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 24118 6984 24124 6996
rect 24079 6956 24124 6984
rect 24118 6944 24124 6956
rect 24176 6944 24182 6996
rect 7190 6916 7196 6928
rect 7151 6888 7196 6916
rect 7190 6876 7196 6888
rect 7248 6916 7254 6928
rect 7837 6919 7895 6925
rect 7837 6916 7849 6919
rect 7248 6888 7849 6916
rect 7248 6876 7254 6888
rect 7837 6885 7849 6888
rect 7883 6885 7895 6919
rect 13538 6916 13544 6928
rect 13499 6888 13544 6916
rect 7837 6879 7895 6885
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 1670 6848 1676 6860
rect 1631 6820 1676 6848
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 1857 6851 1915 6857
rect 1857 6817 1869 6851
rect 1903 6848 1915 6851
rect 1946 6848 1952 6860
rect 1903 6820 1952 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 6546 6848 6552 6860
rect 6507 6820 6552 6848
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 8018 6848 8024 6860
rect 7979 6820 8024 6848
rect 8018 6808 8024 6820
rect 8076 6808 8082 6860
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 8846 6848 8852 6860
rect 8619 6820 8852 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 11149 6851 11207 6857
rect 11149 6817 11161 6851
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 8754 6780 8760 6792
rect 2271 6752 4154 6780
rect 8667 6752 8760 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 4126 6712 4154 6752
rect 8754 6740 8760 6752
rect 8812 6780 8818 6792
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8812 6752 9045 6780
rect 8812 6740 8818 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 10226 6712 10232 6724
rect 4126 6684 10232 6712
rect 10226 6672 10232 6684
rect 10284 6712 10290 6724
rect 10778 6712 10784 6724
rect 10284 6684 10784 6712
rect 10284 6672 10290 6684
rect 10778 6672 10784 6684
rect 10836 6712 10842 6724
rect 11164 6712 11192 6811
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 14332 6820 15301 6848
rect 14332 6808 14338 6820
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 15654 6848 15660 6860
rect 15335 6820 15660 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6848 15899 6851
rect 15930 6848 15936 6860
rect 15887 6820 15936 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 23934 6808 23940 6860
rect 23992 6848 23998 6860
rect 24486 6848 24492 6860
rect 23992 6820 24492 6848
rect 23992 6808 23998 6820
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 25409 6851 25467 6857
rect 25409 6817 25421 6851
rect 25455 6848 25467 6851
rect 25498 6848 25504 6860
rect 25455 6820 25504 6848
rect 25455 6817 25467 6820
rect 25409 6811 25467 6817
rect 25498 6808 25504 6820
rect 25556 6808 25562 6860
rect 11238 6740 11244 6792
rect 11296 6780 11302 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11296 6752 11529 6780
rect 11296 6740 11302 6752
rect 11517 6749 11529 6752
rect 11563 6780 11575 6783
rect 11882 6780 11888 6792
rect 11563 6752 11888 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 14090 6780 14096 6792
rect 13495 6752 13814 6780
rect 14051 6752 14096 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 11422 6712 11428 6724
rect 10836 6684 11192 6712
rect 11383 6684 11428 6712
rect 10836 6672 10842 6684
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 13786 6712 13814 6752
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 13998 6712 14004 6724
rect 13786 6684 14004 6712
rect 13998 6672 14004 6684
rect 14056 6712 14062 6724
rect 22094 6712 22100 6724
rect 14056 6684 22100 6712
rect 14056 6672 14062 6684
rect 22094 6672 22100 6684
rect 22152 6672 22158 6724
rect 24026 6672 24032 6724
rect 24084 6712 24090 6724
rect 25547 6715 25605 6721
rect 25547 6712 25559 6715
rect 24084 6684 25559 6712
rect 24084 6672 24090 6684
rect 25547 6681 25559 6684
rect 25593 6681 25605 6715
rect 25547 6675 25605 6681
rect 7558 6644 7564 6656
rect 7519 6616 7564 6644
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 10962 6644 10968 6656
rect 10919 6616 10968 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11330 6653 11336 6656
rect 11314 6647 11336 6653
rect 11314 6613 11326 6647
rect 11314 6607 11336 6613
rect 11330 6604 11336 6607
rect 11388 6604 11394 6656
rect 11606 6644 11612 6656
rect 11567 6616 11612 6644
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 24854 6644 24860 6656
rect 24815 6616 24860 6644
rect 24854 6604 24860 6616
rect 24912 6604 24918 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 8018 6440 8024 6452
rect 5040 6412 8024 6440
rect 5040 6400 5046 6412
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 9398 6440 9404 6452
rect 9359 6412 9404 6440
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 10226 6440 10232 6452
rect 10187 6412 10232 6440
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11480 6412 11805 6440
rect 11480 6400 11486 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 11793 6403 11851 6409
rect 13786 6412 14565 6440
rect 6181 6375 6239 6381
rect 6181 6341 6193 6375
rect 6227 6372 6239 6375
rect 8846 6372 8852 6384
rect 6227 6344 8852 6372
rect 6227 6341 6239 6344
rect 6181 6335 6239 6341
rect 1854 6304 1860 6316
rect 1688 6276 1860 6304
rect 1688 6245 1716 6276
rect 1854 6264 1860 6276
rect 1912 6304 1918 6316
rect 3145 6307 3203 6313
rect 3145 6304 3157 6307
rect 1912 6276 3157 6304
rect 1912 6264 1918 6276
rect 3145 6273 3157 6276
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6205 1731 6239
rect 1673 6199 1731 6205
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 1946 6236 1952 6248
rect 1820 6208 1865 6236
rect 1907 6208 1952 6236
rect 1820 6196 1826 6208
rect 1946 6196 1952 6208
rect 2004 6236 2010 6248
rect 2409 6239 2467 6245
rect 2409 6236 2421 6239
rect 2004 6208 2421 6236
rect 2004 6196 2010 6208
rect 2409 6205 2421 6208
rect 2455 6236 2467 6239
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 2455 6208 2789 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2777 6205 2789 6208
rect 2823 6205 2835 6239
rect 6914 6236 6920 6248
rect 6875 6208 6920 6236
rect 2777 6199 2835 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7484 6245 7512 6344
rect 8846 6332 8852 6344
rect 8904 6372 8910 6384
rect 9677 6375 9735 6381
rect 9677 6372 9689 6375
rect 8904 6344 9689 6372
rect 8904 6332 8910 6344
rect 9677 6341 9689 6344
rect 9723 6341 9735 6375
rect 9677 6335 9735 6341
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 13357 6375 13415 6381
rect 13357 6372 13369 6375
rect 12768 6344 13369 6372
rect 12768 6332 12774 6344
rect 13357 6341 13369 6344
rect 13403 6372 13415 6375
rect 13538 6372 13544 6384
rect 13403 6344 13544 6372
rect 13403 6341 13415 6344
rect 13357 6335 13415 6341
rect 13538 6332 13544 6344
rect 13596 6372 13602 6384
rect 13633 6375 13691 6381
rect 13633 6372 13645 6375
rect 13596 6344 13645 6372
rect 13596 6332 13602 6344
rect 13633 6341 13645 6344
rect 13679 6341 13691 6375
rect 13633 6335 13691 6341
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6304 8539 6307
rect 8754 6304 8760 6316
rect 8527 6276 8760 6304
rect 8527 6273 8539 6276
rect 8481 6267 8539 6273
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 12066 6304 12072 6316
rect 10796 6276 12072 6304
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 9674 6236 9680 6248
rect 7469 6199 7527 6205
rect 7944 6208 9680 6236
rect 7650 6168 7656 6180
rect 7611 6140 7656 6168
rect 7650 6128 7656 6140
rect 7708 6128 7714 6180
rect 6546 6100 6552 6112
rect 6507 6072 6552 6100
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7944 6100 7972 6208
rect 9674 6196 9680 6208
rect 9732 6236 9738 6248
rect 10796 6245 10824 6276
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12308 6276 12449 6304
rect 12308 6264 12314 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 9732 6208 10609 6236
rect 9732 6196 9738 6208
rect 10597 6205 10609 6208
rect 10643 6236 10655 6239
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10643 6208 10793 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 10870 6196 10876 6248
rect 10928 6236 10934 6248
rect 11241 6239 11299 6245
rect 11241 6236 11253 6239
rect 10928 6208 11253 6236
rect 10928 6196 10934 6208
rect 11241 6205 11253 6208
rect 11287 6236 11299 6239
rect 11606 6236 11612 6248
rect 11287 6208 11612 6236
rect 11287 6205 11299 6208
rect 11241 6199 11299 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 8843 6171 8901 6177
rect 8843 6137 8855 6171
rect 8889 6168 8901 6171
rect 8938 6168 8944 6180
rect 8889 6140 8944 6168
rect 8889 6137 8901 6140
rect 8843 6131 8901 6137
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 11514 6168 11520 6180
rect 11475 6140 11520 6168
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 12758 6171 12816 6177
rect 12758 6137 12770 6171
rect 12804 6168 12816 6171
rect 13786 6168 13814 6412
rect 14553 6409 14565 6412
rect 14599 6440 14611 6443
rect 14826 6440 14832 6452
rect 14599 6412 14832 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 14826 6400 14832 6412
rect 14884 6440 14890 6452
rect 15562 6440 15568 6452
rect 14884 6412 15568 6440
rect 14884 6400 14890 6412
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 15841 6443 15899 6449
rect 15841 6440 15853 6443
rect 15712 6412 15853 6440
rect 15712 6400 15718 6412
rect 15841 6409 15853 6412
rect 15887 6409 15899 6443
rect 15841 6403 15899 6409
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 15988 6412 16221 6440
rect 15988 6400 15994 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 23934 6440 23940 6452
rect 23895 6412 23940 6440
rect 16209 6403 16267 6409
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 13998 6372 14004 6384
rect 13959 6344 14004 6372
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 25498 6372 25504 6384
rect 25411 6344 25504 6372
rect 25498 6332 25504 6344
rect 25556 6372 25562 6384
rect 27614 6372 27620 6384
rect 25556 6344 27620 6372
rect 25556 6332 25562 6344
rect 27614 6332 27620 6344
rect 27672 6332 27678 6384
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6304 14703 6307
rect 14734 6304 14740 6316
rect 14691 6276 14740 6304
rect 14691 6273 14703 6276
rect 14645 6267 14703 6273
rect 14734 6264 14740 6276
rect 14792 6304 14798 6316
rect 15378 6304 15384 6316
rect 14792 6276 15384 6304
rect 14792 6264 14798 6276
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 23290 6264 23296 6316
rect 23348 6304 23354 6316
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 23348 6276 24133 6304
rect 23348 6264 23354 6276
rect 24121 6273 24133 6276
rect 24167 6304 24179 6307
rect 25041 6307 25099 6313
rect 25041 6304 25053 6307
rect 24167 6276 25053 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 25041 6273 25053 6276
rect 25087 6273 25099 6307
rect 25041 6267 25099 6273
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6236 15623 6239
rect 15611 6208 19334 6236
rect 15611 6205 15623 6208
rect 15565 6199 15623 6205
rect 12804 6140 13814 6168
rect 12804 6137 12816 6140
rect 12758 6131 12816 6137
rect 12158 6100 12164 6112
rect 6972 6072 7972 6100
rect 12119 6072 12164 6100
rect 6972 6060 6978 6072
rect 12158 6060 12164 6072
rect 12216 6100 12222 6112
rect 12773 6100 12801 6131
rect 14826 6128 14832 6180
rect 14884 6168 14890 6180
rect 14966 6171 15024 6177
rect 14966 6168 14978 6171
rect 14884 6140 14978 6168
rect 14884 6128 14890 6140
rect 14966 6137 14978 6140
rect 15012 6137 15024 6171
rect 19306 6168 19334 6208
rect 23385 6171 23443 6177
rect 23385 6168 23397 6171
rect 19306 6140 23397 6168
rect 14966 6131 15024 6137
rect 23385 6137 23397 6140
rect 23431 6168 23443 6171
rect 23842 6168 23848 6180
rect 23431 6140 23848 6168
rect 23431 6137 23443 6140
rect 23385 6131 23443 6137
rect 23842 6128 23848 6140
rect 23900 6168 23906 6180
rect 24213 6171 24271 6177
rect 24213 6168 24225 6171
rect 23900 6140 24225 6168
rect 23900 6128 23906 6140
rect 24213 6137 24225 6140
rect 24259 6137 24271 6171
rect 24762 6168 24768 6180
rect 24723 6140 24768 6168
rect 24213 6131 24271 6137
rect 24762 6128 24768 6140
rect 24820 6128 24826 6180
rect 18230 6100 18236 6112
rect 12216 6072 12801 6100
rect 18191 6072 18236 6100
rect 12216 6060 12222 6072
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1670 5896 1676 5908
rect 1631 5868 1676 5896
rect 1670 5856 1676 5868
rect 1728 5896 1734 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 1728 5868 2421 5896
rect 1728 5856 1734 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 2409 5859 2467 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 10870 5896 10876 5908
rect 10831 5868 10876 5896
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11238 5896 11244 5908
rect 11199 5868 11244 5896
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 11517 5899 11575 5905
rect 11517 5896 11529 5899
rect 11388 5868 11529 5896
rect 11388 5856 11394 5868
rect 11517 5865 11529 5868
rect 11563 5865 11575 5899
rect 11517 5859 11575 5865
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 12437 5899 12495 5905
rect 12437 5896 12449 5899
rect 12308 5868 12449 5896
rect 12308 5856 12314 5868
rect 12437 5865 12449 5868
rect 12483 5865 12495 5899
rect 12437 5859 12495 5865
rect 14090 5856 14096 5908
rect 14148 5896 14154 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14148 5868 14289 5896
rect 14148 5856 14154 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14734 5896 14740 5908
rect 14695 5868 14740 5896
rect 14277 5859 14335 5865
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 15620 5868 15669 5896
rect 15620 5856 15626 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 8110 5828 8116 5840
rect 8071 5800 8116 5828
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 9398 5828 9404 5840
rect 8260 5800 9404 5828
rect 8260 5788 8266 5800
rect 9398 5788 9404 5800
rect 9456 5788 9462 5840
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 9824 5800 9873 5828
rect 9824 5788 9830 5800
rect 9861 5797 9873 5800
rect 9907 5797 9919 5831
rect 9861 5791 9919 5797
rect 12158 5788 12164 5840
rect 12216 5828 12222 5840
rect 13034 5831 13092 5837
rect 13034 5828 13046 5831
rect 12216 5800 13046 5828
rect 12216 5788 12222 5800
rect 13034 5797 13046 5800
rect 13080 5797 13092 5831
rect 13034 5791 13092 5797
rect 18598 5788 18604 5840
rect 18656 5828 18662 5840
rect 18693 5831 18751 5837
rect 18693 5828 18705 5831
rect 18656 5800 18705 5828
rect 18656 5788 18662 5800
rect 18693 5797 18705 5800
rect 18739 5797 18751 5831
rect 18693 5791 18751 5797
rect 1854 5760 1860 5772
rect 1815 5732 1860 5760
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 11514 5720 11520 5772
rect 11572 5760 11578 5772
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 11572 5732 12725 5760
rect 11572 5720 11578 5732
rect 12713 5729 12725 5732
rect 12759 5760 12771 5763
rect 13722 5760 13728 5772
rect 12759 5732 13728 5760
rect 12759 5729 12771 5732
rect 12713 5723 12771 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 14240 5732 15301 5760
rect 14240 5720 14246 5732
rect 15289 5729 15301 5732
rect 15335 5760 15347 5763
rect 16850 5760 16856 5772
rect 15335 5732 16856 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 23842 5760 23848 5772
rect 23803 5732 23848 5760
rect 23842 5720 23848 5732
rect 23900 5720 23906 5772
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5692 9827 5695
rect 9950 5692 9956 5704
rect 9815 5664 9956 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 8665 5627 8723 5633
rect 8665 5593 8677 5627
rect 8711 5624 8723 5627
rect 9858 5624 9864 5636
rect 8711 5596 9864 5624
rect 8711 5593 8723 5596
rect 8665 5587 8723 5593
rect 9858 5584 9864 5596
rect 9916 5624 9922 5636
rect 10060 5624 10088 5655
rect 17862 5652 17868 5704
rect 17920 5692 17926 5704
rect 18230 5692 18236 5704
rect 17920 5664 18236 5692
rect 17920 5652 17926 5664
rect 18230 5652 18236 5664
rect 18288 5692 18294 5704
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 18288 5664 18613 5692
rect 18288 5652 18294 5664
rect 18601 5661 18613 5664
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 19150 5624 19156 5636
rect 9916 5596 10088 5624
rect 19111 5596 19156 5624
rect 9916 5584 9922 5596
rect 19150 5584 19156 5596
rect 19208 5584 19214 5636
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9033 5559 9091 5565
rect 9033 5556 9045 5559
rect 8996 5528 9045 5556
rect 8996 5516 9002 5528
rect 9033 5525 9045 5528
rect 9079 5525 9091 5559
rect 13630 5556 13636 5568
rect 13591 5528 13636 5556
rect 9033 5519 9091 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 16209 5559 16267 5565
rect 16209 5525 16221 5559
rect 16255 5556 16267 5559
rect 18230 5556 18236 5568
rect 16255 5528 18236 5556
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 24026 5556 24032 5568
rect 23987 5528 24032 5556
rect 24026 5516 24032 5528
rect 24084 5516 24090 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 1854 5352 1860 5364
rect 1360 5324 1860 5352
rect 1360 5312 1366 5324
rect 1854 5312 1860 5324
rect 1912 5352 1918 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 1912 5324 2237 5352
rect 1912 5312 1918 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5352 7803 5355
rect 8110 5352 8116 5364
rect 7791 5324 8116 5352
rect 7791 5321 7803 5324
rect 7745 5315 7803 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 9861 5355 9919 5361
rect 9861 5352 9873 5355
rect 9824 5324 9873 5352
rect 9824 5312 9830 5324
rect 9861 5321 9873 5324
rect 9907 5321 9919 5355
rect 9861 5315 9919 5321
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 11514 5352 11520 5364
rect 10008 5324 11520 5352
rect 10008 5312 10014 5324
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 13630 5312 13636 5364
rect 13688 5352 13694 5364
rect 14093 5355 14151 5361
rect 14093 5352 14105 5355
rect 13688 5324 14105 5352
rect 13688 5312 13694 5324
rect 14093 5321 14105 5324
rect 14139 5352 14151 5355
rect 14458 5352 14464 5364
rect 14139 5324 14464 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15562 5352 15568 5364
rect 15427 5324 15568 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17862 5352 17868 5364
rect 17823 5324 17868 5352
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 23477 5355 23535 5361
rect 23477 5321 23489 5355
rect 23523 5352 23535 5355
rect 23842 5352 23848 5364
rect 23523 5324 23848 5352
rect 23523 5321 23535 5324
rect 23477 5315 23535 5321
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 24026 5352 24032 5364
rect 23987 5324 24032 5352
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 8021 5287 8079 5293
rect 8021 5253 8033 5287
rect 8067 5284 8079 5287
rect 8202 5284 8208 5296
rect 8067 5256 8208 5284
rect 8067 5253 8079 5256
rect 8021 5247 8079 5253
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 8938 5244 8944 5296
rect 8996 5284 9002 5296
rect 12158 5284 12164 5296
rect 8996 5256 12164 5284
rect 8996 5244 9002 5256
rect 12158 5244 12164 5256
rect 12216 5244 12222 5296
rect 13722 5284 13728 5296
rect 13683 5256 13728 5284
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 19797 5287 19855 5293
rect 19797 5284 19809 5287
rect 18800 5256 19809 5284
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 7708 5188 8677 5216
rect 7708 5176 7714 5188
rect 8665 5185 8677 5188
rect 8711 5216 8723 5219
rect 9030 5216 9036 5228
rect 8711 5188 9036 5216
rect 8711 5185 8723 5188
rect 8665 5179 8723 5185
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 10778 5216 10784 5228
rect 10739 5188 10784 5216
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12492 5188 12817 5216
rect 12492 5176 12498 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5216 13507 5219
rect 14090 5216 14096 5228
rect 13495 5188 14096 5216
rect 13495 5185 13507 5188
rect 13449 5179 13507 5185
rect 14090 5176 14096 5188
rect 14148 5216 14154 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 14148 5188 14381 5216
rect 14148 5176 14154 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5216 15071 5219
rect 15378 5216 15384 5228
rect 15059 5188 15384 5216
rect 15059 5185 15071 5188
rect 15013 5179 15071 5185
rect 15378 5176 15384 5188
rect 15436 5216 15442 5228
rect 18800 5225 18828 5256
rect 19797 5253 19809 5256
rect 19843 5284 19855 5287
rect 24762 5284 24768 5296
rect 19843 5256 24768 5284
rect 19843 5253 19855 5256
rect 19797 5247 19855 5253
rect 16209 5219 16267 5225
rect 16209 5216 16221 5219
rect 15436 5188 16221 5216
rect 15436 5176 15442 5188
rect 16209 5185 16221 5188
rect 16255 5185 16267 5219
rect 16209 5179 16267 5185
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 19150 5216 19156 5228
rect 19111 5188 19156 5216
rect 18785 5179 18843 5185
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 24504 5225 24532 5256
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 24489 5219 24547 5225
rect 24489 5185 24501 5219
rect 24535 5185 24547 5219
rect 24489 5179 24547 5185
rect 106 5108 112 5160
rect 164 5148 170 5160
rect 1432 5151 1490 5157
rect 1432 5148 1444 5151
rect 164 5120 1444 5148
rect 164 5108 170 5120
rect 1432 5117 1444 5120
rect 1478 5148 1490 5151
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1478 5120 1869 5148
rect 1478 5117 1490 5120
rect 1432 5111 1490 5117
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 8938 5080 8944 5092
rect 8896 5052 8944 5080
rect 8938 5040 8944 5052
rect 8996 5089 9002 5092
rect 8996 5083 9044 5089
rect 8996 5049 8998 5083
rect 9032 5049 9044 5083
rect 8996 5043 9044 5049
rect 8996 5040 9029 5043
rect 10042 5040 10048 5092
rect 10100 5080 10106 5092
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 10100 5052 10517 5080
rect 10100 5040 10106 5052
rect 10505 5049 10517 5052
rect 10551 5049 10563 5083
rect 10505 5043 10563 5049
rect 10597 5083 10655 5089
rect 10597 5049 10609 5083
rect 10643 5049 10655 5083
rect 10597 5043 10655 5049
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12618 5080 12624 5092
rect 11931 5052 12624 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 1535 5015 1593 5021
rect 1535 4981 1547 5015
rect 1581 5012 1593 5015
rect 2130 5012 2136 5024
rect 1581 4984 2136 5012
rect 1581 4981 1593 4984
rect 1535 4975 1593 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 8481 5015 8539 5021
rect 8481 5012 8493 5015
rect 3476 4984 8493 5012
rect 3476 4972 3482 4984
rect 8481 4981 8493 4984
rect 8527 5012 8539 5015
rect 9001 5012 9029 5040
rect 9582 5012 9588 5024
rect 8527 4984 9029 5012
rect 9543 4984 9588 5012
rect 8527 4981 8539 4984
rect 8481 4975 8539 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 10192 4984 10241 5012
rect 10192 4972 10198 4984
rect 10229 4981 10241 4984
rect 10275 5012 10287 5015
rect 10612 5012 10640 5043
rect 12618 5040 12624 5052
rect 12676 5080 12682 5092
rect 12874 5083 12932 5089
rect 12874 5080 12886 5083
rect 12676 5052 12886 5080
rect 12676 5040 12682 5052
rect 12874 5049 12886 5052
rect 12920 5049 12932 5083
rect 12874 5043 12932 5049
rect 14458 5040 14464 5092
rect 14516 5080 14522 5092
rect 15930 5080 15936 5092
rect 14516 5052 14561 5080
rect 15891 5052 15936 5080
rect 14516 5040 14522 5052
rect 15930 5040 15936 5052
rect 15988 5040 15994 5092
rect 16025 5083 16083 5089
rect 16025 5049 16037 5083
rect 16071 5049 16083 5083
rect 16025 5043 16083 5049
rect 11514 5012 11520 5024
rect 10275 4984 10640 5012
rect 11475 4984 11520 5012
rect 10275 4981 10287 4984
rect 10229 4975 10287 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 15654 5012 15660 5024
rect 15615 4984 15660 5012
rect 15654 4972 15660 4984
rect 15712 5012 15718 5024
rect 16040 5012 16068 5043
rect 18230 5040 18236 5092
rect 18288 5080 18294 5092
rect 18877 5083 18935 5089
rect 18877 5080 18889 5083
rect 18288 5052 18889 5080
rect 18288 5040 18294 5052
rect 18877 5049 18889 5052
rect 18923 5049 18935 5083
rect 24210 5080 24216 5092
rect 24171 5052 24216 5080
rect 18877 5043 18935 5049
rect 24210 5040 24216 5052
rect 24268 5040 24274 5092
rect 24305 5083 24363 5089
rect 24305 5049 24317 5083
rect 24351 5049 24363 5083
rect 24305 5043 24363 5049
rect 18598 5012 18604 5024
rect 15712 4984 16068 5012
rect 18559 4984 18604 5012
rect 15712 4972 15718 4984
rect 18598 4972 18604 4984
rect 18656 4972 18662 5024
rect 24026 4972 24032 5024
rect 24084 5012 24090 5024
rect 24320 5012 24348 5043
rect 24084 4984 24348 5012
rect 24084 4972 24090 4984
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 10042 4808 10048 4820
rect 8619 4780 10048 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 10042 4768 10048 4780
rect 10100 4808 10106 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10100 4780 10701 4808
rect 10100 4768 10106 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 10689 4771 10747 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 18598 4808 18604 4820
rect 18559 4780 18604 4808
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 18690 4768 18696 4820
rect 18748 4808 18754 4820
rect 22879 4811 22937 4817
rect 22879 4808 22891 4811
rect 18748 4780 22891 4808
rect 18748 4768 18754 4780
rect 22879 4777 22891 4780
rect 22925 4777 22937 4811
rect 24210 4808 24216 4820
rect 24171 4780 24216 4808
rect 22879 4771 22937 4777
rect 24210 4768 24216 4780
rect 24268 4808 24274 4820
rect 24719 4811 24777 4817
rect 24719 4808 24731 4811
rect 24268 4780 24731 4808
rect 24268 4768 24274 4780
rect 24719 4777 24731 4780
rect 24765 4777 24777 4811
rect 24719 4771 24777 4777
rect 9030 4740 9036 4752
rect 8991 4712 9036 4740
rect 9030 4700 9036 4712
rect 9088 4700 9094 4752
rect 9582 4700 9588 4752
rect 9640 4740 9646 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9640 4712 9873 4740
rect 9640 4700 9646 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 9861 4703 9919 4709
rect 10413 4743 10471 4749
rect 10413 4709 10425 4743
rect 10459 4740 10471 4743
rect 10778 4740 10784 4752
rect 10459 4712 10784 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 12618 4740 12624 4752
rect 12579 4712 12624 4740
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 14185 4743 14243 4749
rect 14185 4709 14197 4743
rect 14231 4740 14243 4743
rect 15841 4743 15899 4749
rect 15841 4740 15853 4743
rect 14231 4712 15853 4740
rect 14231 4709 14243 4712
rect 14185 4703 14243 4709
rect 15841 4709 15853 4712
rect 15887 4740 15899 4743
rect 15930 4740 15936 4752
rect 15887 4712 15936 4740
rect 15887 4709 15899 4712
rect 15841 4703 15899 4709
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 12710 4672 12716 4684
rect 12671 4644 12716 4672
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4672 15255 4675
rect 15378 4672 15384 4684
rect 15243 4644 15384 4672
rect 15243 4641 15255 4644
rect 15197 4635 15255 4641
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 18230 4672 18236 4684
rect 18191 4644 18236 4672
rect 18230 4632 18236 4644
rect 18288 4672 18294 4684
rect 19153 4675 19211 4681
rect 19153 4672 19165 4675
rect 18288 4644 19165 4672
rect 18288 4632 18294 4644
rect 19153 4641 19165 4644
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 22808 4675 22866 4681
rect 22808 4641 22820 4675
rect 22854 4672 22866 4675
rect 22922 4672 22928 4684
rect 22854 4644 22928 4672
rect 22854 4641 22866 4644
rect 22808 4635 22866 4641
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 24670 4681 24676 4684
rect 24648 4675 24676 4681
rect 24648 4672 24660 4675
rect 24583 4644 24660 4672
rect 24648 4641 24660 4644
rect 24728 4672 24734 4684
rect 27614 4672 27620 4684
rect 24728 4644 27620 4672
rect 24648 4635 24676 4641
rect 24670 4632 24676 4635
rect 24728 4632 24734 4644
rect 27614 4632 27620 4644
rect 27672 4632 27678 4684
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 9858 4604 9864 4616
rect 9815 4576 9864 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 9858 4564 9864 4576
rect 9916 4604 9922 4616
rect 10410 4604 10416 4616
rect 9916 4576 10416 4604
rect 9916 4564 9922 4576
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 15427 4471 15485 4477
rect 15427 4437 15439 4471
rect 15473 4468 15485 4471
rect 15746 4468 15752 4480
rect 15473 4440 15752 4468
rect 15473 4437 15485 4440
rect 15427 4431 15485 4437
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1210 4224 1216 4276
rect 1268 4264 1274 4276
rect 1535 4267 1593 4273
rect 1535 4264 1547 4267
rect 1268 4236 1547 4264
rect 1268 4224 1274 4236
rect 1535 4233 1547 4236
rect 1581 4233 1593 4267
rect 1535 4227 1593 4233
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 10045 4267 10103 4273
rect 10045 4264 10057 4267
rect 9732 4236 10057 4264
rect 9732 4224 9738 4236
rect 10045 4233 10057 4236
rect 10091 4233 10103 4267
rect 10410 4264 10416 4276
rect 10371 4236 10416 4264
rect 10045 4227 10103 4233
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 12710 4264 12716 4276
rect 12671 4236 12716 4264
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 13630 4264 13636 4276
rect 13591 4236 13636 4264
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 15378 4264 15384 4276
rect 15339 4236 15384 4264
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 18230 4264 18236 4276
rect 18191 4236 18236 4264
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 19150 4224 19156 4276
rect 19208 4264 19214 4276
rect 19245 4267 19303 4273
rect 19245 4264 19257 4267
rect 19208 4236 19257 4264
rect 19208 4224 19214 4236
rect 19245 4233 19257 4236
rect 19291 4233 19303 4267
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 19245 4227 19303 4233
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 15654 4128 15660 4140
rect 14599 4100 15660 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 22830 4128 22836 4140
rect 22791 4100 22836 4128
rect 22830 4088 22836 4100
rect 22888 4088 22894 4140
rect 106 4020 112 4072
rect 164 4060 170 4072
rect 1432 4063 1490 4069
rect 1432 4060 1444 4063
rect 164 4032 1444 4060
rect 164 4020 170 4032
rect 1432 4029 1444 4032
rect 1478 4060 1490 4063
rect 1857 4063 1915 4069
rect 1857 4060 1869 4063
rect 1478 4032 1869 4060
rect 1478 4029 1490 4032
rect 1432 4023 1490 4029
rect 1857 4029 1869 4032
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4060 8999 4063
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8987 4032 9137 4060
rect 8987 4029 8999 4032
rect 8941 4023 8999 4029
rect 9125 4029 9137 4032
rect 9171 4060 9183 4063
rect 9582 4060 9588 4072
rect 9171 4032 9588 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13688 4032 13921 4060
rect 13688 4020 13694 4032
rect 13909 4029 13921 4032
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 18852 4063 18910 4069
rect 18852 4029 18864 4063
rect 18898 4060 18910 4063
rect 19150 4060 19156 4072
rect 18898 4032 19156 4060
rect 18898 4029 18910 4032
rect 18852 4023 18910 4029
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 9769 3995 9827 4001
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 10134 3992 10140 4004
rect 9815 3964 10140 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 18923 3927 18981 3933
rect 18923 3893 18935 3927
rect 18969 3924 18981 3927
rect 19150 3924 19156 3936
rect 18969 3896 19156 3924
rect 18969 3893 18981 3896
rect 18923 3887 18981 3893
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 22830 3884 22836 3936
rect 22888 3924 22894 3936
rect 24762 3924 24768 3936
rect 22888 3896 24768 3924
rect 22888 3884 22894 3896
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 9728 3587 9786 3593
rect 9728 3553 9740 3587
rect 9774 3584 9786 3587
rect 9950 3584 9956 3596
rect 9774 3556 9956 3584
rect 9774 3553 9786 3556
rect 9728 3547 9786 3553
rect 8496 3516 8524 3547
rect 9950 3544 9956 3556
rect 10008 3584 10014 3596
rect 10778 3584 10784 3596
rect 10008 3556 10784 3584
rect 10008 3544 10014 3556
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 16206 3584 16212 3596
rect 15804 3556 16212 3584
rect 15804 3544 15810 3556
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 19150 3584 19156 3596
rect 19111 3556 19156 3584
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 8570 3516 8576 3528
rect 8483 3488 8576 3516
rect 8570 3476 8576 3488
rect 8628 3516 8634 3528
rect 9815 3519 9873 3525
rect 9815 3516 9827 3519
rect 8628 3488 9827 3516
rect 8628 3476 8634 3488
rect 9815 3485 9827 3488
rect 9861 3485 9873 3519
rect 9815 3479 9873 3485
rect 8665 3383 8723 3389
rect 8665 3349 8677 3383
rect 8711 3380 8723 3383
rect 9674 3380 9680 3392
rect 8711 3352 9680 3380
rect 8711 3349 8723 3352
rect 8665 3343 8723 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 16393 3383 16451 3389
rect 16393 3349 16405 3383
rect 16439 3380 16451 3383
rect 18322 3380 18328 3392
rect 16439 3352 18328 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 19337 3383 19395 3389
rect 19337 3349 19349 3383
rect 19383 3380 19395 3383
rect 20162 3380 20168 3392
rect 19383 3352 20168 3380
rect 19383 3349 19395 3352
rect 19337 3343 19395 3349
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 8570 3176 8576 3188
rect 8531 3148 8576 3176
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 9769 3179 9827 3185
rect 9769 3145 9781 3179
rect 9815 3176 9827 3179
rect 9950 3176 9956 3188
rect 9815 3148 9956 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 16206 3176 16212 3188
rect 16167 3148 16212 3176
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 19150 3176 19156 3188
rect 19111 3148 19156 3176
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 12897 2635 12955 2641
rect 12897 2632 12909 2635
rect 12860 2604 12909 2632
rect 12860 2592 12866 2604
rect 12897 2601 12909 2604
rect 12943 2601 12955 2635
rect 12897 2595 12955 2601
rect 15703 2635 15761 2641
rect 15703 2601 15715 2635
rect 15749 2632 15761 2635
rect 16298 2632 16304 2644
rect 15749 2604 16304 2632
rect 15749 2601 15761 2604
rect 15703 2595 15761 2601
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 24719 2635 24777 2641
rect 24719 2601 24731 2635
rect 24765 2632 24777 2635
rect 24854 2632 24860 2644
rect 24765 2604 24860 2632
rect 24765 2601 24777 2604
rect 24719 2595 24777 2601
rect 24854 2592 24860 2604
rect 24912 2592 24918 2644
rect 7834 2524 7840 2576
rect 7892 2564 7898 2576
rect 14231 2567 14289 2573
rect 14231 2564 14243 2567
rect 7892 2536 14243 2564
rect 7892 2524 7898 2536
rect 14231 2533 14243 2536
rect 14277 2533 14289 2567
rect 14231 2527 14289 2533
rect 10042 2456 10048 2508
rect 10100 2496 10106 2508
rect 10505 2499 10563 2505
rect 10505 2496 10517 2499
rect 10100 2468 10517 2496
rect 10100 2456 10106 2468
rect 10505 2465 10517 2468
rect 10551 2496 10563 2499
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 10551 2468 11069 2496
rect 10551 2465 10563 2468
rect 10505 2459 10563 2465
rect 11057 2465 11069 2468
rect 11103 2465 11115 2499
rect 11057 2459 11115 2465
rect 12688 2499 12746 2505
rect 12688 2465 12700 2499
rect 12734 2496 12746 2499
rect 14144 2499 14202 2505
rect 12734 2468 13216 2496
rect 12734 2465 12746 2468
rect 12688 2459 12746 2465
rect 10689 2363 10747 2369
rect 10689 2329 10701 2363
rect 10735 2360 10747 2363
rect 11422 2360 11428 2372
rect 10735 2332 11428 2360
rect 10735 2329 10747 2332
rect 10689 2323 10747 2329
rect 11422 2320 11428 2332
rect 11480 2320 11486 2372
rect 13188 2301 13216 2468
rect 14144 2465 14156 2499
rect 14190 2496 14202 2499
rect 15632 2499 15690 2505
rect 14190 2468 14688 2496
rect 14190 2465 14202 2468
rect 14144 2459 14202 2465
rect 13173 2295 13231 2301
rect 13173 2261 13185 2295
rect 13219 2292 13231 2295
rect 13722 2292 13728 2304
rect 13219 2264 13728 2292
rect 13219 2261 13231 2264
rect 13173 2255 13231 2261
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14660 2301 14688 2468
rect 15632 2465 15644 2499
rect 15678 2496 15690 2499
rect 24648 2499 24706 2505
rect 15678 2468 16160 2496
rect 15678 2465 15690 2468
rect 15632 2459 15690 2465
rect 14645 2295 14703 2301
rect 14645 2261 14657 2295
rect 14691 2292 14703 2295
rect 15654 2292 15660 2304
rect 14691 2264 15660 2292
rect 14691 2261 14703 2264
rect 14645 2255 14703 2261
rect 15654 2252 15660 2264
rect 15712 2252 15718 2304
rect 16132 2301 16160 2468
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 24694 2468 25176 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 16117 2295 16175 2301
rect 16117 2261 16129 2295
rect 16163 2292 16175 2295
rect 22094 2292 22100 2304
rect 16163 2264 22100 2292
rect 16163 2261 16175 2264
rect 16117 2255 16175 2261
rect 22094 2252 22100 2264
rect 22152 2252 22158 2304
rect 25148 2301 25176 2468
rect 25133 2295 25191 2301
rect 25133 2261 25145 2295
rect 25179 2292 25191 2295
rect 26510 2292 26516 2304
rect 25179 2264 26516 2292
rect 25179 2261 25191 2264
rect 25133 2255 25191 2261
rect 26510 2252 26516 2264
rect 26568 2252 26574 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 13084 24352 13136 24404
rect 2228 24216 2280 24268
rect 9404 24216 9456 24268
rect 10784 24259 10836 24268
rect 10784 24225 10793 24259
rect 10793 24225 10827 24259
rect 10827 24225 10836 24259
rect 10784 24216 10836 24225
rect 16488 24259 16540 24268
rect 16488 24225 16506 24259
rect 16506 24225 16540 24259
rect 16488 24216 16540 24225
rect 18328 24216 18380 24268
rect 25136 24216 25188 24268
rect 3424 24012 3476 24064
rect 8392 24055 8444 24064
rect 8392 24021 8401 24055
rect 8401 24021 8435 24055
rect 8435 24021 8444 24055
rect 8392 24012 8444 24021
rect 9220 24012 9272 24064
rect 10048 24055 10100 24064
rect 10048 24021 10057 24055
rect 10057 24021 10091 24055
rect 10091 24021 10100 24055
rect 10048 24012 10100 24021
rect 14280 24012 14332 24064
rect 19984 24012 20036 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2228 23851 2280 23860
rect 2228 23817 2237 23851
rect 2237 23817 2271 23851
rect 2271 23817 2280 23851
rect 2228 23808 2280 23817
rect 4252 23851 4304 23860
rect 4252 23817 4261 23851
rect 4261 23817 4295 23851
rect 4295 23817 4304 23851
rect 4252 23808 4304 23817
rect 9404 23851 9456 23860
rect 9404 23817 9413 23851
rect 9413 23817 9447 23851
rect 9447 23817 9456 23851
rect 9404 23808 9456 23817
rect 10784 23808 10836 23860
rect 10968 23851 11020 23860
rect 10968 23817 10977 23851
rect 10977 23817 11011 23851
rect 11011 23817 11020 23851
rect 10968 23808 11020 23817
rect 14832 23808 14884 23860
rect 848 23604 900 23656
rect 4252 23604 4304 23656
rect 5448 23604 5500 23656
rect 3700 23468 3752 23520
rect 4436 23536 4488 23588
rect 4712 23579 4764 23588
rect 4712 23545 4721 23579
rect 4721 23545 4755 23579
rect 4755 23545 4764 23579
rect 4712 23536 4764 23545
rect 6460 23468 6512 23520
rect 8392 23604 8444 23656
rect 8760 23647 8812 23656
rect 8760 23613 8769 23647
rect 8769 23613 8803 23647
rect 8803 23613 8812 23647
rect 8760 23604 8812 23613
rect 9680 23604 9732 23656
rect 10048 23604 10100 23656
rect 11980 23604 12032 23656
rect 16580 23808 16632 23860
rect 16488 23783 16540 23792
rect 16488 23749 16497 23783
rect 16497 23749 16531 23783
rect 16531 23749 16540 23783
rect 16488 23740 16540 23749
rect 17224 23647 17276 23656
rect 8576 23511 8628 23520
rect 8576 23477 8585 23511
rect 8585 23477 8619 23511
rect 8619 23477 8628 23511
rect 8576 23468 8628 23477
rect 10048 23511 10100 23520
rect 10048 23477 10057 23511
rect 10057 23477 10091 23511
rect 10091 23477 10100 23511
rect 10048 23468 10100 23477
rect 17224 23613 17233 23647
rect 17233 23613 17267 23647
rect 17267 23613 17276 23647
rect 17224 23604 17276 23613
rect 21824 23808 21876 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 27068 23808 27120 23860
rect 25504 23783 25556 23792
rect 25504 23749 25513 23783
rect 25513 23749 25547 23783
rect 25547 23749 25556 23783
rect 25504 23740 25556 23749
rect 14648 23536 14700 23588
rect 16304 23536 16356 23588
rect 16948 23536 17000 23588
rect 16028 23468 16080 23520
rect 23296 23468 23348 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 10968 23264 11020 23316
rect 15936 23264 15988 23316
rect 16948 23264 17000 23316
rect 13728 23239 13780 23248
rect 13728 23205 13737 23239
rect 13737 23205 13771 23239
rect 13771 23205 13780 23239
rect 13728 23196 13780 23205
rect 1032 23128 1084 23180
rect 1584 23128 1636 23180
rect 2596 23128 2648 23180
rect 5356 23171 5408 23180
rect 5356 23137 5365 23171
rect 5365 23137 5399 23171
rect 5399 23137 5408 23171
rect 5356 23128 5408 23137
rect 8208 23171 8260 23180
rect 8208 23137 8217 23171
rect 8217 23137 8251 23171
rect 8251 23137 8260 23171
rect 8208 23128 8260 23137
rect 9588 23171 9640 23180
rect 9588 23137 9597 23171
rect 9597 23137 9631 23171
rect 9631 23137 9640 23171
rect 9588 23128 9640 23137
rect 11336 23171 11388 23180
rect 11336 23137 11345 23171
rect 11345 23137 11379 23171
rect 11379 23137 11388 23171
rect 11336 23128 11388 23137
rect 15476 23128 15528 23180
rect 24676 23128 24728 23180
rect 14556 23103 14608 23112
rect 14556 23069 14565 23103
rect 14565 23069 14599 23103
rect 14599 23069 14608 23103
rect 14556 23060 14608 23069
rect 16212 22992 16264 23044
rect 1860 22924 1912 22976
rect 2320 22924 2372 22976
rect 4620 22967 4672 22976
rect 4620 22933 4629 22967
rect 4629 22933 4663 22967
rect 4663 22933 4672 22967
rect 4620 22924 4672 22933
rect 5172 22967 5224 22976
rect 5172 22933 5181 22967
rect 5181 22933 5215 22967
rect 5215 22933 5224 22967
rect 5172 22924 5224 22933
rect 8300 22967 8352 22976
rect 8300 22933 8309 22967
rect 8309 22933 8343 22967
rect 8343 22933 8352 22967
rect 8300 22924 8352 22933
rect 11520 22967 11572 22976
rect 11520 22933 11529 22967
rect 11529 22933 11563 22967
rect 11563 22933 11572 22967
rect 11520 22924 11572 22933
rect 13544 22924 13596 22976
rect 15384 22924 15436 22976
rect 15752 22924 15804 22976
rect 22100 22924 22152 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 2596 22720 2648 22772
rect 8208 22763 8260 22772
rect 8208 22729 8217 22763
rect 8217 22729 8251 22763
rect 8251 22729 8260 22763
rect 8208 22720 8260 22729
rect 11336 22763 11388 22772
rect 11336 22729 11345 22763
rect 11345 22729 11379 22763
rect 11379 22729 11388 22763
rect 11336 22720 11388 22729
rect 15476 22763 15528 22772
rect 15476 22729 15485 22763
rect 15485 22729 15519 22763
rect 15519 22729 15528 22763
rect 15476 22720 15528 22729
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 2320 22559 2372 22568
rect 2320 22525 2329 22559
rect 2329 22525 2363 22559
rect 2363 22525 2372 22559
rect 2320 22516 2372 22525
rect 3332 22516 3384 22568
rect 4712 22491 4764 22500
rect 4712 22457 4721 22491
rect 4721 22457 4755 22491
rect 4755 22457 4764 22491
rect 4712 22448 4764 22457
rect 5264 22491 5316 22500
rect 5264 22457 5273 22491
rect 5273 22457 5307 22491
rect 5307 22457 5316 22491
rect 5264 22448 5316 22457
rect 8668 22584 8720 22636
rect 9588 22584 9640 22636
rect 8852 22491 8904 22500
rect 8852 22457 8861 22491
rect 8861 22457 8895 22491
rect 8895 22457 8904 22491
rect 8852 22448 8904 22457
rect 2228 22423 2280 22432
rect 2228 22389 2237 22423
rect 2237 22389 2271 22423
rect 2271 22389 2280 22423
rect 2228 22380 2280 22389
rect 5356 22380 5408 22432
rect 7564 22380 7616 22432
rect 9588 22448 9640 22500
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 12808 22516 12860 22568
rect 13912 22652 13964 22704
rect 13728 22627 13780 22636
rect 13728 22593 13737 22627
rect 13737 22593 13771 22627
rect 13771 22593 13780 22627
rect 13728 22584 13780 22593
rect 14556 22584 14608 22636
rect 15016 22491 15068 22500
rect 14096 22423 14148 22432
rect 10140 22380 10192 22389
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 15016 22457 15025 22491
rect 15025 22457 15059 22491
rect 15059 22457 15068 22491
rect 15016 22448 15068 22457
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 16212 22627 16264 22636
rect 16212 22593 16221 22627
rect 16221 22593 16255 22627
rect 16255 22593 16264 22627
rect 16212 22584 16264 22593
rect 20076 22720 20128 22772
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 15752 22448 15804 22500
rect 14096 22380 14148 22389
rect 15844 22380 15896 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5264 22176 5316 22228
rect 2228 22108 2280 22160
rect 5448 22151 5500 22160
rect 5448 22117 5457 22151
rect 5457 22117 5491 22151
rect 5491 22117 5500 22151
rect 5448 22108 5500 22117
rect 8852 22176 8904 22228
rect 9496 22176 9548 22228
rect 8300 22108 8352 22160
rect 9220 22108 9272 22160
rect 9772 22151 9824 22160
rect 9772 22117 9781 22151
rect 9781 22117 9815 22151
rect 9815 22117 9824 22151
rect 9772 22108 9824 22117
rect 10140 22176 10192 22228
rect 12808 22219 12860 22228
rect 12808 22185 12817 22219
rect 12817 22185 12851 22219
rect 12851 22185 12860 22219
rect 12808 22176 12860 22185
rect 13544 22219 13596 22228
rect 13544 22185 13553 22219
rect 13553 22185 13587 22219
rect 13587 22185 13596 22219
rect 13544 22176 13596 22185
rect 14096 22219 14148 22228
rect 14096 22185 14105 22219
rect 14105 22185 14139 22219
rect 14139 22185 14148 22219
rect 14096 22176 14148 22185
rect 15016 22176 15068 22228
rect 15752 22176 15804 22228
rect 11520 22108 11572 22160
rect 15384 22151 15436 22160
rect 15384 22117 15393 22151
rect 15393 22117 15427 22151
rect 15427 22117 15436 22151
rect 15384 22108 15436 22117
rect 15476 22151 15528 22160
rect 15476 22117 15485 22151
rect 15485 22117 15519 22151
rect 15519 22117 15528 22151
rect 15476 22108 15528 22117
rect 7104 22040 7156 22092
rect 1216 21972 1268 22024
rect 3516 21972 3568 22024
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 6184 21972 6236 22024
rect 7564 21972 7616 22024
rect 9588 21972 9640 22024
rect 11796 21972 11848 22024
rect 2780 21904 2832 21956
rect 7840 21947 7892 21956
rect 7840 21913 7849 21947
rect 7849 21913 7883 21947
rect 7883 21913 7892 21947
rect 7840 21904 7892 21913
rect 8668 21947 8720 21956
rect 8668 21913 8677 21947
rect 8677 21913 8711 21947
rect 8711 21913 8720 21947
rect 8668 21904 8720 21913
rect 12256 21904 12308 21956
rect 13728 21972 13780 22024
rect 24676 22040 24728 22092
rect 14464 21972 14516 22024
rect 15476 21972 15528 22024
rect 15844 21904 15896 21956
rect 4344 21836 4396 21888
rect 5540 21836 5592 21888
rect 6828 21836 6880 21888
rect 10876 21879 10928 21888
rect 10876 21845 10885 21879
rect 10885 21845 10919 21879
rect 10919 21845 10928 21879
rect 10876 21836 10928 21845
rect 18604 21836 18656 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2228 21632 2280 21684
rect 3516 21675 3568 21684
rect 3516 21641 3525 21675
rect 3525 21641 3559 21675
rect 3559 21641 3568 21675
rect 3516 21632 3568 21641
rect 3884 21675 3936 21684
rect 3884 21641 3893 21675
rect 3893 21641 3927 21675
rect 3927 21641 3936 21675
rect 3884 21632 3936 21641
rect 5448 21632 5500 21684
rect 7656 21632 7708 21684
rect 8300 21632 8352 21684
rect 2780 21607 2832 21616
rect 2780 21573 2789 21607
rect 2789 21573 2823 21607
rect 2823 21573 2832 21607
rect 2780 21564 2832 21573
rect 7564 21607 7616 21616
rect 7564 21573 7573 21607
rect 7573 21573 7607 21607
rect 7607 21573 7616 21607
rect 7564 21564 7616 21573
rect 8668 21607 8720 21616
rect 8668 21573 8677 21607
rect 8677 21573 8711 21607
rect 8711 21573 8720 21607
rect 8668 21564 8720 21573
rect 11060 21632 11112 21684
rect 11520 21632 11572 21684
rect 13728 21675 13780 21684
rect 13728 21641 13737 21675
rect 13737 21641 13771 21675
rect 13771 21641 13780 21675
rect 13728 21632 13780 21641
rect 15384 21632 15436 21684
rect 15476 21632 15528 21684
rect 16028 21632 16080 21684
rect 24676 21675 24728 21684
rect 24676 21641 24685 21675
rect 24685 21641 24719 21675
rect 24719 21641 24728 21675
rect 24676 21632 24728 21641
rect 1860 21496 1912 21548
rect 5264 21496 5316 21548
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 7840 21496 7892 21548
rect 3700 21471 3752 21480
rect 3700 21437 3709 21471
rect 3709 21437 3743 21471
rect 3743 21437 3752 21471
rect 3700 21428 3752 21437
rect 6828 21471 6880 21480
rect 6828 21437 6837 21471
rect 6837 21437 6871 21471
rect 6871 21437 6880 21471
rect 6828 21428 6880 21437
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 2320 21403 2372 21412
rect 2320 21369 2329 21403
rect 2329 21369 2363 21403
rect 2363 21369 2372 21403
rect 2320 21360 2372 21369
rect 3332 21360 3384 21412
rect 5264 21403 5316 21412
rect 5264 21369 5273 21403
rect 5273 21369 5307 21403
rect 5307 21369 5316 21403
rect 5264 21360 5316 21369
rect 8208 21403 8260 21412
rect 8208 21369 8217 21403
rect 8217 21369 8251 21403
rect 8251 21369 8260 21403
rect 8208 21360 8260 21369
rect 11336 21360 11388 21412
rect 12256 21360 12308 21412
rect 12900 21471 12952 21480
rect 12900 21437 12909 21471
rect 12909 21437 12943 21471
rect 12943 21437 12952 21471
rect 12900 21428 12952 21437
rect 14832 21360 14884 21412
rect 15660 21403 15712 21412
rect 7104 21292 7156 21344
rect 9496 21292 9548 21344
rect 12348 21292 12400 21344
rect 12532 21335 12584 21344
rect 12532 21301 12541 21335
rect 12541 21301 12575 21335
rect 12575 21301 12584 21335
rect 12532 21292 12584 21301
rect 15660 21369 15669 21403
rect 15669 21369 15703 21403
rect 15703 21369 15712 21403
rect 15660 21360 15712 21369
rect 15568 21292 15620 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5448 21088 5500 21140
rect 6828 21088 6880 21140
rect 7932 21131 7984 21140
rect 7932 21097 7941 21131
rect 7941 21097 7975 21131
rect 7975 21097 7984 21131
rect 7932 21088 7984 21097
rect 8208 21088 8260 21140
rect 8576 21088 8628 21140
rect 9772 21088 9824 21140
rect 11336 21088 11388 21140
rect 11796 21131 11848 21140
rect 11796 21097 11805 21131
rect 11805 21097 11839 21131
rect 11839 21097 11848 21131
rect 11796 21088 11848 21097
rect 13912 21131 13964 21140
rect 13912 21097 13921 21131
rect 13921 21097 13955 21131
rect 13955 21097 13964 21131
rect 13912 21088 13964 21097
rect 2044 21063 2096 21072
rect 2044 21029 2053 21063
rect 2053 21029 2087 21063
rect 2087 21029 2096 21063
rect 2044 21020 2096 21029
rect 5356 21020 5408 21072
rect 10600 21020 10652 21072
rect 13452 21020 13504 21072
rect 15476 21063 15528 21072
rect 15476 21029 15485 21063
rect 15485 21029 15519 21063
rect 15519 21029 15528 21063
rect 15476 21020 15528 21029
rect 15568 21020 15620 21072
rect 2964 20995 3016 21004
rect 2964 20961 2973 20995
rect 2973 20961 3007 20995
rect 3007 20961 3016 20995
rect 2964 20952 3016 20961
rect 8484 20952 8536 21004
rect 10232 20952 10284 21004
rect 12532 20952 12584 21004
rect 17224 20952 17276 21004
rect 1952 20927 2004 20936
rect 1952 20893 1961 20927
rect 1961 20893 1995 20927
rect 1995 20893 2004 20927
rect 1952 20884 2004 20893
rect 2596 20927 2648 20936
rect 2596 20893 2605 20927
rect 2605 20893 2639 20927
rect 2639 20893 2648 20927
rect 2596 20884 2648 20893
rect 4896 20927 4948 20936
rect 4896 20893 4905 20927
rect 4905 20893 4939 20927
rect 4939 20893 4948 20927
rect 4896 20884 4948 20893
rect 7564 20927 7616 20936
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 12992 20927 13044 20936
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 15384 20927 15436 20936
rect 15384 20893 15393 20927
rect 15393 20893 15427 20927
rect 15427 20893 15436 20927
rect 15384 20884 15436 20893
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 1676 20791 1728 20800
rect 1676 20757 1685 20791
rect 1685 20757 1719 20791
rect 1719 20757 1728 20791
rect 1676 20748 1728 20757
rect 5540 20748 5592 20800
rect 6184 20791 6236 20800
rect 6184 20757 6193 20791
rect 6193 20757 6227 20791
rect 6227 20757 6236 20791
rect 6184 20748 6236 20757
rect 7472 20748 7524 20800
rect 11980 20748 12032 20800
rect 12900 20748 12952 20800
rect 14188 20748 14240 20800
rect 14832 20748 14884 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 3332 20587 3384 20596
rect 3332 20553 3341 20587
rect 3341 20553 3375 20587
rect 3375 20553 3384 20587
rect 3332 20544 3384 20553
rect 5264 20544 5316 20596
rect 9496 20587 9548 20596
rect 9496 20553 9505 20587
rect 9505 20553 9539 20587
rect 9539 20553 9548 20587
rect 9496 20544 9548 20553
rect 10232 20587 10284 20596
rect 10232 20553 10241 20587
rect 10241 20553 10275 20587
rect 10275 20553 10284 20587
rect 10232 20544 10284 20553
rect 14464 20587 14516 20596
rect 14464 20553 14473 20587
rect 14473 20553 14507 20587
rect 14507 20553 14516 20587
rect 14464 20544 14516 20553
rect 17224 20587 17276 20596
rect 17224 20553 17233 20587
rect 17233 20553 17267 20587
rect 17267 20553 17276 20587
rect 17224 20544 17276 20553
rect 4896 20476 4948 20528
rect 7932 20519 7984 20528
rect 7932 20485 7941 20519
rect 7941 20485 7975 20519
rect 7975 20485 7984 20519
rect 7932 20476 7984 20485
rect 2964 20408 3016 20460
rect 8576 20451 8628 20460
rect 8576 20417 8585 20451
rect 8585 20417 8619 20451
rect 8619 20417 8628 20451
rect 8576 20408 8628 20417
rect 1676 20340 1728 20392
rect 2044 20340 2096 20392
rect 4804 20340 4856 20392
rect 2412 20272 2464 20324
rect 1676 20247 1728 20256
rect 1676 20213 1685 20247
rect 1685 20213 1719 20247
rect 1719 20213 1728 20247
rect 1676 20204 1728 20213
rect 5356 20272 5408 20324
rect 7472 20340 7524 20392
rect 7932 20272 7984 20324
rect 10600 20476 10652 20528
rect 16304 20451 16356 20460
rect 16304 20417 16313 20451
rect 16313 20417 16347 20451
rect 16347 20417 16356 20451
rect 16304 20408 16356 20417
rect 11336 20340 11388 20392
rect 13360 20340 13412 20392
rect 10600 20315 10652 20324
rect 10600 20281 10609 20315
rect 10609 20281 10643 20315
rect 10643 20281 10652 20315
rect 10600 20272 10652 20281
rect 15384 20272 15436 20324
rect 10968 20247 11020 20256
rect 10968 20213 10977 20247
rect 10977 20213 11011 20247
rect 11011 20213 11020 20247
rect 10968 20204 11020 20213
rect 11060 20204 11112 20256
rect 13452 20247 13504 20256
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 14832 20204 14884 20256
rect 15476 20204 15528 20256
rect 16396 20315 16448 20324
rect 16396 20281 16405 20315
rect 16405 20281 16439 20315
rect 16439 20281 16448 20315
rect 16396 20272 16448 20281
rect 17592 20272 17644 20324
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 4896 20000 4948 20052
rect 7564 20043 7616 20052
rect 7564 20009 7573 20043
rect 7573 20009 7607 20043
rect 7607 20009 7616 20043
rect 7564 20000 7616 20009
rect 10048 20000 10100 20052
rect 2504 19932 2556 19984
rect 4252 19932 4304 19984
rect 4988 19975 5040 19984
rect 4988 19941 4997 19975
rect 4997 19941 5031 19975
rect 5031 19941 5040 19975
rect 4988 19932 5040 19941
rect 5172 19932 5224 19984
rect 6460 19907 6512 19916
rect 6460 19873 6469 19907
rect 6469 19873 6503 19907
rect 6503 19873 6512 19907
rect 6460 19864 6512 19873
rect 7472 19864 7524 19916
rect 8024 19907 8076 19916
rect 8024 19873 8033 19907
rect 8033 19873 8067 19907
rect 8067 19873 8076 19907
rect 8024 19864 8076 19873
rect 2320 19839 2372 19848
rect 2320 19805 2329 19839
rect 2329 19805 2363 19839
rect 2363 19805 2372 19839
rect 2320 19796 2372 19805
rect 2596 19839 2648 19848
rect 2596 19805 2605 19839
rect 2605 19805 2639 19839
rect 2639 19805 2648 19839
rect 2596 19796 2648 19805
rect 8852 19864 8904 19916
rect 10692 20000 10744 20052
rect 11336 20043 11388 20052
rect 11336 20009 11345 20043
rect 11345 20009 11379 20043
rect 11379 20009 11388 20043
rect 11336 20000 11388 20009
rect 12992 20000 13044 20052
rect 14188 20043 14240 20052
rect 14188 20009 14197 20043
rect 14197 20009 14231 20043
rect 14231 20009 14240 20043
rect 14188 20000 14240 20009
rect 15384 19932 15436 19984
rect 17132 19932 17184 19984
rect 18696 19907 18748 19916
rect 18696 19873 18705 19907
rect 18705 19873 18739 19907
rect 18739 19873 18748 19907
rect 18696 19864 18748 19873
rect 24676 19864 24728 19916
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 15292 19839 15344 19848
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 15292 19796 15344 19805
rect 17500 19796 17552 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 5540 19771 5592 19780
rect 5540 19737 5549 19771
rect 5549 19737 5583 19771
rect 5583 19737 5592 19771
rect 5540 19728 5592 19737
rect 1400 19660 1452 19712
rect 1952 19660 2004 19712
rect 3332 19703 3384 19712
rect 3332 19669 3341 19703
rect 3341 19669 3375 19703
rect 3375 19669 3384 19703
rect 3332 19660 3384 19669
rect 4436 19703 4488 19712
rect 4436 19669 4445 19703
rect 4445 19669 4479 19703
rect 4479 19669 4488 19703
rect 4436 19660 4488 19669
rect 13360 19660 13412 19712
rect 14004 19703 14056 19712
rect 14004 19669 14013 19703
rect 14013 19669 14047 19703
rect 14047 19669 14056 19703
rect 14004 19660 14056 19669
rect 16396 19660 16448 19712
rect 18696 19660 18748 19712
rect 23388 19660 23440 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 2412 19499 2464 19508
rect 2412 19465 2421 19499
rect 2421 19465 2455 19499
rect 2455 19465 2464 19499
rect 2412 19456 2464 19465
rect 5172 19456 5224 19508
rect 6460 19499 6512 19508
rect 6460 19465 6469 19499
rect 6469 19465 6503 19499
rect 6503 19465 6512 19499
rect 6460 19456 6512 19465
rect 4988 19388 5040 19440
rect 7472 19388 7524 19440
rect 10048 19456 10100 19508
rect 10692 19456 10744 19508
rect 11336 19456 11388 19508
rect 14832 19456 14884 19508
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 18696 19499 18748 19508
rect 18696 19465 18705 19499
rect 18705 19465 18739 19499
rect 18739 19465 18748 19499
rect 18696 19456 18748 19465
rect 24676 19499 24728 19508
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 2320 19320 2372 19372
rect 6828 19320 6880 19372
rect 1676 19252 1728 19304
rect 2228 19252 2280 19304
rect 13452 19388 13504 19440
rect 13912 19388 13964 19440
rect 11060 19320 11112 19372
rect 11704 19320 11756 19372
rect 12532 19320 12584 19372
rect 14004 19363 14056 19372
rect 14004 19329 14013 19363
rect 14013 19329 14047 19363
rect 14047 19329 14056 19363
rect 14004 19320 14056 19329
rect 15568 19320 15620 19372
rect 8852 19295 8904 19304
rect 8852 19261 8861 19295
rect 8861 19261 8895 19295
rect 8895 19261 8904 19295
rect 8852 19252 8904 19261
rect 12348 19252 12400 19304
rect 2504 19184 2556 19236
rect 3056 19184 3108 19236
rect 3332 19184 3384 19236
rect 4252 19184 4304 19236
rect 4436 19227 4488 19236
rect 4436 19193 4445 19227
rect 4445 19193 4479 19227
rect 4479 19193 4488 19227
rect 4436 19184 4488 19193
rect 3516 19159 3568 19168
rect 3516 19125 3525 19159
rect 3525 19125 3559 19159
rect 3559 19125 3568 19159
rect 3516 19116 3568 19125
rect 4160 19159 4212 19168
rect 4160 19125 4169 19159
rect 4169 19125 4203 19159
rect 4203 19125 4212 19159
rect 4804 19184 4856 19236
rect 7932 19159 7984 19168
rect 4160 19116 4212 19125
rect 7932 19125 7941 19159
rect 7941 19125 7975 19159
rect 7975 19125 7984 19159
rect 7932 19116 7984 19125
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 10968 19184 11020 19236
rect 12532 19184 12584 19236
rect 13728 19252 13780 19304
rect 13176 19227 13228 19236
rect 13176 19193 13185 19227
rect 13185 19193 13219 19227
rect 13219 19193 13228 19227
rect 13176 19184 13228 19193
rect 12992 19116 13044 19168
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 15384 19184 15436 19236
rect 15568 19227 15620 19236
rect 15568 19193 15577 19227
rect 15577 19193 15611 19227
rect 15611 19193 15620 19227
rect 15568 19184 15620 19193
rect 16304 19295 16356 19304
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 13912 19116 13964 19125
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2044 18844 2096 18896
rect 2228 18844 2280 18896
rect 4252 18844 4304 18896
rect 11060 18955 11112 18964
rect 11060 18921 11069 18955
rect 11069 18921 11103 18955
rect 11103 18921 11112 18955
rect 11060 18912 11112 18921
rect 12256 18912 12308 18964
rect 13176 18912 13228 18964
rect 15292 18912 15344 18964
rect 6552 18887 6604 18896
rect 6552 18853 6561 18887
rect 6561 18853 6595 18887
rect 6595 18853 6604 18887
rect 6552 18844 6604 18853
rect 6828 18844 6880 18896
rect 12532 18844 12584 18896
rect 13728 18887 13780 18896
rect 4160 18819 4212 18828
rect 4160 18785 4169 18819
rect 4169 18785 4203 18819
rect 4203 18785 4212 18819
rect 7932 18819 7984 18828
rect 4160 18776 4212 18785
rect 7932 18785 7941 18819
rect 7941 18785 7975 18819
rect 7975 18785 7984 18819
rect 7932 18776 7984 18785
rect 8024 18776 8076 18828
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 11704 18776 11756 18828
rect 12716 18776 12768 18828
rect 13728 18853 13737 18887
rect 13737 18853 13771 18887
rect 13771 18853 13780 18887
rect 13728 18844 13780 18853
rect 16120 18912 16172 18964
rect 15936 18844 15988 18896
rect 1860 18708 1912 18760
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 3424 18708 3476 18760
rect 5264 18708 5316 18760
rect 7104 18751 7156 18760
rect 1676 18683 1728 18692
rect 1676 18649 1685 18683
rect 1685 18649 1719 18683
rect 1719 18649 1728 18683
rect 1676 18640 1728 18649
rect 2596 18640 2648 18692
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 6000 18572 6052 18624
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 15752 18708 15804 18760
rect 16212 18708 16264 18760
rect 9864 18640 9916 18692
rect 10140 18572 10192 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 14832 18572 14884 18624
rect 16304 18572 16356 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2044 18411 2096 18420
rect 2044 18377 2053 18411
rect 2053 18377 2087 18411
rect 2087 18377 2096 18411
rect 2044 18368 2096 18377
rect 4068 18368 4120 18420
rect 4160 18368 4212 18420
rect 6092 18368 6144 18420
rect 7932 18411 7984 18420
rect 7932 18377 7941 18411
rect 7941 18377 7975 18411
rect 7975 18377 7984 18411
rect 7932 18368 7984 18377
rect 11704 18411 11756 18420
rect 11704 18377 11713 18411
rect 11713 18377 11747 18411
rect 11747 18377 11756 18411
rect 11704 18368 11756 18377
rect 3700 18300 3752 18352
rect 7104 18300 7156 18352
rect 9680 18300 9732 18352
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 8392 18232 8444 18284
rect 9588 18232 9640 18284
rect 10876 18232 10928 18284
rect 1676 18164 1728 18216
rect 2964 18164 3016 18216
rect 4804 18164 4856 18216
rect 7656 18164 7708 18216
rect 16120 18300 16172 18352
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14096 18232 14148 18241
rect 15936 18275 15988 18284
rect 15936 18241 15945 18275
rect 15945 18241 15979 18275
rect 15979 18241 15988 18275
rect 15936 18232 15988 18241
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 12716 18164 12768 18216
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 3056 18028 3108 18080
rect 5264 18096 5316 18148
rect 4068 18071 4120 18080
rect 4068 18037 4077 18071
rect 4077 18037 4111 18071
rect 4111 18037 4120 18071
rect 4068 18028 4120 18037
rect 6000 18096 6052 18148
rect 6368 18028 6420 18080
rect 10232 18139 10284 18148
rect 10232 18105 10241 18139
rect 10241 18105 10275 18139
rect 10275 18105 10284 18139
rect 10784 18139 10836 18148
rect 10232 18096 10284 18105
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 10784 18096 10836 18105
rect 13452 18096 13504 18148
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 12716 18028 12768 18080
rect 13820 18028 13872 18080
rect 15752 18071 15804 18080
rect 15752 18037 15761 18071
rect 15761 18037 15795 18071
rect 15795 18037 15804 18071
rect 15752 18028 15804 18037
rect 16120 18028 16172 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1400 17867 1452 17876
rect 1400 17833 1409 17867
rect 1409 17833 1443 17867
rect 1443 17833 1452 17867
rect 1400 17824 1452 17833
rect 6552 17824 6604 17876
rect 7656 17824 7708 17876
rect 8024 17867 8076 17876
rect 8024 17833 8033 17867
rect 8033 17833 8067 17867
rect 8067 17833 8076 17867
rect 8024 17824 8076 17833
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 10048 17867 10100 17876
rect 10048 17833 10057 17867
rect 10057 17833 10091 17867
rect 10091 17833 10100 17867
rect 10048 17824 10100 17833
rect 11060 17824 11112 17876
rect 13360 17867 13412 17876
rect 13360 17833 13369 17867
rect 13369 17833 13403 17867
rect 13403 17833 13412 17867
rect 13360 17824 13412 17833
rect 15476 17824 15528 17876
rect 15752 17867 15804 17876
rect 15752 17833 15761 17867
rect 15761 17833 15795 17867
rect 15795 17833 15804 17867
rect 15752 17824 15804 17833
rect 2228 17756 2280 17808
rect 5356 17756 5408 17808
rect 6644 17756 6696 17808
rect 10876 17799 10928 17808
rect 10876 17765 10885 17799
rect 10885 17765 10919 17799
rect 10919 17765 10928 17799
rect 10876 17756 10928 17765
rect 12532 17756 12584 17808
rect 12992 17756 13044 17808
rect 8944 17688 8996 17740
rect 11244 17688 11296 17740
rect 12348 17688 12400 17740
rect 13820 17756 13872 17808
rect 5172 17620 5224 17672
rect 6184 17620 6236 17672
rect 11888 17663 11940 17672
rect 2688 17552 2740 17604
rect 7012 17552 7064 17604
rect 9496 17552 9548 17604
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 16120 17688 16172 17740
rect 17224 17688 17276 17740
rect 17592 17688 17644 17740
rect 13912 17620 13964 17672
rect 1400 17484 1452 17536
rect 1860 17527 1912 17536
rect 1860 17493 1869 17527
rect 1869 17493 1903 17527
rect 1903 17493 1912 17527
rect 1860 17484 1912 17493
rect 4528 17484 4580 17536
rect 8576 17484 8628 17536
rect 11336 17527 11388 17536
rect 11336 17493 11345 17527
rect 11345 17493 11379 17527
rect 11379 17493 11388 17527
rect 11336 17484 11388 17493
rect 11796 17527 11848 17536
rect 11796 17493 11805 17527
rect 11805 17493 11839 17527
rect 11839 17493 11848 17527
rect 11796 17484 11848 17493
rect 12164 17484 12216 17536
rect 12992 17484 13044 17536
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 5356 17280 5408 17332
rect 8024 17280 8076 17332
rect 10140 17323 10192 17332
rect 10140 17289 10149 17323
rect 10149 17289 10183 17323
rect 10183 17289 10192 17323
rect 10140 17280 10192 17289
rect 12348 17280 12400 17332
rect 13912 17280 13964 17332
rect 16212 17280 16264 17332
rect 17224 17323 17276 17332
rect 6644 17255 6696 17264
rect 6644 17221 6653 17255
rect 6653 17221 6687 17255
rect 6687 17221 6696 17255
rect 6644 17212 6696 17221
rect 8392 17212 8444 17264
rect 2504 17144 2556 17196
rect 2688 17187 2740 17196
rect 2688 17153 2697 17187
rect 2697 17153 2731 17187
rect 2731 17153 2740 17187
rect 2688 17144 2740 17153
rect 4620 17144 4672 17196
rect 4528 17119 4580 17128
rect 4528 17085 4537 17119
rect 4537 17085 4571 17119
rect 4571 17085 4580 17119
rect 4528 17076 4580 17085
rect 6000 17144 6052 17196
rect 9220 17212 9272 17264
rect 11796 17212 11848 17264
rect 2136 17008 2188 17060
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 2504 17051 2556 17060
rect 2504 17017 2513 17051
rect 2513 17017 2547 17051
rect 2547 17017 2556 17051
rect 2504 17008 2556 17017
rect 3516 17008 3568 17060
rect 6460 17076 6512 17128
rect 9312 17144 9364 17196
rect 10048 17144 10100 17196
rect 10692 17144 10744 17196
rect 16120 17144 16172 17196
rect 13452 17119 13504 17128
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 14096 17076 14148 17128
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 24768 17255 24820 17264
rect 24768 17221 24777 17255
rect 24777 17221 24811 17255
rect 24811 17221 24820 17255
rect 24768 17212 24820 17221
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 17224 17076 17276 17128
rect 5540 17008 5592 17060
rect 5172 16983 5224 16992
rect 5172 16949 5181 16983
rect 5181 16949 5215 16983
rect 5215 16949 5224 16983
rect 5172 16940 5224 16949
rect 6184 16983 6236 16992
rect 6184 16949 6193 16983
rect 6193 16949 6227 16983
rect 6227 16949 6236 16983
rect 6184 16940 6236 16949
rect 7012 17051 7064 17060
rect 7012 17017 7021 17051
rect 7021 17017 7055 17051
rect 7055 17017 7064 17051
rect 7012 17008 7064 17017
rect 8576 17008 8628 17060
rect 7564 16940 7616 16992
rect 10140 16940 10192 16992
rect 10784 17008 10836 17060
rect 12072 17008 12124 17060
rect 14004 17008 14056 17060
rect 11152 16940 11204 16992
rect 12440 16983 12492 16992
rect 12440 16949 12449 16983
rect 12449 16949 12483 16983
rect 12483 16949 12492 16983
rect 12440 16940 12492 16949
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 17592 16983 17644 16992
rect 17592 16949 17601 16983
rect 17601 16949 17635 16983
rect 17635 16949 17644 16983
rect 17592 16940 17644 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 4344 16779 4396 16788
rect 4344 16745 4353 16779
rect 4353 16745 4387 16779
rect 4387 16745 4396 16779
rect 4344 16736 4396 16745
rect 5172 16779 5224 16788
rect 5172 16745 5181 16779
rect 5181 16745 5215 16779
rect 5215 16745 5224 16779
rect 5172 16736 5224 16745
rect 6184 16779 6236 16788
rect 6184 16745 6193 16779
rect 6193 16745 6227 16779
rect 6227 16745 6236 16779
rect 6184 16736 6236 16745
rect 7012 16736 7064 16788
rect 9496 16779 9548 16788
rect 9496 16745 9505 16779
rect 9505 16745 9539 16779
rect 9539 16745 9548 16779
rect 9496 16736 9548 16745
rect 10692 16736 10744 16788
rect 12440 16736 12492 16788
rect 13452 16736 13504 16788
rect 14004 16779 14056 16788
rect 14004 16745 14013 16779
rect 14013 16745 14047 16779
rect 14047 16745 14056 16779
rect 14004 16736 14056 16745
rect 2412 16668 2464 16720
rect 3056 16668 3108 16720
rect 5356 16668 5408 16720
rect 4252 16600 4304 16652
rect 4528 16600 4580 16652
rect 2320 16532 2372 16584
rect 5540 16600 5592 16652
rect 6000 16600 6052 16652
rect 11980 16668 12032 16720
rect 12164 16711 12216 16720
rect 12164 16677 12173 16711
rect 12173 16677 12207 16711
rect 12207 16677 12216 16711
rect 12164 16668 12216 16677
rect 12716 16668 12768 16720
rect 16028 16736 16080 16788
rect 7196 16600 7248 16652
rect 9772 16600 9824 16652
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 6184 16532 6236 16584
rect 10140 16532 10192 16584
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 11152 16532 11204 16584
rect 11888 16600 11940 16652
rect 12808 16600 12860 16652
rect 15752 16668 15804 16720
rect 11704 16532 11756 16584
rect 13084 16600 13136 16652
rect 14832 16600 14884 16652
rect 24676 16643 24728 16652
rect 24676 16609 24694 16643
rect 24694 16609 24728 16643
rect 24676 16600 24728 16609
rect 25044 16600 25096 16652
rect 13268 16532 13320 16584
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 2504 16464 2556 16516
rect 6368 16464 6420 16516
rect 8392 16464 8444 16516
rect 11336 16464 11388 16516
rect 11888 16464 11940 16516
rect 8668 16396 8720 16448
rect 10048 16396 10100 16448
rect 11796 16396 11848 16448
rect 18420 16396 18472 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2412 16192 2464 16244
rect 4620 16235 4672 16244
rect 4620 16201 4629 16235
rect 4629 16201 4663 16235
rect 4663 16201 4672 16235
rect 4620 16192 4672 16201
rect 4712 16192 4764 16244
rect 8852 16235 8904 16244
rect 7932 16124 7984 16176
rect 8392 16124 8444 16176
rect 8852 16201 8861 16235
rect 8861 16201 8895 16235
rect 8895 16201 8904 16235
rect 8852 16192 8904 16201
rect 10048 16192 10100 16244
rect 10876 16192 10928 16244
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 13084 16235 13136 16244
rect 13084 16201 13093 16235
rect 13093 16201 13127 16235
rect 13127 16201 13136 16235
rect 13084 16192 13136 16201
rect 13268 16192 13320 16244
rect 15752 16235 15804 16244
rect 15752 16201 15761 16235
rect 15761 16201 15795 16235
rect 15795 16201 15804 16235
rect 15752 16192 15804 16201
rect 16028 16192 16080 16244
rect 24676 16235 24728 16244
rect 24676 16201 24685 16235
rect 24685 16201 24719 16235
rect 24719 16201 24728 16235
rect 24676 16192 24728 16201
rect 10232 16124 10284 16176
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 3056 16031 3108 16040
rect 3056 15997 3065 16031
rect 3065 15997 3099 16031
rect 3099 15997 3108 16031
rect 3056 15988 3108 15997
rect 3516 15988 3568 16040
rect 7104 16056 7156 16108
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 9496 16056 9548 16108
rect 11888 16124 11940 16176
rect 12808 16099 12860 16108
rect 5356 15988 5408 16040
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 15660 16056 15712 16108
rect 6552 15920 6604 15972
rect 6920 15963 6972 15972
rect 6920 15929 6929 15963
rect 6929 15929 6963 15963
rect 6963 15929 6972 15963
rect 6920 15920 6972 15929
rect 7012 15963 7064 15972
rect 7012 15929 7021 15963
rect 7021 15929 7055 15963
rect 7055 15929 7064 15963
rect 7012 15920 7064 15929
rect 8576 15920 8628 15972
rect 8852 15920 8904 15972
rect 9404 15920 9456 15972
rect 10692 15920 10744 15972
rect 11336 15920 11388 15972
rect 12440 15963 12492 15972
rect 12440 15929 12449 15963
rect 12449 15929 12483 15963
rect 12483 15929 12492 15963
rect 12440 15920 12492 15929
rect 14832 15963 14884 15972
rect 14832 15929 14841 15963
rect 14841 15929 14875 15963
rect 14875 15929 14884 15963
rect 14832 15920 14884 15929
rect 2320 15852 2372 15904
rect 4252 15895 4304 15904
rect 4252 15861 4261 15895
rect 4261 15861 4295 15895
rect 4295 15861 4304 15895
rect 4252 15852 4304 15861
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 5172 15852 5224 15904
rect 6000 15852 6052 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 7932 15895 7984 15904
rect 7932 15861 7941 15895
rect 7941 15861 7975 15895
rect 7975 15861 7984 15895
rect 7932 15852 7984 15861
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 9680 15852 9732 15904
rect 11704 15852 11756 15904
rect 15476 15920 15528 15972
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2136 15648 2188 15700
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 3056 15648 3108 15700
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 7196 15691 7248 15700
rect 2228 15580 2280 15632
rect 6092 15580 6144 15632
rect 6276 15623 6328 15632
rect 6276 15589 6285 15623
rect 6285 15589 6319 15623
rect 6319 15589 6328 15623
rect 6276 15580 6328 15589
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 10140 15648 10192 15700
rect 11888 15691 11940 15700
rect 11888 15657 11897 15691
rect 11897 15657 11931 15691
rect 11931 15657 11940 15691
rect 11888 15648 11940 15657
rect 13084 15648 13136 15700
rect 14832 15691 14884 15700
rect 14832 15657 14841 15691
rect 14841 15657 14875 15691
rect 14875 15657 14884 15691
rect 14832 15648 14884 15657
rect 1308 15512 1360 15564
rect 2504 15555 2556 15564
rect 2504 15521 2513 15555
rect 2513 15521 2547 15555
rect 2547 15521 2556 15555
rect 2504 15512 2556 15521
rect 4528 15512 4580 15564
rect 9312 15580 9364 15632
rect 11152 15580 11204 15632
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 12808 15555 12860 15564
rect 12808 15521 12817 15555
rect 12817 15521 12851 15555
rect 12851 15521 12860 15555
rect 12808 15512 12860 15521
rect 15660 15512 15712 15564
rect 16304 15555 16356 15564
rect 16304 15521 16348 15555
rect 16348 15521 16356 15555
rect 16304 15512 16356 15521
rect 4344 15444 4396 15496
rect 7012 15444 7064 15496
rect 11244 15444 11296 15496
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 6552 15376 6604 15428
rect 9404 15419 9456 15428
rect 9404 15385 9413 15419
rect 9413 15385 9447 15419
rect 9447 15385 9456 15419
rect 9404 15376 9456 15385
rect 11060 15376 11112 15428
rect 11428 15376 11480 15428
rect 12440 15376 12492 15428
rect 4712 15308 4764 15360
rect 5540 15308 5592 15360
rect 6000 15351 6052 15360
rect 6000 15317 6009 15351
rect 6009 15317 6043 15351
rect 6043 15317 6052 15351
rect 6000 15308 6052 15317
rect 6276 15308 6328 15360
rect 6920 15308 6972 15360
rect 7104 15308 7156 15360
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 8852 15351 8904 15360
rect 8852 15317 8861 15351
rect 8861 15317 8895 15351
rect 8895 15317 8904 15351
rect 8852 15308 8904 15317
rect 9772 15308 9824 15360
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 16672 15308 16724 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1308 15104 1360 15156
rect 2504 15104 2556 15156
rect 4344 15147 4396 15156
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 4712 15147 4764 15156
rect 4712 15113 4721 15147
rect 4721 15113 4755 15147
rect 4755 15113 4764 15147
rect 4712 15104 4764 15113
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 9312 15104 9364 15156
rect 9680 15104 9732 15156
rect 9956 15104 10008 15156
rect 11152 15147 11204 15156
rect 11152 15113 11161 15147
rect 11161 15113 11195 15147
rect 11195 15113 11204 15147
rect 11152 15104 11204 15113
rect 11244 15104 11296 15156
rect 14648 15104 14700 15156
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 10692 15036 10744 15088
rect 12808 15036 12860 15088
rect 5724 14968 5776 15020
rect 9680 14968 9732 15020
rect 2964 14900 3016 14952
rect 7380 14900 7432 14952
rect 9956 14900 10008 14952
rect 3884 14832 3936 14884
rect 5356 14875 5408 14884
rect 5356 14841 5365 14875
rect 5365 14841 5399 14875
rect 5399 14841 5408 14875
rect 5356 14832 5408 14841
rect 6092 14832 6144 14884
rect 6184 14832 6236 14884
rect 7012 14832 7064 14884
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 6368 14764 6420 14816
rect 6644 14764 6696 14816
rect 7288 14832 7340 14884
rect 10048 14832 10100 14884
rect 12348 14900 12400 14952
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 4528 14603 4580 14612
rect 4528 14569 4537 14603
rect 4537 14569 4571 14603
rect 4571 14569 4580 14603
rect 4528 14560 4580 14569
rect 5356 14560 5408 14612
rect 2872 14492 2924 14544
rect 3792 14492 3844 14544
rect 3884 14492 3936 14544
rect 6368 14492 6420 14544
rect 8024 14560 8076 14612
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 12808 14603 12860 14612
rect 12808 14569 12817 14603
rect 12817 14569 12851 14603
rect 12851 14569 12860 14603
rect 12808 14560 12860 14569
rect 16856 14603 16908 14612
rect 16856 14569 16865 14603
rect 16865 14569 16899 14603
rect 16899 14569 16908 14603
rect 16856 14560 16908 14569
rect 10048 14492 10100 14544
rect 10232 14492 10284 14544
rect 11980 14535 12032 14544
rect 11980 14501 11989 14535
rect 11989 14501 12023 14535
rect 12023 14501 12032 14535
rect 11980 14492 12032 14501
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 5264 14424 5316 14476
rect 5724 14467 5776 14476
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 7288 14424 7340 14476
rect 7748 14424 7800 14476
rect 16672 14467 16724 14476
rect 16672 14433 16681 14467
rect 16681 14433 16715 14467
rect 16715 14433 16724 14467
rect 16672 14424 16724 14433
rect 2228 14356 2280 14408
rect 2688 14356 2740 14408
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 6552 14356 6604 14408
rect 10048 14399 10100 14408
rect 10048 14365 10057 14399
rect 10057 14365 10091 14399
rect 10091 14365 10100 14399
rect 10048 14356 10100 14365
rect 11336 14356 11388 14408
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 10692 14220 10744 14272
rect 11336 14263 11388 14272
rect 11336 14229 11345 14263
rect 11345 14229 11379 14263
rect 11379 14229 11388 14263
rect 11336 14220 11388 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2872 14016 2924 14068
rect 3516 13948 3568 14000
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 5540 14016 5592 14068
rect 6184 14016 6236 14068
rect 6368 14016 6420 14068
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 7748 14016 7800 14068
rect 8024 14016 8076 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 6092 13948 6144 14000
rect 10140 14016 10192 14068
rect 10692 14016 10744 14068
rect 11980 14016 12032 14068
rect 16672 14059 16724 14068
rect 16672 14025 16681 14059
rect 16681 14025 16715 14059
rect 16715 14025 16724 14059
rect 16672 14016 16724 14025
rect 4528 13880 4580 13932
rect 5172 13855 5224 13864
rect 5172 13821 5181 13855
rect 5181 13821 5215 13855
rect 5215 13821 5224 13855
rect 5172 13812 5224 13821
rect 5264 13812 5316 13864
rect 5540 13812 5592 13864
rect 1860 13719 1912 13728
rect 1860 13685 1869 13719
rect 1869 13685 1903 13719
rect 1903 13685 1912 13719
rect 1860 13676 1912 13685
rect 2412 13719 2464 13728
rect 2412 13685 2421 13719
rect 2421 13685 2455 13719
rect 2455 13685 2464 13719
rect 2412 13676 2464 13685
rect 2964 13719 3016 13728
rect 2964 13685 2973 13719
rect 2973 13685 3007 13719
rect 3007 13685 3016 13719
rect 2964 13676 3016 13685
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 4712 13676 4764 13685
rect 4988 13676 5040 13728
rect 7380 13880 7432 13932
rect 11612 13948 11664 14000
rect 12164 13948 12216 14000
rect 8760 13880 8812 13932
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 10232 13880 10284 13932
rect 11336 13880 11388 13932
rect 6920 13787 6972 13796
rect 6920 13753 6929 13787
rect 6929 13753 6963 13787
rect 6963 13753 6972 13787
rect 6920 13744 6972 13753
rect 7012 13787 7064 13796
rect 7012 13753 7021 13787
rect 7021 13753 7055 13787
rect 7055 13753 7064 13787
rect 7012 13744 7064 13753
rect 8024 13744 8076 13796
rect 7196 13676 7248 13728
rect 9220 13812 9272 13864
rect 9956 13812 10008 13864
rect 8944 13787 8996 13796
rect 8944 13753 8953 13787
rect 8953 13753 8987 13787
rect 8987 13753 8996 13787
rect 8944 13744 8996 13753
rect 11336 13744 11388 13796
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2228 13515 2280 13524
rect 2228 13481 2237 13515
rect 2237 13481 2271 13515
rect 2271 13481 2280 13515
rect 2228 13472 2280 13481
rect 3516 13515 3568 13524
rect 1676 13336 1728 13388
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 6000 13472 6052 13524
rect 6920 13472 6972 13524
rect 7472 13472 7524 13524
rect 9220 13472 9272 13524
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 2596 13447 2648 13456
rect 2596 13413 2605 13447
rect 2605 13413 2639 13447
rect 2639 13413 2648 13447
rect 2596 13404 2648 13413
rect 3148 13447 3200 13456
rect 3148 13413 3157 13447
rect 3157 13413 3191 13447
rect 3191 13413 3200 13447
rect 3148 13404 3200 13413
rect 11336 13447 11388 13456
rect 11336 13413 11345 13447
rect 11345 13413 11379 13447
rect 11379 13413 11388 13447
rect 11336 13404 11388 13413
rect 4896 13336 4948 13388
rect 6092 13336 6144 13388
rect 7012 13336 7064 13388
rect 7104 13336 7156 13388
rect 8300 13336 8352 13388
rect 8944 13336 8996 13388
rect 10692 13379 10744 13388
rect 10692 13345 10701 13379
rect 10701 13345 10735 13379
rect 10735 13345 10744 13379
rect 10692 13336 10744 13345
rect 12072 13336 12124 13388
rect 1860 13268 1912 13320
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 4252 13200 4304 13252
rect 7932 13200 7984 13252
rect 8392 13200 8444 13252
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 6276 13132 6328 13184
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 7748 13175 7800 13184
rect 7748 13141 7757 13175
rect 7757 13141 7791 13175
rect 7791 13141 7800 13175
rect 7748 13132 7800 13141
rect 10048 13175 10100 13184
rect 10048 13141 10057 13175
rect 10057 13141 10091 13175
rect 10091 13141 10100 13175
rect 10048 13132 10100 13141
rect 18604 13132 18656 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 1860 12928 1912 12980
rect 4896 12928 4948 12980
rect 6092 12971 6144 12980
rect 6092 12937 6101 12971
rect 6101 12937 6135 12971
rect 6135 12937 6144 12971
rect 6092 12928 6144 12937
rect 6276 12928 6328 12980
rect 10692 12971 10744 12980
rect 10692 12937 10701 12971
rect 10701 12937 10735 12971
rect 10735 12937 10744 12971
rect 10692 12928 10744 12937
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 12072 12928 12124 12980
rect 7196 12860 7248 12912
rect 7748 12903 7800 12912
rect 7748 12869 7757 12903
rect 7757 12869 7791 12903
rect 7791 12869 7800 12903
rect 7748 12860 7800 12869
rect 2596 12792 2648 12844
rect 7288 12792 7340 12844
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 7748 12724 7800 12776
rect 9588 12767 9640 12776
rect 9588 12733 9597 12767
rect 9597 12733 9631 12767
rect 9631 12733 9640 12767
rect 9588 12724 9640 12733
rect 9680 12724 9732 12776
rect 11612 12724 11664 12776
rect 7380 12656 7432 12708
rect 8208 12656 8260 12708
rect 8300 12656 8352 12708
rect 10968 12656 11020 12708
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 9588 12588 9640 12640
rect 10048 12588 10100 12640
rect 12440 12588 12492 12640
rect 13820 12724 13872 12776
rect 13544 12699 13596 12708
rect 13544 12665 13553 12699
rect 13553 12665 13587 12699
rect 13587 12665 13596 12699
rect 13544 12656 13596 12665
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2872 12427 2924 12436
rect 2872 12393 2881 12427
rect 2881 12393 2915 12427
rect 2915 12393 2924 12427
rect 2872 12384 2924 12393
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 9680 12384 9732 12436
rect 9956 12316 10008 12368
rect 1584 12248 1636 12300
rect 2228 12248 2280 12300
rect 5080 12248 5132 12300
rect 7748 12291 7800 12300
rect 7748 12257 7792 12291
rect 7792 12257 7800 12291
rect 10232 12291 10284 12300
rect 7748 12248 7800 12257
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 10876 12248 10928 12300
rect 10968 12248 11020 12300
rect 12164 12248 12216 12300
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 13820 12291 13872 12300
rect 13820 12257 13829 12291
rect 13829 12257 13863 12291
rect 13863 12257 13872 12291
rect 13820 12248 13872 12257
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 14004 12223 14056 12232
rect 14004 12189 14013 12223
rect 14013 12189 14047 12223
rect 14047 12189 14056 12223
rect 14004 12180 14056 12189
rect 7288 12112 7340 12164
rect 8484 12112 8536 12164
rect 112 12044 164 12096
rect 8116 12044 8168 12096
rect 8392 12044 8444 12096
rect 10140 12044 10192 12096
rect 10784 12044 10836 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14372 12044 14424 12053
rect 15844 12087 15896 12096
rect 15844 12053 15853 12087
rect 15853 12053 15887 12087
rect 15887 12053 15896 12087
rect 15844 12044 15896 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2228 11883 2280 11892
rect 2228 11849 2237 11883
rect 2237 11849 2271 11883
rect 2271 11849 2280 11883
rect 2228 11840 2280 11849
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 9956 11840 10008 11892
rect 11980 11840 12032 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 27620 11840 27672 11892
rect 8760 11772 8812 11824
rect 10692 11772 10744 11824
rect 8944 11704 8996 11756
rect 1124 11636 1176 11688
rect 15844 11747 15896 11756
rect 15844 11713 15853 11747
rect 15853 11713 15887 11747
rect 15887 11713 15896 11747
rect 15844 11704 15896 11713
rect 16212 11747 16264 11756
rect 16212 11713 16221 11747
rect 16221 11713 16255 11747
rect 16255 11713 16264 11747
rect 16212 11704 16264 11713
rect 8760 11568 8812 11620
rect 10232 11568 10284 11620
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 8484 11500 8536 11509
rect 9956 11500 10008 11552
rect 10784 11636 10836 11688
rect 10968 11636 11020 11688
rect 12072 11636 12124 11688
rect 12624 11679 12676 11688
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 14372 11679 14424 11688
rect 14372 11645 14381 11679
rect 14381 11645 14415 11679
rect 14415 11645 14424 11679
rect 14372 11636 14424 11645
rect 15660 11636 15712 11688
rect 24216 11636 24268 11688
rect 11336 11568 11388 11620
rect 13176 11611 13228 11620
rect 13176 11577 13185 11611
rect 13185 11577 13219 11611
rect 13219 11577 13228 11611
rect 13176 11568 13228 11577
rect 10968 11500 11020 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 12900 11500 12952 11552
rect 13268 11500 13320 11552
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 10692 11339 10744 11348
rect 10692 11305 10701 11339
rect 10701 11305 10735 11339
rect 10735 11305 10744 11339
rect 10692 11296 10744 11305
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 14372 11339 14424 11348
rect 14372 11305 14381 11339
rect 14381 11305 14415 11339
rect 14415 11305 14424 11339
rect 14372 11296 14424 11305
rect 15844 11296 15896 11348
rect 13912 11228 13964 11280
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 10140 11160 10192 11212
rect 11152 11160 11204 11212
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 13544 11160 13596 11212
rect 14280 11160 14332 11212
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 16948 11024 17000 11076
rect 11336 10956 11388 11008
rect 12164 10956 12216 11008
rect 16304 10999 16356 11008
rect 16304 10965 16313 10999
rect 16313 10965 16347 10999
rect 16347 10965 16356 10999
rect 16304 10956 16356 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 12624 10752 12676 10804
rect 11888 10684 11940 10736
rect 13912 10752 13964 10804
rect 15476 10795 15528 10804
rect 10416 10616 10468 10668
rect 10968 10616 11020 10668
rect 12716 10616 12768 10668
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 14004 10616 14056 10668
rect 14372 10548 14424 10600
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 15660 10752 15712 10804
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 24952 10752 25004 10804
rect 15844 10684 15896 10736
rect 16304 10616 16356 10668
rect 11888 10480 11940 10532
rect 12624 10523 12676 10532
rect 12624 10489 12633 10523
rect 12633 10489 12667 10523
rect 12667 10489 12676 10523
rect 12624 10480 12676 10489
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 15292 10412 15344 10464
rect 15660 10412 15712 10464
rect 25228 10455 25280 10464
rect 25228 10421 25237 10455
rect 25237 10421 25271 10455
rect 25271 10421 25280 10455
rect 25228 10412 25280 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 10968 10251 11020 10260
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 11888 10251 11940 10260
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 12532 10208 12584 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 27620 10208 27672 10260
rect 13176 10140 13228 10192
rect 14004 10140 14056 10192
rect 15292 10140 15344 10192
rect 16212 10183 16264 10192
rect 16212 10149 16221 10183
rect 16221 10149 16255 10183
rect 16255 10149 16264 10183
rect 16212 10140 16264 10149
rect 10140 10072 10192 10124
rect 17040 10115 17092 10124
rect 17040 10081 17084 10115
rect 17084 10081 17092 10115
rect 24584 10115 24636 10124
rect 17040 10072 17092 10081
rect 24584 10081 24593 10115
rect 24593 10081 24627 10115
rect 24627 10081 24636 10115
rect 24584 10072 24636 10081
rect 10232 10004 10284 10056
rect 12348 10004 12400 10056
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 12716 9936 12768 9988
rect 15660 10004 15712 10056
rect 18880 9936 18932 9988
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 10140 9664 10192 9716
rect 11888 9707 11940 9716
rect 11888 9673 11897 9707
rect 11897 9673 11931 9707
rect 11931 9673 11940 9707
rect 11888 9664 11940 9673
rect 12532 9664 12584 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 10692 9596 10744 9648
rect 12808 9664 12860 9716
rect 13176 9664 13228 9716
rect 15292 9664 15344 9716
rect 15568 9707 15620 9716
rect 15568 9673 15577 9707
rect 15577 9673 15611 9707
rect 15611 9673 15620 9707
rect 15568 9664 15620 9673
rect 17040 9707 17092 9716
rect 17040 9673 17049 9707
rect 17049 9673 17083 9707
rect 17083 9673 17092 9707
rect 17040 9664 17092 9673
rect 24676 9707 24728 9716
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 25228 9664 25280 9716
rect 12716 9596 12768 9648
rect 13360 9596 13412 9648
rect 23388 9596 23440 9648
rect 12808 9528 12860 9580
rect 15292 9460 15344 9512
rect 10876 9435 10928 9444
rect 10876 9401 10885 9435
rect 10885 9401 10919 9435
rect 10919 9401 10928 9435
rect 10876 9392 10928 9401
rect 9496 9324 9548 9376
rect 10140 9324 10192 9376
rect 11244 9392 11296 9444
rect 12624 9435 12676 9444
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 24584 9460 24636 9512
rect 23480 9367 23532 9376
rect 23480 9333 23489 9367
rect 23489 9333 23523 9367
rect 23523 9333 23532 9367
rect 23480 9324 23532 9333
rect 24124 9367 24176 9376
rect 24124 9333 24133 9367
rect 24133 9333 24167 9367
rect 24167 9333 24176 9367
rect 24124 9324 24176 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 9496 9120 9548 9172
rect 10876 9163 10928 9172
rect 10876 9129 10885 9163
rect 10885 9129 10919 9163
rect 10919 9129 10928 9163
rect 10876 9120 10928 9129
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 15660 9120 15712 9172
rect 8208 9052 8260 9104
rect 11336 9095 11388 9104
rect 11336 9061 11345 9095
rect 11345 9061 11379 9095
rect 11379 9061 11388 9095
rect 11336 9052 11388 9061
rect 24124 9052 24176 9104
rect 24584 9095 24636 9104
rect 24584 9061 24593 9095
rect 24593 9061 24627 9095
rect 24627 9061 24636 9095
rect 24584 9052 24636 9061
rect 7380 8984 7432 9036
rect 7564 8984 7616 9036
rect 10692 8984 10744 9036
rect 8760 8916 8812 8968
rect 11888 8916 11940 8968
rect 23388 8916 23440 8968
rect 8392 8848 8444 8900
rect 8208 8780 8260 8832
rect 11244 8780 11296 8832
rect 11612 8823 11664 8832
rect 11612 8789 11621 8823
rect 11621 8789 11655 8823
rect 11655 8789 11664 8823
rect 11612 8780 11664 8789
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 14464 8823 14516 8832
rect 14464 8789 14473 8823
rect 14473 8789 14507 8823
rect 14507 8789 14516 8823
rect 14464 8780 14516 8789
rect 24860 8823 24912 8832
rect 24860 8789 24869 8823
rect 24869 8789 24903 8823
rect 24903 8789 24912 8823
rect 24860 8780 24912 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 10692 8576 10744 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 14372 8619 14424 8628
rect 14372 8585 14381 8619
rect 14381 8585 14415 8619
rect 14415 8585 14424 8619
rect 14372 8576 14424 8585
rect 23388 8619 23440 8628
rect 23388 8585 23397 8619
rect 23397 8585 23431 8619
rect 23431 8585 23440 8619
rect 23388 8576 23440 8585
rect 24124 8576 24176 8628
rect 8024 8508 8076 8560
rect 24676 8551 24728 8560
rect 24676 8517 24685 8551
rect 24685 8517 24719 8551
rect 24719 8517 24728 8551
rect 24676 8508 24728 8517
rect 8760 8440 8812 8492
rect 10876 8440 10928 8492
rect 14464 8483 14516 8492
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 24860 8440 24912 8492
rect 2044 8372 2096 8424
rect 13360 8415 13412 8424
rect 1768 8304 1820 8356
rect 2412 8304 2464 8356
rect 8208 8347 8260 8356
rect 8208 8313 8217 8347
rect 8217 8313 8251 8347
rect 8251 8313 8260 8347
rect 8208 8304 8260 8313
rect 8576 8304 8628 8356
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13360 8372 13412 8381
rect 14372 8304 14424 8356
rect 15660 8304 15712 8356
rect 23480 8304 23532 8356
rect 2044 8279 2096 8288
rect 2044 8245 2053 8279
rect 2053 8245 2087 8279
rect 2087 8245 2096 8279
rect 2044 8236 2096 8245
rect 6552 8236 6604 8288
rect 7380 8236 7432 8288
rect 7564 8279 7616 8288
rect 7564 8245 7573 8279
rect 7573 8245 7607 8279
rect 7607 8245 7616 8279
rect 7564 8236 7616 8245
rect 8024 8279 8076 8288
rect 8024 8245 8033 8279
rect 8033 8245 8067 8279
rect 8067 8245 8076 8279
rect 8024 8236 8076 8245
rect 8852 8279 8904 8288
rect 8852 8245 8861 8279
rect 8861 8245 8895 8279
rect 8895 8245 8904 8279
rect 8852 8236 8904 8245
rect 11244 8236 11296 8288
rect 11428 8236 11480 8288
rect 11612 8236 11664 8288
rect 12900 8236 12952 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 6184 8032 6236 8084
rect 8760 8032 8812 8084
rect 11336 8075 11388 8084
rect 11336 8041 11345 8075
rect 11345 8041 11379 8075
rect 11379 8041 11388 8075
rect 11336 8032 11388 8041
rect 11980 8032 12032 8084
rect 13360 8032 13412 8084
rect 15660 8075 15712 8084
rect 15660 8041 15669 8075
rect 15669 8041 15703 8075
rect 15703 8041 15712 8075
rect 15660 8032 15712 8041
rect 7196 7896 7248 7948
rect 11520 7939 11572 7948
rect 11520 7905 11529 7939
rect 11529 7905 11563 7939
rect 11563 7905 11572 7939
rect 11520 7896 11572 7905
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 14464 7896 14516 7948
rect 23204 7939 23256 7948
rect 23204 7905 23222 7939
rect 23222 7905 23256 7939
rect 27620 8032 27672 8084
rect 24676 7964 24728 8016
rect 24860 8007 24912 8016
rect 24860 7973 24869 8007
rect 24869 7973 24903 8007
rect 24903 7973 24912 8007
rect 24860 7964 24912 7973
rect 23204 7896 23256 7905
rect 6644 7828 6696 7880
rect 8484 7828 8536 7880
rect 10968 7828 11020 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 15660 7828 15712 7880
rect 7564 7760 7616 7812
rect 24768 7760 24820 7812
rect 7012 7692 7064 7744
rect 8024 7692 8076 7744
rect 8576 7735 8628 7744
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 12164 7692 12216 7744
rect 14372 7735 14424 7744
rect 14372 7701 14381 7735
rect 14381 7701 14415 7735
rect 14415 7701 14424 7735
rect 14372 7692 14424 7701
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 24124 7692 24176 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1400 7488 1452 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 8576 7488 8628 7540
rect 10784 7488 10836 7540
rect 11520 7488 11572 7540
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 14280 7488 14332 7540
rect 14464 7531 14516 7540
rect 14464 7497 14473 7531
rect 14473 7497 14507 7531
rect 14507 7497 14516 7531
rect 14464 7488 14516 7497
rect 15660 7531 15712 7540
rect 15660 7497 15669 7531
rect 15669 7497 15703 7531
rect 15703 7497 15712 7531
rect 15660 7488 15712 7497
rect 23204 7531 23256 7540
rect 23204 7497 23213 7531
rect 23213 7497 23247 7531
rect 23247 7497 23256 7531
rect 23204 7488 23256 7497
rect 8024 7420 8076 7472
rect 9956 7420 10008 7472
rect 11428 7420 11480 7472
rect 15568 7420 15620 7472
rect 24860 7463 24912 7472
rect 24860 7429 24869 7463
rect 24869 7429 24903 7463
rect 24903 7429 24912 7463
rect 24860 7420 24912 7429
rect 10968 7352 11020 7404
rect 204 7284 256 7336
rect 4988 7284 5040 7336
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 7656 7284 7708 7336
rect 9404 7284 9456 7336
rect 12900 7284 12952 7336
rect 24124 7352 24176 7404
rect 14372 7284 14424 7336
rect 15936 7284 15988 7336
rect 6920 7216 6972 7268
rect 9772 7259 9824 7268
rect 9772 7225 9781 7259
rect 9781 7225 9815 7259
rect 9815 7225 9824 7259
rect 9772 7216 9824 7225
rect 10784 7259 10836 7268
rect 10784 7225 10793 7259
rect 10793 7225 10827 7259
rect 10827 7225 10836 7259
rect 10784 7216 10836 7225
rect 11612 7216 11664 7268
rect 11980 7216 12032 7268
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 8024 7148 8076 7200
rect 10140 7148 10192 7200
rect 11520 7148 11572 7200
rect 12072 7148 12124 7200
rect 14188 7259 14240 7268
rect 14188 7225 14197 7259
rect 14197 7225 14231 7259
rect 14231 7225 14240 7259
rect 14188 7216 14240 7225
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 24492 7148 24544 7200
rect 24676 7148 24728 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 15384 6987 15436 6996
rect 15384 6953 15393 6987
rect 15393 6953 15427 6987
rect 15427 6953 15436 6987
rect 15384 6944 15436 6953
rect 24124 6987 24176 6996
rect 24124 6953 24133 6987
rect 24133 6953 24167 6987
rect 24167 6953 24176 6987
rect 24124 6944 24176 6953
rect 7196 6919 7248 6928
rect 7196 6885 7205 6919
rect 7205 6885 7239 6919
rect 7239 6885 7248 6919
rect 7196 6876 7248 6885
rect 13544 6919 13596 6928
rect 13544 6885 13553 6919
rect 13553 6885 13587 6919
rect 13587 6885 13596 6919
rect 13544 6876 13596 6885
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 1952 6808 2004 6860
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 8024 6808 8076 6817
rect 8852 6808 8904 6860
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 10232 6672 10284 6724
rect 10784 6672 10836 6724
rect 14280 6808 14332 6860
rect 15660 6808 15712 6860
rect 15936 6808 15988 6860
rect 23940 6808 23992 6860
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 25504 6808 25556 6860
rect 11244 6740 11296 6792
rect 11888 6740 11940 6792
rect 14096 6783 14148 6792
rect 11428 6715 11480 6724
rect 11428 6681 11437 6715
rect 11437 6681 11471 6715
rect 11471 6681 11480 6715
rect 11428 6672 11480 6681
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 14004 6672 14056 6724
rect 22100 6672 22152 6724
rect 24032 6672 24084 6724
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 10968 6604 11020 6656
rect 11336 6647 11388 6656
rect 11336 6613 11360 6647
rect 11360 6613 11388 6647
rect 11336 6604 11388 6613
rect 11612 6647 11664 6656
rect 11612 6613 11621 6647
rect 11621 6613 11655 6647
rect 11655 6613 11664 6647
rect 11612 6604 11664 6613
rect 24860 6647 24912 6656
rect 24860 6613 24869 6647
rect 24869 6613 24903 6647
rect 24903 6613 24912 6647
rect 24860 6604 24912 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 4988 6400 5040 6452
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10232 6443 10284 6452
rect 10232 6409 10241 6443
rect 10241 6409 10275 6443
rect 10275 6409 10284 6443
rect 10232 6400 10284 6409
rect 11428 6400 11480 6452
rect 1860 6264 1912 6316
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1952 6239 2004 6248
rect 1768 6196 1820 6205
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 6920 6196 6972 6205
rect 8852 6332 8904 6384
rect 12716 6332 12768 6384
rect 13544 6332 13596 6384
rect 8760 6264 8812 6316
rect 7656 6171 7708 6180
rect 7656 6137 7665 6171
rect 7665 6137 7699 6171
rect 7699 6137 7708 6171
rect 7656 6128 7708 6137
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 6920 6060 6972 6112
rect 9680 6196 9732 6248
rect 12072 6264 12124 6316
rect 12256 6264 12308 6316
rect 10876 6196 10928 6248
rect 11612 6196 11664 6248
rect 8944 6128 8996 6180
rect 11520 6171 11572 6180
rect 11520 6137 11529 6171
rect 11529 6137 11563 6171
rect 11563 6137 11572 6171
rect 11520 6128 11572 6137
rect 14832 6400 14884 6452
rect 15568 6400 15620 6452
rect 15660 6400 15712 6452
rect 15936 6400 15988 6452
rect 23940 6443 23992 6452
rect 23940 6409 23949 6443
rect 23949 6409 23983 6443
rect 23983 6409 23992 6443
rect 23940 6400 23992 6409
rect 14004 6375 14056 6384
rect 14004 6341 14013 6375
rect 14013 6341 14047 6375
rect 14047 6341 14056 6375
rect 14004 6332 14056 6341
rect 25504 6375 25556 6384
rect 25504 6341 25513 6375
rect 25513 6341 25547 6375
rect 25547 6341 25556 6375
rect 25504 6332 25556 6341
rect 27620 6332 27672 6384
rect 14740 6264 14792 6316
rect 15384 6264 15436 6316
rect 23296 6264 23348 6316
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 14832 6128 14884 6180
rect 23848 6128 23900 6180
rect 24768 6171 24820 6180
rect 24768 6137 24777 6171
rect 24777 6137 24811 6171
rect 24811 6137 24820 6171
rect 24768 6128 24820 6137
rect 18236 6103 18288 6112
rect 12164 6060 12216 6069
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1676 5899 1728 5908
rect 1676 5865 1685 5899
rect 1685 5865 1719 5899
rect 1719 5865 1728 5899
rect 1676 5856 1728 5865
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 11244 5899 11296 5908
rect 11244 5865 11253 5899
rect 11253 5865 11287 5899
rect 11287 5865 11296 5899
rect 11244 5856 11296 5865
rect 11336 5856 11388 5908
rect 12256 5856 12308 5908
rect 14096 5856 14148 5908
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 15568 5856 15620 5908
rect 8116 5831 8168 5840
rect 8116 5797 8125 5831
rect 8125 5797 8159 5831
rect 8159 5797 8168 5831
rect 8116 5788 8168 5797
rect 8208 5831 8260 5840
rect 8208 5797 8217 5831
rect 8217 5797 8251 5831
rect 8251 5797 8260 5831
rect 8208 5788 8260 5797
rect 9404 5788 9456 5840
rect 9772 5788 9824 5840
rect 12164 5788 12216 5840
rect 18604 5788 18656 5840
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 11520 5720 11572 5772
rect 13728 5720 13780 5772
rect 14188 5720 14240 5772
rect 16856 5720 16908 5772
rect 23848 5763 23900 5772
rect 23848 5729 23857 5763
rect 23857 5729 23891 5763
rect 23891 5729 23900 5763
rect 23848 5720 23900 5729
rect 9956 5652 10008 5704
rect 9864 5584 9916 5636
rect 17868 5652 17920 5704
rect 18236 5652 18288 5704
rect 19156 5627 19208 5636
rect 19156 5593 19165 5627
rect 19165 5593 19199 5627
rect 19199 5593 19208 5627
rect 19156 5584 19208 5593
rect 8944 5516 8996 5568
rect 13636 5559 13688 5568
rect 13636 5525 13645 5559
rect 13645 5525 13679 5559
rect 13679 5525 13688 5559
rect 13636 5516 13688 5525
rect 18236 5516 18288 5568
rect 24032 5559 24084 5568
rect 24032 5525 24041 5559
rect 24041 5525 24075 5559
rect 24075 5525 24084 5559
rect 24032 5516 24084 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1308 5312 1360 5364
rect 1860 5312 1912 5364
rect 8116 5312 8168 5364
rect 9772 5312 9824 5364
rect 9956 5312 10008 5364
rect 11520 5312 11572 5364
rect 13636 5312 13688 5364
rect 14464 5312 14516 5364
rect 15568 5312 15620 5364
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 17868 5355 17920 5364
rect 17868 5321 17877 5355
rect 17877 5321 17911 5355
rect 17911 5321 17920 5355
rect 17868 5312 17920 5321
rect 23848 5312 23900 5364
rect 24032 5355 24084 5364
rect 24032 5321 24041 5355
rect 24041 5321 24075 5355
rect 24075 5321 24084 5355
rect 24032 5312 24084 5321
rect 8208 5244 8260 5296
rect 8944 5244 8996 5296
rect 12164 5287 12216 5296
rect 12164 5253 12173 5287
rect 12173 5253 12207 5287
rect 12207 5253 12216 5287
rect 12164 5244 12216 5253
rect 13728 5287 13780 5296
rect 13728 5253 13737 5287
rect 13737 5253 13771 5287
rect 13771 5253 13780 5287
rect 13728 5244 13780 5253
rect 7656 5176 7708 5228
rect 9036 5176 9088 5228
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 12440 5176 12492 5228
rect 14096 5176 14148 5228
rect 15384 5176 15436 5228
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 24768 5244 24820 5296
rect 112 5108 164 5160
rect 8944 5040 8996 5092
rect 10048 5040 10100 5092
rect 2136 4972 2188 5024
rect 3424 4972 3476 5024
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 10140 4972 10192 5024
rect 12624 5040 12676 5092
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 15936 5083 15988 5092
rect 14464 5040 14516 5049
rect 15936 5049 15945 5083
rect 15945 5049 15979 5083
rect 15979 5049 15988 5083
rect 15936 5040 15988 5049
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 15660 5015 15712 5024
rect 15660 4981 15669 5015
rect 15669 4981 15703 5015
rect 15703 4981 15712 5015
rect 18236 5040 18288 5092
rect 24216 5083 24268 5092
rect 24216 5049 24225 5083
rect 24225 5049 24259 5083
rect 24259 5049 24268 5083
rect 24216 5040 24268 5049
rect 18604 5015 18656 5024
rect 15660 4972 15712 4981
rect 18604 4981 18613 5015
rect 18613 4981 18647 5015
rect 18647 4981 18656 5015
rect 18604 4972 18656 4981
rect 24032 4972 24084 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 10048 4768 10100 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 18696 4768 18748 4820
rect 24216 4811 24268 4820
rect 24216 4777 24225 4811
rect 24225 4777 24259 4811
rect 24259 4777 24268 4811
rect 24216 4768 24268 4777
rect 9036 4743 9088 4752
rect 9036 4709 9045 4743
rect 9045 4709 9079 4743
rect 9079 4709 9088 4743
rect 9036 4700 9088 4709
rect 9588 4700 9640 4752
rect 10784 4700 10836 4752
rect 12624 4743 12676 4752
rect 12624 4709 12633 4743
rect 12633 4709 12667 4743
rect 12667 4709 12676 4743
rect 12624 4700 12676 4709
rect 15936 4700 15988 4752
rect 12716 4675 12768 4684
rect 12716 4641 12725 4675
rect 12725 4641 12759 4675
rect 12759 4641 12768 4675
rect 12716 4632 12768 4641
rect 15384 4632 15436 4684
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 22928 4632 22980 4684
rect 24676 4675 24728 4684
rect 24676 4641 24694 4675
rect 24694 4641 24728 4675
rect 24676 4632 24728 4641
rect 27620 4632 27672 4684
rect 9864 4564 9916 4616
rect 10416 4564 10468 4616
rect 15752 4428 15804 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1216 4224 1268 4276
rect 9680 4224 9732 4276
rect 10416 4267 10468 4276
rect 10416 4233 10425 4267
rect 10425 4233 10459 4267
rect 10459 4233 10468 4267
rect 10416 4224 10468 4233
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 13636 4267 13688 4276
rect 13636 4233 13645 4267
rect 13645 4233 13679 4267
rect 13679 4233 13688 4267
rect 13636 4224 13688 4233
rect 15384 4267 15436 4276
rect 15384 4233 15393 4267
rect 15393 4233 15427 4267
rect 15427 4233 15436 4267
rect 15384 4224 15436 4233
rect 18236 4267 18288 4276
rect 18236 4233 18245 4267
rect 18245 4233 18279 4267
rect 18279 4233 18288 4267
rect 18236 4224 18288 4233
rect 19156 4224 19208 4276
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 15660 4088 15712 4140
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 112 4020 164 4072
rect 9588 4020 9640 4072
rect 13636 4020 13688 4072
rect 19156 4020 19208 4072
rect 10140 3952 10192 4004
rect 19156 3884 19208 3936
rect 22836 3884 22888 3936
rect 24768 3884 24820 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 9956 3544 10008 3596
rect 10784 3544 10836 3596
rect 15752 3544 15804 3596
rect 16212 3587 16264 3596
rect 16212 3553 16221 3587
rect 16221 3553 16255 3587
rect 16255 3553 16264 3587
rect 16212 3544 16264 3553
rect 19156 3587 19208 3596
rect 19156 3553 19165 3587
rect 19165 3553 19199 3587
rect 19199 3553 19208 3587
rect 19156 3544 19208 3553
rect 8576 3476 8628 3528
rect 9680 3340 9732 3392
rect 18328 3340 18380 3392
rect 20168 3340 20220 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 9956 3136 10008 3188
rect 16212 3179 16264 3188
rect 16212 3145 16221 3179
rect 16221 3145 16255 3179
rect 16255 3145 16264 3179
rect 16212 3136 16264 3145
rect 19156 3179 19208 3188
rect 19156 3145 19165 3179
rect 19165 3145 19199 3179
rect 19199 3145 19208 3179
rect 19156 3136 19208 3145
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 12808 2592 12860 2644
rect 16304 2592 16356 2644
rect 24860 2592 24912 2644
rect 7840 2524 7892 2576
rect 10048 2456 10100 2508
rect 11428 2320 11480 2372
rect 13728 2252 13780 2304
rect 15660 2252 15712 2304
rect 22100 2252 22152 2304
rect 26516 2252 26568 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 846 27520 902 28000
rect 2594 27520 2650 28000
rect 4342 27554 4398 28000
rect 4264 27526 4398 27554
rect 860 23662 888 27520
rect 1030 26616 1086 26625
rect 1030 26551 1086 26560
rect 848 23656 900 23662
rect 848 23598 900 23604
rect 1044 23186 1072 26551
rect 2226 25120 2282 25129
rect 2226 25055 2282 25064
rect 2240 24274 2268 25055
rect 2228 24268 2280 24274
rect 2228 24210 2280 24216
rect 2240 23866 2268 24210
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2608 23186 2636 27520
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3330 23488 3386 23497
rect 3330 23423 3386 23432
rect 1032 23180 1084 23186
rect 1032 23122 1084 23128
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 1596 22778 1624 23122
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1216 22024 1268 22030
rect 1216 21966 1268 21972
rect 1122 12608 1178 12617
rect 1122 12543 1178 12552
rect 112 12096 164 12102
rect 112 12038 164 12044
rect 124 11665 152 12038
rect 1136 11694 1164 12543
rect 1124 11688 1176 11694
rect 110 11656 166 11665
rect 1124 11630 1176 11636
rect 110 11591 166 11600
rect 204 7336 256 7342
rect 204 7278 256 7284
rect 216 7177 244 7278
rect 202 7168 258 7177
rect 202 7103 258 7112
rect 110 5400 166 5409
rect 110 5335 166 5344
rect 124 5166 152 5335
rect 112 5160 164 5166
rect 112 5102 164 5108
rect 1228 4282 1256 21966
rect 1872 21554 1900 22918
rect 2332 22574 2360 22918
rect 2608 22778 2636 23122
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 3344 22574 3372 23423
rect 2320 22568 2372 22574
rect 2320 22510 2372 22516
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2240 22166 2268 22374
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 2240 21690 2268 22102
rect 2228 21684 2280 21690
rect 2228 21626 2280 21632
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 2332 21418 2360 22510
rect 2780 21956 2832 21962
rect 2780 21898 2832 21904
rect 2792 21622 2820 21898
rect 2780 21616 2832 21622
rect 2780 21558 2832 21564
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 3332 21412 3384 21418
rect 3332 21354 3384 21360
rect 2044 21072 2096 21078
rect 2044 21014 2096 21020
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1676 20800 1728 20806
rect 1676 20742 1728 20748
rect 1688 20398 1716 20742
rect 1676 20392 1728 20398
rect 1582 20360 1638 20369
rect 1676 20334 1728 20340
rect 1582 20295 1638 20304
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 1306 18864 1362 18873
rect 1306 18799 1362 18808
rect 1320 15570 1348 18799
rect 1412 17882 1440 19654
rect 1596 19514 1624 20295
rect 1676 20256 1728 20262
rect 1676 20198 1728 20204
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1688 19310 1716 20198
rect 1964 19718 1992 20878
rect 2056 20398 2084 21014
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2412 20324 2464 20330
rect 2412 20266 2464 20272
rect 2320 19848 2372 19854
rect 2320 19790 2372 19796
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 2332 19378 2360 19790
rect 2424 19514 2452 20266
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 18902 2268 19246
rect 2044 18896 2096 18902
rect 2044 18838 2096 18844
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 1676 18692 1728 18698
rect 1676 18634 1728 18640
rect 1688 18222 1716 18634
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1400 17876 1452 17882
rect 1400 17818 1452 17824
rect 1872 17542 1900 18702
rect 2056 18426 2084 18838
rect 2332 18766 2360 19314
rect 2516 19242 2544 19926
rect 2608 19854 2636 20878
rect 2976 20466 3004 20946
rect 3344 20602 3372 21354
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2608 18698 2636 19790
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3344 19242 3372 19654
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 3332 19236 3384 19242
rect 3332 19178 3384 19184
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 2976 18222 3004 18566
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 3068 18086 3096 19178
rect 3436 18766 3464 24006
rect 4264 23866 4292 27526
rect 4342 27520 4398 27526
rect 5552 27526 6040 27554
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4264 23662 4292 23802
rect 4252 23656 4304 23662
rect 4252 23598 4304 23604
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 4436 23588 4488 23594
rect 4436 23530 4488 23536
rect 4712 23588 4764 23594
rect 4712 23530 4764 23536
rect 3700 23520 3752 23526
rect 3700 23462 3752 23468
rect 3712 23089 3740 23462
rect 4448 23225 4476 23530
rect 4434 23216 4490 23225
rect 4434 23151 4490 23160
rect 3698 23080 3754 23089
rect 3698 23015 3754 23024
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4632 22642 4660 22918
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4724 22506 4752 23530
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 3516 22024 3568 22030
rect 4252 22024 4304 22030
rect 3516 21966 3568 21972
rect 3882 21992 3938 22001
rect 3528 21690 3556 21966
rect 4252 21966 4304 21972
rect 3882 21927 3938 21936
rect 3896 21690 3924 21927
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 3700 21480 3752 21486
rect 3700 21422 3752 21428
rect 3514 19272 3570 19281
rect 3514 19207 3570 19216
rect 3528 19174 3556 19207
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3712 18358 3740 21422
rect 4264 19990 4292 21966
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4252 19984 4304 19990
rect 4252 19926 4304 19932
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4172 18834 4200 19110
rect 4264 18902 4292 19178
rect 4252 18896 4304 18902
rect 4252 18838 4304 18844
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4172 18426 4200 18770
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 4080 18086 4108 18362
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 2228 17808 2280 17814
rect 2228 17750 2280 17756
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15162 1348 15506
rect 1308 15156 1360 15162
rect 1308 15098 1360 15104
rect 1412 7546 1440 17478
rect 1858 17232 1914 17241
rect 1858 17167 1914 17176
rect 1872 16046 1900 17167
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 2148 15706 2176 17002
rect 2240 16998 2268 17750
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2700 17202 2728 17546
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2516 17066 2544 17138
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2240 15638 2268 16934
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2332 15910 2360 16526
rect 2424 16250 2452 16662
rect 2516 16522 2544 17002
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 15706 2360 15846
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2228 15632 2280 15638
rect 2228 15574 2280 15580
rect 2516 15570 2544 16458
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2516 15162 2544 15506
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2700 14414 2728 17138
rect 3068 16726 3096 18022
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3528 16794 3556 17002
rect 4356 16794 4384 21830
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4908 20534 4936 20878
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4434 19816 4490 19825
rect 4434 19751 4490 19760
rect 4448 19718 4476 19751
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4448 19242 4476 19654
rect 4816 19242 4844 20334
rect 4908 20058 4936 20470
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 5184 19990 5212 22918
rect 5264 22500 5316 22506
rect 5264 22442 5316 22448
rect 5276 22234 5304 22442
rect 5368 22438 5396 23122
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5276 21554 5304 22170
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5264 21412 5316 21418
rect 5368 21400 5396 22374
rect 5460 22166 5488 23598
rect 5448 22160 5500 22166
rect 5448 22102 5500 22108
rect 5460 21690 5488 22102
rect 5552 21894 5580 27526
rect 6012 27520 6040 27526
rect 6090 27520 6146 28000
rect 7838 27554 7894 28000
rect 9586 27554 9642 28000
rect 11334 27554 11390 28000
rect 7668 27526 7894 27554
rect 6012 27492 6132 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5316 21372 5396 21400
rect 5264 21354 5316 21360
rect 5276 20602 5304 21354
rect 5460 21146 5488 21626
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5356 21072 5408 21078
rect 5356 21014 5408 21020
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5368 20330 5396 21014
rect 5552 20806 5580 21490
rect 6196 20806 6224 21966
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5000 19446 5028 19926
rect 5184 19514 5212 19926
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 4988 19440 5040 19446
rect 4988 19382 5040 19388
rect 4436 19236 4488 19242
rect 4436 19178 4488 19184
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5276 18290 5304 18702
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4540 17134 4568 17478
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 3528 16046 3556 16730
rect 4540 16658 4568 17070
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3068 15706 3096 15982
rect 4264 15910 4292 16594
rect 4632 16250 4660 17138
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12306 1624 13126
rect 1688 12986 1716 13330
rect 1872 13326 1900 13670
rect 2240 13530 2268 14350
rect 2884 14074 2912 14486
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 12986 1900 13262
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 11898 2268 12242
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1596 9654 1624 9687
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1582 8800 1638 8809
rect 1582 8735 1638 8744
rect 1596 8634 1624 8735
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2044 8424 2096 8430
rect 2042 8392 2044 8401
rect 2096 8392 2098 8401
rect 1768 8356 1820 8362
rect 2424 8362 2452 13670
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2608 12850 2636 13398
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2884 12782 2912 14010
rect 2976 13734 3004 14894
rect 3068 13870 3096 15642
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 14550 3832 14758
rect 3896 14550 3924 14826
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3884 14544 3936 14550
rect 3884 14486 3936 14492
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 3160 13462 3188 14350
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3528 13530 3556 13942
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 4264 13258 4292 15846
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4356 15162 4384 15438
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4540 14618 4568 15506
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4540 13938 4568 14554
rect 4632 14482 4660 16186
rect 4724 15366 4752 16186
rect 4816 15910 4844 18158
rect 5264 18148 5316 18154
rect 5368 18136 5396 20266
rect 5552 19786 5580 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6196 20505 6224 20742
rect 6182 20496 6238 20505
rect 6182 20431 6238 20440
rect 6472 19922 6500 23462
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6840 21486 6868 21830
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6840 21146 6868 21422
rect 7116 21350 7144 22034
rect 7576 22030 7604 22374
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7576 21622 7604 21966
rect 7668 21690 7696 27526
rect 7838 27520 7894 27526
rect 9416 27526 9642 27554
rect 9416 24274 9444 27526
rect 9586 27520 9642 27526
rect 11072 27526 11390 27554
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 10784 24268 10836 24274
rect 10784 24210 10836 24216
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 9220 24064 9272 24070
rect 9220 24006 9272 24012
rect 8404 23662 8432 24006
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8760 23656 8812 23662
rect 8760 23598 8812 23604
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8220 22778 8248 23122
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7852 21554 7880 21898
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 8220 21418 8248 22714
rect 8312 22166 8340 22918
rect 8300 22160 8352 22166
rect 8300 22102 8352 22108
rect 8312 21690 8340 22102
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6472 19514 6500 19858
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18154 6040 18566
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 5316 18108 5396 18136
rect 5264 18090 5316 18096
rect 5368 17814 5396 18108
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 16998 5212 17614
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16794 5212 16934
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5368 16726 5396 17274
rect 6012 17202 6040 18090
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5262 16552 5318 16561
rect 5262 16487 5318 16496
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5078 15736 5134 15745
rect 5078 15671 5134 15680
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4724 15162 4752 15302
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4620 14476 4672 14482
rect 4672 14436 4752 14464
rect 4620 14418 4672 14424
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4724 13734 4752 14436
rect 4894 14240 4950 14249
rect 4894 14175 4950 14184
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4908 13394 4936 14175
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4908 12986 4936 13330
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12442 2912 12718
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2042 8327 2098 8336
rect 2412 8356 2464 8362
rect 1768 8298 1820 8304
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1688 5914 1716 6802
rect 1780 6254 1808 8298
rect 2056 8294 2084 8327
rect 2412 8298 2464 8304
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 5000 7342 5028 13670
rect 5092 12306 5120 15671
rect 5184 13870 5212 15846
rect 5276 15706 5304 16487
rect 5368 16046 5396 16662
rect 5552 16658 5580 17002
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 6000 16652 6052 16658
rect 6104 16640 6132 18362
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6196 16998 6224 17614
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 16794 6224 16934
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6052 16612 6132 16640
rect 6000 16594 6052 16600
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5552 15366 5580 16594
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 15910 6040 16594
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 15910 6224 16526
rect 6380 16522 6408 18022
rect 6472 17134 6500 19450
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6840 19281 6868 19314
rect 6826 19272 6882 19281
rect 6826 19207 6882 19216
rect 6840 18902 6868 19207
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6564 17882 6592 18838
rect 7116 18766 7144 21286
rect 8220 21146 8248 21354
rect 8588 21146 8616 23462
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8680 21962 8708 22578
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8680 21622 8708 21898
rect 8668 21616 8720 21622
rect 8668 21558 8720 21564
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7484 20398 7512 20742
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7484 19922 7512 20334
rect 7576 20058 7604 20878
rect 7944 20534 7972 21082
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 7932 20528 7984 20534
rect 7932 20470 7984 20476
rect 7932 20324 7984 20330
rect 7932 20266 7984 20272
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7944 19904 7972 20266
rect 8024 19916 8076 19922
rect 7944 19876 8024 19904
rect 7484 19446 7512 19858
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 18358 7144 18702
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6656 17270 6684 17750
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6552 15972 6604 15978
rect 6552 15914 6604 15920
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6092 15632 6144 15638
rect 6196 15620 6224 15846
rect 6144 15592 6224 15620
rect 6092 15574 6144 15580
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5368 14618 5396 14826
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 13870 5304 14418
rect 5552 14074 5580 15302
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5736 14482 5764 14962
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5552 13190 5580 13806
rect 6012 13530 6040 15302
rect 6196 14890 6224 15592
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6288 15366 6316 15574
rect 6564 15434 6592 15914
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6656 15162 6684 17206
rect 7024 17066 7052 17546
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 7024 16794 7052 17002
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 6918 16144 6974 16153
rect 6918 16079 6974 16088
rect 7104 16108 7156 16114
rect 6932 15978 6960 16079
rect 7104 16050 7156 16056
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7024 15502 7052 15914
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7116 15366 7144 16050
rect 7208 15706 7236 16594
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6104 14006 6132 14826
rect 6656 14822 6684 15098
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6380 14550 6408 14758
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6380 14074 6408 14486
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6564 14074 6592 14350
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6104 13394 6132 13942
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6104 12986 6132 13330
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6196 8090 6224 14010
rect 6932 13802 6960 15302
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7024 14090 7052 14826
rect 7300 14482 7328 14826
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7392 14278 7420 14894
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7024 14062 7144 14090
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 6932 13530 6960 13738
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7024 13394 7052 13738
rect 7116 13394 7144 14062
rect 7392 13938 7420 14214
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12986 6316 13126
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 7208 12918 7236 13670
rect 7484 13530 7512 19382
rect 7944 19174 7972 19876
rect 8024 19858 8076 19864
rect 8496 19174 8524 20946
rect 8588 20466 8616 21082
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 7944 18834 7972 19110
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 7944 18426 7972 18770
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 17882 7696 18158
rect 8036 17882 8064 18770
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8404 17882 8432 18226
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8036 17338 8064 17818
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 15366 7604 16934
rect 8404 16522 8432 17206
rect 8588 17066 8616 17478
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8404 16182 8432 16458
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8482 16144 8538 16153
rect 7944 15910 7972 16118
rect 8482 16079 8538 16088
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7208 12442 7236 12854
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7300 12646 7328 12786
rect 7392 12714 7420 13126
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7300 12170 7328 12582
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7576 9674 7604 15302
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14482 7788 14758
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14074 7788 14418
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7838 13968 7894 13977
rect 7838 13903 7894 13912
rect 7852 13326 7880 13903
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12918 7788 13126
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 7760 12782 7788 12854
rect 7852 12850 7880 13262
rect 7944 13258 7972 15846
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8036 15162 8064 15506
rect 8496 15162 8524 16079
rect 8588 15978 8616 17002
rect 8772 16561 8800 23598
rect 8852 22500 8904 22506
rect 8852 22442 8904 22448
rect 8864 22234 8892 22442
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 9232 22166 9260 24006
rect 9416 23866 9444 24210
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 10060 23662 10088 24006
rect 10796 23866 10824 24210
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10968 23860 11020 23866
rect 10968 23802 11020 23808
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9600 22642 9628 23122
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9220 22160 9272 22166
rect 9220 22102 9272 22108
rect 9508 21350 9536 22170
rect 9600 22030 9628 22442
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9508 20602 9536 21286
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8864 19310 8892 19858
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8758 16552 8814 16561
rect 8758 16487 8814 16496
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8680 16096 8708 16390
rect 8864 16250 8892 19246
rect 9600 18290 9628 21966
rect 9692 18358 9720 23598
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9784 21146 9812 22102
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 10060 20058 10088 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10980 23322 11008 23802
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22234 10180 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10888 21554 10916 21830
rect 11072 21690 11100 27526
rect 11334 27520 11390 27526
rect 13082 27520 13138 28000
rect 14830 27520 14886 28000
rect 16578 27520 16634 28000
rect 18326 27520 18382 28000
rect 20074 27520 20130 28000
rect 21822 27520 21878 28000
rect 23570 27520 23626 28000
rect 25318 27520 25374 28000
rect 27066 27520 27122 28000
rect 13096 24410 13124 27520
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11348 22778 11376 23122
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 11348 21418 11376 22714
rect 11532 22166 11560 22918
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11532 21690 11560 22102
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 11348 21146 11376 21354
rect 11808 21146 11836 21966
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10244 20602 10272 20946
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10612 20534 10640 21014
rect 11992 20806 12020 23598
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 13542 23080 13598 23089
rect 13542 23015 13598 23024
rect 13556 22982 13584 23015
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12820 22234 12848 22510
rect 13556 22234 13584 22918
rect 13740 22642 13768 23190
rect 13912 22704 13964 22710
rect 13912 22646 13964 22652
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12268 21418 12296 21898
rect 13740 21690 13768 21966
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10612 20330 10640 20470
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 10600 20324 10652 20330
rect 10652 20284 10732 20312
rect 10600 20266 10652 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20284
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10704 19514 10732 19994
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8956 17649 8984 17682
rect 8942 17640 8998 17649
rect 8942 17575 8998 17584
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8760 16108 8812 16114
rect 8680 16068 8760 16096
rect 8760 16050 8812 16056
rect 8576 15972 8628 15978
rect 8576 15914 8628 15920
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8864 15366 8892 15914
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8036 14618 8064 15098
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8036 13802 8064 14010
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8206 13832 8262 13841
rect 8024 13796 8076 13802
rect 8206 13767 8262 13776
rect 8024 13738 8076 13744
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 8220 12714 8248 13767
rect 8772 13734 8800 13874
rect 8864 13841 8892 15302
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8850 13832 8906 13841
rect 8956 13802 8984 14214
rect 9232 14074 9260 17206
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9324 15638 9352 17138
rect 9508 16794 9536 17546
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9404 15972 9456 15978
rect 9404 15914 9456 15920
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 9324 15162 9352 15574
rect 9416 15434 9444 15914
rect 9508 15910 9536 16050
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9404 15428 9456 15434
rect 9404 15370 9456 15376
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9232 13870 9260 14010
rect 9324 13938 9352 15098
rect 9508 13977 9536 15846
rect 9692 15162 9720 15846
rect 9784 15366 9812 16594
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9494 13968 9550 13977
rect 9312 13932 9364 13938
rect 9692 13938 9720 14962
rect 9494 13903 9550 13912
rect 9680 13932 9732 13938
rect 9312 13874 9364 13880
rect 9680 13874 9732 13880
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 8850 13767 8906 13776
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8312 12714 8340 13330
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7760 11898 7788 12242
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7576 9646 7788 9674
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7392 8294 7420 8978
rect 7576 8294 7604 8978
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1872 5778 1900 6258
rect 1964 6254 1992 6802
rect 5000 6458 5028 7278
rect 6564 6866 6592 8230
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6656 7546 6684 7822
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5370 1900 5714
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1216 4276 1268 4282
rect 1216 4218 1268 4224
rect 112 4072 164 4078
rect 112 4014 164 4020
rect 124 3777 152 4014
rect 110 3768 166 3777
rect 110 3703 166 3712
rect 1030 82 1086 480
rect 1320 82 1348 5306
rect 1964 1329 1992 6190
rect 2134 5128 2190 5137
rect 2134 5063 2190 5072
rect 2148 5030 2176 5063
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 1950 1320 2006 1329
rect 1950 1255 2006 1264
rect 1030 54 1348 82
rect 3146 82 3202 480
rect 3436 82 3464 4966
rect 3146 54 3464 82
rect 5000 82 5028 6394
rect 6564 6118 6592 6802
rect 6932 6254 6960 7210
rect 7024 7206 7052 7686
rect 7208 7342 7236 7890
rect 7576 7818 7604 8230
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7576 7324 7604 7754
rect 7656 7336 7708 7342
rect 7576 7296 7656 7324
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 6118 6960 6190
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6564 1601 6592 6054
rect 6932 5914 6960 6054
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 2825 7052 7142
rect 7208 6934 7236 7278
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7576 6662 7604 7296
rect 7656 7278 7708 7284
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7010 2816 7066 2825
rect 7010 2751 7066 2760
rect 6550 1592 6606 1601
rect 6550 1527 6606 1536
rect 5262 82 5318 480
rect 5000 54 5318 82
rect 1030 0 1086 54
rect 3146 0 3202 54
rect 5262 0 5318 54
rect 7470 82 7526 480
rect 7576 82 7604 6598
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7668 5234 7696 6122
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7760 4154 7788 9646
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8036 8294 8064 8502
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7750 8064 8230
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8036 6866 8064 7142
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8036 6458 8064 6802
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8128 5846 8156 12038
rect 8220 9110 8248 12650
rect 8404 12102 8432 13194
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8220 8838 8248 9046
rect 8404 8906 8432 12038
rect 8496 11558 8524 12106
rect 8772 11830 8800 13670
rect 8956 13394 8984 13738
rect 9232 13530 9260 13806
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 9692 12782 9720 13874
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9600 12646 9628 12718
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8772 11626 8800 11766
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8956 11665 8984 11698
rect 8942 11656 8998 11665
rect 8760 11620 8812 11626
rect 8942 11591 8998 11600
rect 8760 11562 8812 11568
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8362 8248 8774
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8496 7886 8524 11494
rect 8772 8974 8800 11562
rect 9600 11200 9628 12582
rect 9692 12442 9720 12718
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 11212 9732 11218
rect 9600 11172 9680 11200
rect 9680 11154 9732 11160
rect 9692 10470 9720 11154
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 9178 9536 9318
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8498 8800 8910
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8588 7750 8616 8298
rect 8772 8090 8800 8434
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8588 7546 8616 7686
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8864 6866 8892 8230
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8772 6322 8800 6734
rect 8864 6390 8892 6802
rect 9416 6458 9444 7278
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8128 5370 8156 5782
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8220 5302 8248 5782
rect 8956 5574 8984 6122
rect 9416 5846 9444 6394
rect 9692 6254 9720 10406
rect 9876 8401 9904 18634
rect 10060 17882 10088 19450
rect 10980 19242 11008 20198
rect 11072 19378 11100 20198
rect 11348 20058 11376 20334
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11348 19514 11376 19994
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 11072 18970 11100 19314
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 11716 18834 11744 19314
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10060 17202 10088 17818
rect 10152 17338 10180 18566
rect 10244 18154 10272 18770
rect 11716 18426 11744 18770
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 17196 10100 17202
rect 9968 17156 10048 17184
rect 9968 15162 9996 17156
rect 10048 17138 10100 17144
rect 10152 16998 10180 17274
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16794 10732 17138
rect 10796 17066 10824 18090
rect 10888 17814 10916 18226
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17882 11100 18022
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 11164 16590 11192 16934
rect 11256 16658 11284 17682
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16250 10088 16390
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10152 15706 10180 16526
rect 10244 16182 10272 16526
rect 11348 16522 11376 17478
rect 11808 17270 11836 17478
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9956 15156 10008 15162
rect 10008 15116 10088 15144
rect 9956 15098 10008 15104
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9968 14618 9996 14894
rect 10060 14890 10088 15116
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10060 14550 10088 14826
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9968 12374 9996 13806
rect 10060 13190 10088 14350
rect 10152 14074 10180 15642
rect 10704 15366 10732 15914
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 15094 10732 15302
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12850 10088 13126
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9968 11898 9996 12310
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9862 8392 9918 8401
rect 9862 8327 9918 8336
rect 9968 7478 9996 11494
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9784 5846 9812 7210
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5302 8984 5510
rect 9784 5370 9812 5782
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8956 5098 8984 5238
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 9048 4758 9076 5170
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4758 9628 4966
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9600 4264 9628 4694
rect 9876 4622 9904 5578
rect 9968 5370 9996 5646
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10060 5250 10088 12582
rect 10152 12102 10180 14010
rect 10244 13938 10272 14486
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10704 14074 10732 14214
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13394 10732 14010
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10704 12986 10732 13330
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10888 12306 10916 16186
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 13814 11100 15370
rect 11164 15162 11192 15574
rect 11348 15502 11376 15914
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11256 15162 11284 15438
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11348 14414 11376 15438
rect 11440 15434 11468 16594
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 15910 11744 16526
rect 11808 16454 11836 17206
rect 11900 16658 11928 17614
rect 11992 16726 12020 20742
rect 12268 19854 12296 21354
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12268 18970 12296 19790
rect 12360 19310 12388 21286
rect 12544 21010 12572 21286
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12912 20806 12940 21422
rect 13924 21146 13952 22646
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 22234 14136 22374
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 13004 20058 13032 20878
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 19378 12572 19790
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12360 19145 12388 19246
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12346 19136 12402 19145
rect 12346 19071 12402 19080
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12360 17746 12388 19071
rect 12544 18902 12572 19178
rect 13004 19174 13032 19994
rect 13372 19718 13400 20334
rect 13464 20262 13492 21014
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13176 19236 13228 19242
rect 13176 19178 13228 19184
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13188 18970 13216 19178
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12544 18630 12572 18838
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 17814 12572 18566
rect 12728 18222 12756 18770
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12728 18086 12756 18158
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16250 11836 16390
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11900 16182 11928 16458
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11900 15706 11928 16118
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 13938 11376 14214
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 10980 13786 11100 13814
rect 11336 13796 11388 13802
rect 10980 12714 11008 13786
rect 11336 13738 11388 13744
rect 11348 13462 11376 13738
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11624 12986 11652 13942
rect 11900 13530 11928 14350
rect 11992 14074 12020 14486
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 12084 13394 12112 17002
rect 12176 16726 12204 17478
rect 12360 17338 12388 17682
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12360 14958 12388 17274
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16794 12480 16934
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12728 16726 12756 18022
rect 13004 17814 13032 18158
rect 13372 17882 13400 19654
rect 13464 19446 13492 20198
rect 14200 20058 14228 20742
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13464 18154 13492 19382
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13740 18902 13768 19246
rect 13924 19174 13952 19382
rect 14016 19378 14044 19654
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 13912 19168 13964 19174
rect 13964 19128 14044 19156
rect 13912 19110 13964 19116
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13832 17814 13860 18022
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13004 17542 13032 17750
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13924 17338 13952 17614
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13464 16794 13492 17070
rect 14016 17066 14044 19128
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18290 14136 18566
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14292 17649 14320 24006
rect 14844 23866 14872 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 16500 23798 16528 24210
rect 16592 23866 16620 27520
rect 18340 24274 18368 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 17222 23760 17278 23769
rect 17222 23695 17278 23704
rect 17236 23662 17264 23695
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 14648 23588 14700 23594
rect 14648 23530 14700 23536
rect 16304 23588 16356 23594
rect 16304 23530 16356 23536
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 14554 23216 14610 23225
rect 14554 23151 14610 23160
rect 14568 23118 14596 23151
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14568 22642 14596 23054
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14476 20602 14504 21966
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14278 17640 14334 17649
rect 14278 17575 14334 17584
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14108 17134 14136 17478
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14016 16794 14044 17002
rect 13452 16788 13504 16794
rect 14004 16788 14056 16794
rect 13452 16730 13504 16736
rect 13924 16748 14004 16776
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12820 16114 12848 16594
rect 13096 16250 13124 16594
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13280 16250 13308 16526
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12452 15434 12480 15914
rect 13096 15706 13124 16186
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12820 15094 12848 15506
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 14006 12204 14350
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12360 13814 12388 14894
rect 12820 14618 12848 15030
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12360 13786 12480 13814
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12986 12112 13330
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11624 12782 11652 12922
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10980 12306 11008 12650
rect 12452 12646 12480 13786
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 13280 12306 13308 16186
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10244 11626 10272 12242
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11354 10732 11766
rect 10796 11694 10824 12038
rect 11992 11898 12020 12038
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12084 11694 12112 12174
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10810 10180 11154
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10152 10130 10180 10746
rect 10428 10674 10456 11086
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10152 9722 10180 10066
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10140 9376 10192 9382
rect 10244 9364 10272 9998
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10192 9336 10272 9364
rect 10140 9318 10192 9324
rect 10152 7206 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9042 10732 9590
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10704 8634 10732 8978
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10796 7546 10824 11630
rect 10980 11558 11008 11630
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 11218 11192 11494
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10980 10266 11008 10610
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11256 9450 11284 11086
rect 11348 11014 11376 11562
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 10888 9178 10916 9386
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10888 8498 10916 9114
rect 11348 9110 11376 10950
rect 11532 10810 11560 11154
rect 12176 11014 12204 12242
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12636 11354 12664 11630
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12624 11348 12676 11354
rect 12544 11308 12624 11336
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11900 10538 11928 10678
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 10266 11928 10474
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11900 9722 11928 10202
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11256 8294 11284 8774
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7970 11284 8230
rect 11348 8090 11376 9046
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11624 8294 11652 8774
rect 11900 8634 11928 8910
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11256 7942 11376 7970
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10784 7268 10836 7274
rect 10888 7256 10916 7686
rect 10980 7410 11008 7822
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10836 7228 10916 7256
rect 10784 7210 10836 7216
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 6730 10824 7210
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10244 6458 10272 6666
rect 10980 6662 11008 7346
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10888 5914 10916 6190
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10980 5681 11008 6598
rect 11256 5914 11284 6734
rect 11348 6662 11376 7942
rect 11440 7478 11468 8230
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11532 7546 11560 7890
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11440 6730 11468 7414
rect 11532 7206 11560 7482
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 5914 11376 6598
rect 11440 6458 11468 6666
rect 11624 6662 11652 7210
rect 11900 6798 11928 8570
rect 11992 8090 12020 8774
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7274 12020 7890
rect 12176 7750 12204 10950
rect 12544 10266 12572 11308
rect 12624 11290 12676 11296
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12636 10538 12664 10746
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12728 10266 12756 10610
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12360 9178 12388 9998
rect 12544 9722 12572 10202
rect 12728 9994 12756 10202
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12544 9432 12572 9658
rect 12728 9654 12756 9930
rect 12820 9722 12848 10610
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12624 9444 12676 9450
rect 12544 9404 12624 9432
rect 12624 9386 12676 9392
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12820 8838 12848 9522
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11624 6254 11652 6598
rect 12084 6322 12112 7142
rect 12268 6322 12296 7822
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11532 5778 11560 6122
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 5846 12204 6054
rect 12268 5914 12296 6258
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 9968 5222 10088 5250
rect 10784 5228 10836 5234
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9680 4276 9732 4282
rect 9600 4236 9680 4264
rect 7760 4126 7880 4154
rect 7852 2582 7880 4126
rect 9600 4078 9628 4236
rect 9680 4218 9732 4224
rect 9968 4154 9996 5222
rect 10784 5170 10836 5176
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 10060 4826 10088 5034
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9968 4126 10088 4154
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8588 3194 8616 3470
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7470 54 7604 82
rect 9586 82 9642 480
rect 9692 82 9720 3334
rect 9968 3194 9996 3538
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10060 2514 10088 4126
rect 10152 4010 10180 4966
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10796 4758 10824 5170
rect 11532 5030 11560 5306
rect 12176 5302 12204 5782
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12452 5137 12480 5170
rect 12438 5128 12494 5137
rect 12438 5063 12494 5072
rect 12624 5092 12676 5098
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 10784 4752 10836 4758
rect 11532 4729 11560 4966
rect 12452 4826 12480 5063
rect 12624 5034 12676 5040
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12636 4758 12664 5034
rect 12624 4752 12676 4758
rect 10784 4694 10836 4700
rect 11518 4720 11574 4729
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10428 4282 10456 4558
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10796 3602 10824 4694
rect 12624 4694 12676 4700
rect 12728 4690 12756 6326
rect 11518 4655 11574 4664
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12728 4282 12756 4626
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 12820 2650 12848 8774
rect 12912 8294 12940 11494
rect 13188 10198 13216 11562
rect 13280 11558 13308 12242
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13556 11218 13584 12650
rect 13832 12306 13860 12718
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11898 13860 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13924 11286 13952 16748
rect 14004 16730 14056 16736
rect 14660 15162 14688 23530
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 15936 23316 15988 23322
rect 15936 23258 15988 23264
rect 15474 23216 15530 23225
rect 15474 23151 15476 23160
rect 15528 23151 15530 23160
rect 15476 23122 15528 23128
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15016 22500 15068 22506
rect 15016 22442 15068 22448
rect 15028 22234 15056 22442
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 15396 22166 15424 22918
rect 15488 22778 15516 23122
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15764 22506 15792 22918
rect 15948 22642 15976 23258
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15752 22500 15804 22506
rect 15752 22442 15804 22448
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15384 22160 15436 22166
rect 15384 22102 15436 22108
rect 15476 22160 15528 22166
rect 15476 22102 15528 22108
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15396 21690 15424 22102
rect 15488 22030 15516 22102
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15488 21690 15516 21966
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 14832 21412 14884 21418
rect 14832 21354 14884 21360
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 14844 20806 14872 21354
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15580 21078 15608 21286
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15568 21072 15620 21078
rect 15568 21014 15620 21020
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15396 20330 15424 20878
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15488 20262 15516 21014
rect 15672 20942 15700 21354
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 14844 19514 14872 20198
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15304 18970 15332 19790
rect 15396 19242 15424 19926
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15580 19242 15608 19314
rect 15384 19236 15436 19242
rect 15384 19178 15436 19184
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15580 19145 15608 19178
rect 15566 19136 15622 19145
rect 15566 19071 15622 19080
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15764 18766 15792 22170
rect 15856 21962 15884 22374
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 16040 21690 16068 23462
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 16224 22642 16252 22986
rect 16212 22636 16264 22642
rect 16132 22596 16212 22624
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 16132 19122 16160 22596
rect 16212 22578 16264 22584
rect 16316 20466 16344 23530
rect 16960 23322 16988 23530
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 17236 20602 17264 20946
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 18616 20505 18644 21830
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 18602 20496 18658 20505
rect 16304 20460 16356 20466
rect 18602 20431 18658 20440
rect 16304 20402 16356 20408
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 17592 20324 17644 20330
rect 17592 20266 17644 20272
rect 16408 19718 16436 20266
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 17144 19514 17172 19926
rect 17604 19854 17632 20266
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16040 19094 16160 19122
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 16658 14872 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15488 17882 15516 18702
rect 15948 18290 15976 18838
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 17882 15792 18022
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15488 15978 15516 16934
rect 15764 16726 15792 17070
rect 16040 16794 16068 19094
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16132 18358 16160 18906
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 16132 18086 16160 18294
rect 16224 18290 16252 18702
rect 16316 18630 16344 19246
rect 17512 19174 17540 19790
rect 18708 19718 18736 19858
rect 19996 19825 20024 24006
rect 20088 22778 20116 27520
rect 21836 23866 21864 27520
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 23584 23769 23612 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24674 24848 24730 24857
rect 24674 24783 24730 24792
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 23570 23760 23626 23769
rect 23570 23695 23626 23704
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 19982 19816 20038 19825
rect 19982 19751 20038 19760
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 19514 18736 19654
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16132 17746 16160 18022
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 16132 17202 16160 17682
rect 16224 17338 16252 18226
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17236 17338 17264 17682
rect 17512 17377 17540 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17498 17368 17554 17377
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 17224 17332 17276 17338
rect 17498 17303 17554 17312
rect 17224 17274 17276 17280
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 17224 17128 17276 17134
rect 17314 17096 17370 17105
rect 17276 17076 17314 17082
rect 17224 17070 17314 17076
rect 17236 17054 17314 17070
rect 17314 17031 17370 17040
rect 17604 16998 17632 17682
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15752 16720 15804 16726
rect 15752 16662 15804 16668
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15672 16114 15700 16526
rect 15764 16250 15792 16662
rect 16040 16250 16068 16730
rect 17604 16561 17632 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 17590 16552 17646 16561
rect 17590 16487 17646 16496
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 18432 16153 18460 16390
rect 18418 16144 18474 16153
rect 15660 16108 15712 16114
rect 18418 16079 18474 16088
rect 15660 16050 15712 16056
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 14844 15706 14872 15914
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 15672 15570 15700 16050
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 16316 15162 16344 15506
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16684 14482 16712 15302
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16868 14521 16896 14554
rect 16854 14512 16910 14521
rect 16672 14476 16724 14482
rect 16854 14447 16910 14456
rect 16672 14418 16724 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 16684 14074 16712 14418
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 18616 12345 18644 13126
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 18602 12336 18658 12345
rect 18602 12271 18658 12280
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13924 10810 13952 11222
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14016 10674 14044 12174
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 14384 11694 14412 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15856 11762 15884 12038
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 14372 11688 14424 11694
rect 15660 11688 15712 11694
rect 14372 11630 14424 11636
rect 15382 11656 15438 11665
rect 14384 11354 14412 11630
rect 15660 11630 15712 11636
rect 15382 11591 15438 11600
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10198 14044 10610
rect 14292 10266 14320 11154
rect 15396 11150 15424 11591
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15488 10810 15516 11222
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 13188 9722 13216 10134
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13372 9654 13400 9998
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 14384 8634 14412 10542
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 10198 15332 10406
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 10134
rect 15580 9722 15608 11494
rect 15672 10810 15700 11630
rect 15856 11354 15884 11698
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15672 10470 15700 10746
rect 15764 10724 15792 11086
rect 15844 10736 15896 10742
rect 15764 10696 15844 10724
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15660 10056 15712 10062
rect 15764 10044 15792 10696
rect 15844 10678 15896 10684
rect 16224 10198 16252 11698
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10674 16344 10950
rect 16960 10810 16988 11018
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 15712 10016 15792 10044
rect 15660 9998 15712 10004
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15304 9518 15332 9658
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15672 9178 15700 9998
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 7342 12940 8230
rect 13372 8090 13400 8366
rect 14384 8362 14412 8570
rect 14476 8498 14504 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15672 8090 15700 8298
rect 13360 8084 13412 8090
rect 15660 8084 15712 8090
rect 13360 8026 13412 8032
rect 15580 8044 15660 8072
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 13280 7546 13308 7890
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13556 6390 13584 6870
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6390 14044 6666
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14108 5914 14136 6734
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5370 13676 5510
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13648 4282 13676 5306
rect 13740 5302 13768 5714
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 14108 5234 14136 5850
rect 14200 5778 14228 7210
rect 14292 6866 14320 7482
rect 14384 7342 14412 7686
rect 14476 7546 14504 7890
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 15580 7478 15608 8044
rect 15660 8026 15712 8032
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15672 7546 15700 7822
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 5914 14780 6258
rect 14844 6186 14872 6394
rect 15396 6322 15424 6938
rect 15580 6458 15608 7414
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15948 6866 15976 7278
rect 16224 6905 16252 7686
rect 16210 6896 16266 6905
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15936 6860 15988 6866
rect 16210 6831 16266 6840
rect 15936 6802 15988 6808
rect 15672 6458 15700 6802
rect 15948 6458 15976 6802
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 15580 5914 15608 6394
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15580 5370 15608 5850
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14476 5098 14504 5306
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 15396 4690 15424 5170
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15396 4282 15424 4626
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 13648 4078 13676 4218
rect 15672 4146 15700 4966
rect 15948 4758 15976 5034
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 15764 3602 15792 4422
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 16224 3194 16252 3538
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16316 2650 16344 10610
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17052 9722 17080 10066
rect 18970 10024 19026 10033
rect 18892 9994 18970 10010
rect 18880 9988 18970 9994
rect 18932 9982 18970 9988
rect 18970 9959 19026 9968
rect 18880 9930 18932 9936
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 22112 6730 22140 22918
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23216 7546 23244 7890
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 23308 6322 23336 23462
rect 24688 23186 24716 24783
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25148 23866 25176 24210
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25332 23225 25360 27520
rect 25502 26480 25558 26489
rect 25502 26415 25558 26424
rect 25516 23798 25544 26415
rect 27080 23866 27108 27520
rect 27068 23860 27120 23866
rect 27068 23802 27120 23808
rect 25504 23792 25556 23798
rect 25504 23734 25556 23740
rect 25318 23216 25374 23225
rect 24676 23180 24728 23186
rect 25318 23151 25374 23160
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23122
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24674 22672 24730 22681
rect 24674 22607 24730 22616
rect 24688 22098 24716 22607
rect 24676 22092 24728 22098
rect 24676 22034 24728 22040
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21690 24716 22034
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24674 20904 24730 20913
rect 24674 20839 24730 20848
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 19922 24716 20839
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23400 9654 23428 19654
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 19514 24716 19858
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 25042 19000 25098 19009
rect 25042 18935 25098 18944
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24030 17368 24086 17377
rect 24289 17360 24585 17380
rect 24766 17368 24822 17377
rect 24030 17303 24086 17312
rect 24766 17303 24822 17312
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23400 8634 23428 8910
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23492 8362 23520 9318
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23938 6896 23994 6905
rect 23938 6831 23940 6840
rect 23992 6831 23994 6840
rect 23940 6802 23992 6808
rect 23952 6458 23980 6802
rect 24044 6730 24072 17303
rect 24780 17270 24808 17303
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24504 17105 24532 17138
rect 24490 17096 24546 17105
rect 24490 17031 24546 17040
rect 25056 16658 25084 18935
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16250 24716 16594
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24950 15192 25006 15201
rect 24950 15127 25006 15136
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24214 12336 24270 12345
rect 24214 12271 24270 12280
rect 24228 11694 24256 12271
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24964 10810 24992 15127
rect 27618 12064 27674 12073
rect 27618 11999 27674 12008
rect 27632 11898 27660 11999
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 24596 10033 24624 10066
rect 24582 10024 24638 10033
rect 24638 9982 24716 10010
rect 24582 9959 24638 9968
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9722 24716 9982
rect 25240 9722 25268 10406
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27632 10169 27660 10202
rect 27618 10160 27674 10169
rect 27618 10095 27674 10104
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 24136 9110 24164 9318
rect 24596 9110 24624 9454
rect 24124 9104 24176 9110
rect 24124 9046 24176 9052
rect 24584 9104 24636 9110
rect 24636 9064 24716 9092
rect 24584 9046 24636 9052
rect 24136 8634 24164 9046
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24688 8566 24716 9064
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24872 8498 24900 8774
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24872 8022 24900 8434
rect 27618 8256 27674 8265
rect 27618 8191 27674 8200
rect 27632 8090 27660 8191
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 24860 8016 24912 8022
rect 24860 7958 24912 7964
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7410 24164 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24688 7206 24716 7958
rect 24768 7812 24820 7818
rect 24768 7754 24820 7760
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24136 7002 24164 7142
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 24504 6866 24532 7142
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24032 6724 24084 6730
rect 24032 6666 24084 6672
rect 24780 6644 24808 7754
rect 24872 7478 24900 7958
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 24860 6656 24912 6662
rect 24780 6616 24860 6644
rect 24860 6598 24912 6604
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23848 6180 23900 6186
rect 23848 6122 23900 6128
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 5370 16896 5714
rect 18248 5710 18276 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 17880 5370 17908 5646
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 18248 5098 18276 5510
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18248 4690 18276 5034
rect 18616 5030 18644 5782
rect 23860 5778 23888 6122
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 19156 5636 19208 5642
rect 19156 5578 19208 5584
rect 19168 5234 19196 5578
rect 23860 5370 23888 5714
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24044 5370 24072 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18616 4826 18644 4966
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18708 4729 18736 4762
rect 18694 4720 18750 4729
rect 18236 4684 18288 4690
rect 18694 4655 18750 4664
rect 18236 4626 18288 4632
rect 18248 4282 18276 4626
rect 19168 4282 19196 5170
rect 24044 5030 24072 5306
rect 24780 5302 24808 6122
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 24228 4826 24256 5034
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19168 4078 19196 4218
rect 22940 4154 22968 4626
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4626
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 22848 4146 22968 4154
rect 22836 4140 22968 4146
rect 22888 4126 22968 4140
rect 22836 4082 22888 4088
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 22848 3942 22876 4082
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 19168 3602 19196 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 11428 2372 11480 2378
rect 11428 2314 11480 2320
rect 9586 54 9720 82
rect 11440 82 11468 2314
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 11702 82 11758 480
rect 11440 54 11758 82
rect 13740 82 13768 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 13910 82 13966 480
rect 13740 54 13966 82
rect 15672 82 15700 2246
rect 16026 82 16082 480
rect 15672 54 16082 82
rect 7470 0 7526 54
rect 9586 0 9642 54
rect 11702 0 11758 54
rect 13910 0 13966 54
rect 16026 0 16082 54
rect 18234 82 18290 480
rect 18340 82 18368 3334
rect 19168 3194 19196 3538
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 18234 54 18368 82
rect 20180 82 20208 3334
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 20350 82 20406 480
rect 20180 54 20406 82
rect 22112 82 22140 2246
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 22466 82 22522 480
rect 22112 54 22522 82
rect 18234 0 18290 54
rect 20350 0 20406 54
rect 22466 0 22522 54
rect 24674 82 24730 480
rect 24780 82 24808 3878
rect 24872 2650 24900 6598
rect 25516 6390 25544 6802
rect 27618 6488 27674 6497
rect 27618 6423 27674 6432
rect 27632 6390 27660 6423
rect 25504 6384 25556 6390
rect 25504 6326 25556 6332
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27632 4593 27660 4626
rect 27618 4584 27674 4593
rect 27618 4519 27674 4528
rect 27618 2680 27674 2689
rect 24860 2644 24912 2650
rect 27618 2615 27674 2624
rect 24860 2586 24912 2592
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 24674 54 24808 82
rect 26528 82 26556 2246
rect 27632 1601 27660 2615
rect 27618 1592 27674 1601
rect 27618 1527 27674 1536
rect 26790 82 26846 480
rect 26528 54 26846 82
rect 24674 0 24730 54
rect 26790 0 26846 54
<< via2 >>
rect 1030 26560 1086 26616
rect 2226 25064 2282 25120
rect 3330 23432 3386 23488
rect 1122 12552 1178 12608
rect 110 11600 166 11656
rect 202 7112 258 7168
rect 110 5344 166 5400
rect 1582 20304 1638 20360
rect 1306 18808 1362 18864
rect 4434 23160 4490 23216
rect 3698 23024 3754 23080
rect 3882 21936 3938 21992
rect 3514 19216 3570 19272
rect 1858 17176 1914 17232
rect 4434 19760 4490 19816
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 1582 9696 1638 9752
rect 1582 8744 1638 8800
rect 2042 8372 2044 8392
rect 2044 8372 2096 8392
rect 2096 8372 2098 8392
rect 2042 8336 2098 8372
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 6182 20440 6238 20496
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5262 16496 5318 16552
rect 5078 15680 5134 15736
rect 4894 14184 4950 14240
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6826 19216 6882 19272
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6918 16088 6974 16144
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 8482 16088 8538 16144
rect 7838 13912 7894 13968
rect 8758 16496 8814 16552
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 13542 23024 13598 23080
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 8942 17584 8998 17640
rect 8206 13776 8262 13832
rect 8850 13776 8906 13832
rect 9494 13912 9550 13968
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 110 3712 166 3768
rect 2134 5072 2190 5128
rect 1950 1264 2006 1320
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7010 2760 7066 2816
rect 6550 1536 6606 1592
rect 8942 11600 8998 11656
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9862 8336 9918 8392
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 12346 19080 12402 19136
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 17222 23704 17278 23760
rect 14554 23160 14610 23216
rect 14278 17584 14334 17640
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10966 5616 11022 5672
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 12438 5072 12494 5128
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11518 4664 11574 4720
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 15474 23180 15530 23216
rect 15474 23160 15476 23180
rect 15476 23160 15528 23180
rect 15528 23160 15530 23180
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15566 19080 15622 19136
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 18602 20440 18658 20496
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24792 24730 24848
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 23570 23704 23626 23760
rect 19982 19760 20038 19816
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 17498 17312 17554 17368
rect 17314 17040 17370 17096
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 17590 16496 17646 16552
rect 18418 16088 18474 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 16854 14456 16910 14512
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 18602 12280 18658 12336
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15382 11600 15438 11656
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 16210 6840 16266 6896
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 18970 9968 19026 10024
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 25502 26424 25558 26480
rect 25318 23160 25374 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24674 22616 24730 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24674 20848 24730 20904
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 25042 18944 25098 19000
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24030 17312 24086 17368
rect 24766 17312 24822 17368
rect 23938 6860 23994 6896
rect 23938 6840 23940 6860
rect 23940 6840 23992 6860
rect 23992 6840 23994 6860
rect 24490 17040 24546 17096
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24950 15136 25006 15192
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24214 12280 24270 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 27618 12008 27674 12064
rect 24582 9968 24638 10024
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 27618 10104 27674 10160
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 27618 8200 27674 8256
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 18694 4664 18750 4720
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27618 6432 27674 6488
rect 27618 4528 27674 4584
rect 27618 2624 27674 2680
rect 27618 1536 27674 1592
<< metal3 >>
rect 0 27072 480 27192
rect 62 26618 122 27072
rect 27520 26936 28000 27056
rect 1025 26618 1091 26621
rect 62 26616 1091 26618
rect 62 26560 1030 26616
rect 1086 26560 1091 26616
rect 62 26558 1091 26560
rect 1025 26555 1091 26558
rect 25497 26482 25563 26485
rect 27662 26482 27722 26936
rect 25497 26480 27722 26482
rect 25497 26424 25502 26480
rect 25558 26424 27722 26480
rect 25497 26422 27722 26424
rect 25497 26419 25563 26422
rect 0 25576 480 25696
rect 10277 25600 10597 25601
rect 62 25122 122 25576
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 2221 25122 2287 25125
rect 62 25120 2287 25122
rect 62 25064 2226 25120
rect 2282 25064 2287 25120
rect 62 25062 2287 25064
rect 2221 25059 2287 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 27520 25032 28000 25152
rect 24277 24991 24597 24992
rect 24669 24850 24735 24853
rect 27662 24850 27722 25032
rect 24669 24848 27722 24850
rect 24669 24792 24674 24848
rect 24730 24792 27722 24848
rect 24669 24790 27722 24792
rect 24669 24787 24735 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 23944 480 24064
rect 5610 23968 5930 23969
rect 62 23490 122 23944
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 17217 23762 17283 23765
rect 23565 23762 23631 23765
rect 17217 23760 23631 23762
rect 17217 23704 17222 23760
rect 17278 23704 23570 23760
rect 23626 23704 23631 23760
rect 17217 23702 23631 23704
rect 17217 23699 17283 23702
rect 23565 23699 23631 23702
rect 3325 23490 3391 23493
rect 62 23488 3391 23490
rect 62 23432 3330 23488
rect 3386 23432 3391 23488
rect 62 23430 3391 23432
rect 3325 23427 3391 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 4429 23218 4495 23221
rect 14549 23218 14615 23221
rect 4429 23216 14615 23218
rect 4429 23160 4434 23216
rect 4490 23160 14554 23216
rect 14610 23160 14615 23216
rect 4429 23158 14615 23160
rect 4429 23155 4495 23158
rect 14549 23155 14615 23158
rect 15469 23218 15535 23221
rect 25313 23218 25379 23221
rect 15469 23216 25379 23218
rect 15469 23160 15474 23216
rect 15530 23160 25318 23216
rect 25374 23160 25379 23216
rect 15469 23158 25379 23160
rect 15469 23155 15535 23158
rect 25313 23155 25379 23158
rect 27520 23128 28000 23248
rect 3693 23082 3759 23085
rect 13537 23082 13603 23085
rect 3693 23080 13603 23082
rect 3693 23024 3698 23080
rect 3754 23024 13542 23080
rect 13598 23024 13603 23080
rect 3693 23022 13603 23024
rect 3693 23019 3759 23022
rect 13537 23019 13603 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 24669 22674 24735 22677
rect 27662 22674 27722 23128
rect 24669 22672 27722 22674
rect 24669 22616 24674 22672
rect 24730 22616 27722 22672
rect 24669 22614 27722 22616
rect 24669 22611 24735 22614
rect 0 22448 480 22568
rect 62 21994 122 22448
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 3877 21994 3943 21997
rect 62 21992 3943 21994
rect 62 21936 3882 21992
rect 3938 21936 3943 21992
rect 62 21934 3943 21936
rect 3877 21931 3943 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 27520 21360 28000 21480
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 20816 480 20936
rect 24669 20906 24735 20909
rect 27662 20906 27722 21360
rect 24669 20904 27722 20906
rect 24669 20848 24674 20904
rect 24730 20848 27722 20904
rect 24669 20846 27722 20848
rect 24669 20843 24735 20846
rect 62 20362 122 20816
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 6177 20498 6243 20501
rect 18597 20498 18663 20501
rect 6177 20496 18663 20498
rect 6177 20440 6182 20496
rect 6238 20440 18602 20496
rect 18658 20440 18663 20496
rect 6177 20438 18663 20440
rect 6177 20435 6243 20438
rect 18597 20435 18663 20438
rect 1577 20362 1643 20365
rect 62 20360 1643 20362
rect 62 20304 1582 20360
rect 1638 20304 1643 20360
rect 62 20302 1643 20304
rect 1577 20299 1643 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 4429 19818 4495 19821
rect 19977 19818 20043 19821
rect 4429 19816 20043 19818
rect 4429 19760 4434 19816
rect 4490 19760 19982 19816
rect 20038 19760 20043 19816
rect 4429 19758 20043 19760
rect 4429 19755 4495 19758
rect 19977 19755 20043 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19456 28000 19576
rect 0 19320 480 19440
rect 62 18866 122 19320
rect 3509 19274 3575 19277
rect 6821 19274 6887 19277
rect 3509 19272 6887 19274
rect 3509 19216 3514 19272
rect 3570 19216 6826 19272
rect 6882 19216 6887 19272
rect 3509 19214 6887 19216
rect 3509 19211 3575 19214
rect 6821 19211 6887 19214
rect 12341 19138 12407 19141
rect 15561 19138 15627 19141
rect 12341 19136 15627 19138
rect 12341 19080 12346 19136
rect 12402 19080 15566 19136
rect 15622 19080 15627 19136
rect 12341 19078 15627 19080
rect 12341 19075 12407 19078
rect 15561 19075 15627 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 25037 19002 25103 19005
rect 27662 19002 27722 19456
rect 25037 19000 27722 19002
rect 25037 18944 25042 19000
rect 25098 18944 27722 19000
rect 25037 18942 27722 18944
rect 25037 18939 25103 18942
rect 1301 18866 1367 18869
rect 62 18864 1367 18866
rect 62 18808 1306 18864
rect 1362 18808 1367 18864
rect 62 18806 1367 18808
rect 1301 18803 1367 18806
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 0 17688 480 17808
rect 62 17234 122 17688
rect 8937 17642 9003 17645
rect 14273 17642 14339 17645
rect 8937 17640 14339 17642
rect 8937 17584 8942 17640
rect 8998 17584 14278 17640
rect 14334 17584 14339 17640
rect 8937 17582 14339 17584
rect 8937 17579 9003 17582
rect 14273 17579 14339 17582
rect 27520 17552 28000 17672
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 17493 17370 17559 17373
rect 24025 17370 24091 17373
rect 17493 17368 24091 17370
rect 17493 17312 17498 17368
rect 17554 17312 24030 17368
rect 24086 17312 24091 17368
rect 17493 17310 24091 17312
rect 17493 17307 17559 17310
rect 24025 17307 24091 17310
rect 24761 17370 24827 17373
rect 27662 17370 27722 17552
rect 24761 17368 27722 17370
rect 24761 17312 24766 17368
rect 24822 17312 27722 17368
rect 24761 17310 27722 17312
rect 24761 17307 24827 17310
rect 1853 17234 1919 17237
rect 62 17232 1919 17234
rect 62 17176 1858 17232
rect 1914 17176 1919 17232
rect 62 17174 1919 17176
rect 1853 17171 1919 17174
rect 17309 17098 17375 17101
rect 24485 17098 24551 17101
rect 17309 17096 24551 17098
rect 17309 17040 17314 17096
rect 17370 17040 24490 17096
rect 24546 17040 24551 17096
rect 17309 17038 24551 17040
rect 17309 17035 17375 17038
rect 24485 17035 24551 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5257 16554 5323 16557
rect 8753 16554 8819 16557
rect 17585 16554 17651 16557
rect 5257 16552 17651 16554
rect 5257 16496 5262 16552
rect 5318 16496 8758 16552
rect 8814 16496 17590 16552
rect 17646 16496 17651 16552
rect 5257 16494 17651 16496
rect 5257 16491 5323 16494
rect 8753 16491 8819 16494
rect 17585 16491 17651 16494
rect 5610 16352 5930 16353
rect 0 16192 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 62 15738 122 16192
rect 6913 16146 6979 16149
rect 8477 16146 8543 16149
rect 18413 16146 18479 16149
rect 6913 16144 18479 16146
rect 6913 16088 6918 16144
rect 6974 16088 8482 16144
rect 8538 16088 18418 16144
rect 18474 16088 18479 16144
rect 6913 16086 18479 16088
rect 6913 16083 6979 16086
rect 8477 16083 8543 16086
rect 18413 16083 18479 16086
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 5073 15738 5139 15741
rect 62 15736 5139 15738
rect 62 15680 5078 15736
rect 5134 15680 5139 15736
rect 62 15678 5139 15680
rect 5073 15675 5139 15678
rect 27520 15648 28000 15768
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 24945 15194 25011 15197
rect 27662 15194 27722 15648
rect 24945 15192 27722 15194
rect 24945 15136 24950 15192
rect 25006 15136 27722 15192
rect 24945 15134 27722 15136
rect 24945 15131 25011 15134
rect 0 14696 480 14816
rect 10277 14720 10597 14721
rect 62 14242 122 14696
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 16849 14514 16915 14517
rect 16849 14512 27722 14514
rect 16849 14456 16854 14512
rect 16910 14456 27722 14512
rect 16849 14454 27722 14456
rect 16849 14451 16915 14454
rect 4889 14242 4955 14245
rect 62 14240 4955 14242
rect 62 14184 4894 14240
rect 4950 14184 4955 14240
rect 62 14182 4955 14184
rect 4889 14179 4955 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27662 14000 27722 14454
rect 7833 13970 7899 13973
rect 9489 13970 9555 13973
rect 7833 13968 9555 13970
rect 7833 13912 7838 13968
rect 7894 13912 9494 13968
rect 9550 13912 9555 13968
rect 7833 13910 9555 13912
rect 7833 13907 7899 13910
rect 9489 13907 9555 13910
rect 27520 13880 28000 14000
rect 8201 13834 8267 13837
rect 8845 13834 8911 13837
rect 8201 13832 8911 13834
rect 8201 13776 8206 13832
rect 8262 13776 8850 13832
rect 8906 13776 8911 13832
rect 8201 13774 8911 13776
rect 8201 13771 8267 13774
rect 8845 13771 8911 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 0 13064 480 13184
rect 5610 13088 5930 13089
rect 62 12610 122 13064
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 1117 12610 1183 12613
rect 62 12608 1183 12610
rect 62 12552 1122 12608
rect 1178 12552 1183 12608
rect 62 12550 1183 12552
rect 1117 12547 1183 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 18597 12338 18663 12341
rect 24209 12338 24275 12341
rect 18597 12336 24275 12338
rect 18597 12280 18602 12336
rect 18658 12280 24214 12336
rect 24270 12280 24275 12336
rect 18597 12278 24275 12280
rect 18597 12275 18663 12278
rect 24209 12275 24275 12278
rect 27520 12064 28000 12096
rect 27520 12008 27618 12064
rect 27674 12008 28000 12064
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 27520 11976 28000 12008
rect 24277 11935 24597 11936
rect 0 11656 480 11688
rect 0 11600 110 11656
rect 166 11600 480 11656
rect 0 11568 480 11600
rect 8937 11658 9003 11661
rect 15377 11658 15443 11661
rect 8937 11656 15443 11658
rect 8937 11600 8942 11656
rect 8998 11600 15382 11656
rect 15438 11600 15443 11656
rect 8937 11598 15443 11600
rect 8937 11595 9003 11598
rect 15377 11595 15443 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 27520 10160 28000 10192
rect 27520 10104 27618 10160
rect 27674 10104 28000 10160
rect 27520 10072 28000 10104
rect 0 9936 480 10056
rect 18965 10026 19031 10029
rect 24577 10026 24643 10029
rect 18965 10024 24643 10026
rect 18965 9968 18970 10024
rect 19026 9968 24582 10024
rect 24638 9968 24643 10024
rect 18965 9966 24643 9968
rect 18965 9963 19031 9966
rect 24577 9963 24643 9966
rect 62 9754 122 9936
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1577 9754 1643 9757
rect 62 9752 1643 9754
rect 62 9696 1582 9752
rect 1638 9696 1643 9752
rect 62 9694 1643 9696
rect 1577 9691 1643 9694
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 54 8740 60 8804
rect 124 8802 130 8804
rect 1577 8802 1643 8805
rect 124 8800 1643 8802
rect 124 8744 1582 8800
rect 1638 8744 1643 8800
rect 124 8742 1643 8744
rect 124 8740 130 8742
rect 1577 8739 1643 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 0 8532 480 8560
rect 0 8468 60 8532
rect 124 8468 480 8532
rect 0 8440 480 8468
rect 2037 8394 2103 8397
rect 9857 8394 9923 8397
rect 2037 8392 9923 8394
rect 2037 8336 2042 8392
rect 2098 8336 9862 8392
rect 9918 8336 9923 8392
rect 2037 8334 9923 8336
rect 2037 8331 2103 8334
rect 9857 8331 9923 8334
rect 27520 8256 28000 8288
rect 27520 8200 27618 8256
rect 27674 8200 28000 8256
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8200
rect 19610 8127 19930 8128
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 197 7170 263 7173
rect 62 7168 263 7170
rect 62 7112 202 7168
rect 258 7112 263 7168
rect 62 7110 263 7112
rect 62 6928 122 7110
rect 197 7107 263 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6808 480 6928
rect 16205 6898 16271 6901
rect 23933 6898 23999 6901
rect 16205 6896 23999 6898
rect 16205 6840 16210 6896
rect 16266 6840 23938 6896
rect 23994 6840 23999 6896
rect 16205 6838 23999 6840
rect 16205 6835 16271 6838
rect 23933 6835 23999 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 27520 6488 28000 6520
rect 27520 6432 27618 6488
rect 27674 6432 28000 6488
rect 27520 6400 28000 6432
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 10961 5674 11027 5677
rect 27654 5674 27660 5676
rect 10961 5672 27660 5674
rect 10961 5616 10966 5672
rect 11022 5616 27660 5672
rect 10961 5614 27660 5616
rect 10961 5611 11027 5614
rect 27654 5612 27660 5614
rect 27724 5612 27730 5676
rect 5610 5472 5930 5473
rect 0 5400 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5344 110 5400
rect 166 5344 480 5400
rect 0 5312 480 5344
rect 2129 5130 2195 5133
rect 12433 5130 12499 5133
rect 2129 5128 12499 5130
rect 2129 5072 2134 5128
rect 2190 5072 12438 5128
rect 12494 5072 12499 5128
rect 2129 5070 12499 5072
rect 2129 5067 2195 5070
rect 12433 5067 12499 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 11513 4722 11579 4725
rect 18689 4722 18755 4725
rect 11513 4720 18755 4722
rect 11513 4664 11518 4720
rect 11574 4664 18694 4720
rect 18750 4664 18755 4720
rect 11513 4662 18755 4664
rect 11513 4659 11579 4662
rect 18689 4659 18755 4662
rect 27520 4584 28000 4616
rect 27520 4528 27618 4584
rect 27674 4528 28000 4584
rect 27520 4496 28000 4528
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 0 3768 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3712 110 3768
rect 166 3712 480 3768
rect 0 3680 480 3712
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 7005 2818 7071 2821
rect 62 2816 7071 2818
rect 62 2760 7010 2816
rect 7066 2760 7071 2816
rect 62 2758 7071 2760
rect 62 2304 122 2758
rect 7005 2755 7071 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 27520 2680 28000 2712
rect 27520 2624 27618 2680
rect 27674 2624 28000 2680
rect 27520 2592 28000 2624
rect 0 2184 480 2304
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6545 1594 6611 1597
rect 27613 1594 27679 1597
rect 6545 1592 27679 1594
rect 6545 1536 6550 1592
rect 6606 1536 27618 1592
rect 27674 1536 27679 1592
rect 6545 1534 27679 1536
rect 6545 1531 6611 1534
rect 27613 1531 27679 1534
rect 1945 1322 2011 1325
rect 62 1320 2011 1322
rect 62 1264 1950 1320
rect 2006 1264 2011 1320
rect 62 1262 2011 1264
rect 62 808 122 1262
rect 1945 1259 2011 1262
rect 27520 916 28000 944
rect 27520 852 27660 916
rect 27724 852 28000 916
rect 27520 824 28000 852
rect 0 688 480 808
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 60 8740 124 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 60 8468 124 8532
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 27660 5612 27724 5676
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 27660 852 27724 916
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 59 8804 125 8805
rect 59 8740 60 8804
rect 124 8740 125 8804
rect 59 8739 125 8740
rect 62 8533 122 8739
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 59 8532 125 8533
rect 59 8468 60 8532
rect 124 8468 125 8532
rect 59 8467 125 8468
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 27659 5676 27725 5677
rect 27659 5612 27660 5676
rect 27724 5612 27725 5676
rect 27659 5611 27725 5612
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 27662 917 27722 5611
rect 27659 916 27725 917
rect 27659 852 27660 916
rect 27724 852 27725 916
rect 27659 851 27725 852
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__200__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_82
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_90
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _199_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_110
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_122
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_132
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_140 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_154
timestamp 1586364061
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_163
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_166
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_184
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_234
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_242
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 16192 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_162
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_192
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_200
timestamp 1586364061
transform 1 0 19504 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_212
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_6
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_82
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _111_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _093_
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_188
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_237
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _186_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_134
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 774 592
use scs8hd_conb_1  _195_
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_157
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_194
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_26
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_50
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_188
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_271
timestamp 1586364061
transform 1 0 26036 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use scs8hd_nand2_4  _126_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_12
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_20
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_24
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_28
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 774 592
use scs8hd_nor2_4  _165_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__D
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_111
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__C
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_115
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_137
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_177
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_189
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_198
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_241
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_237
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_245
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _102_
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_255
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_262
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_274
timestamp 1586364061
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_or2_4  _122_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 682 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_13
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_25
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_67
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_71
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_or4_4  _136_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_118
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_175
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_8  _096_
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_256
timestamp 1586364061
transform 1 0 24656 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__173__C
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_49
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 590 592
use scs8hd_nand2_4  _148_
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__D
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 130 592
use scs8hd_inv_8  _112_
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 406 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_238
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_260
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_264
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_268
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_or4_4  _173_
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_242
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_67
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _164_
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_102
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_137
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_262
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 682 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_99
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_103
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 406 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_235
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 130 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_256
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_260
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_35
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_109
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_8  _105_
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_165
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_176
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_188
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_200
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_153
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_157
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_170
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_253
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_8  _115_
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__D
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_119
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_123
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_198
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_6
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_70
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _170_
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _116_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_111
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _106_
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_151
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 774 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_253
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_71
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _155_
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_161
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_185
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_209
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _119_
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_40
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_55
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_44
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__D
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use scs8hd_or4_4  _158_
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 866 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_78
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_82
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_78
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_99
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_112
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_147
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_nor3_4  _176_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_32
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_76
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _167_
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_111
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_115
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_11
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _107_
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_173
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_185
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_197
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_209
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_84
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_106
timestamp 1586364061
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_164
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 590 592
use scs8hd_inv_8  _120_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_or4_4  _161_
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_101
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__C
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__D
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_136
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_157
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_180
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_6
timestamp 1586364061
transform 1 0 1656 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_10
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use scs8hd_nor3_4  _177_
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use scs8hd_or4_4  _127_
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_88
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_108
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 406 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_157
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_161
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_165
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_9
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_26
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 4140 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_37
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_nor3_4  _175_
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 1234 592
use scs8hd_nor3_4  _174_
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 406 592
use scs8hd_inv_8  _118_
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_or4_4  _145_
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_75
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_81
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_88
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_85
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_or4_4  _152_
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__D
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use scs8hd_or4_4  _142_
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 866 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_119
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_145
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _086_
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_166
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_181
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_258
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_270
timestamp 1586364061
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_71
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__D
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 314 592
use scs8hd_or4_4  _133_
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__C
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_122
timestamp 1586364061
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _097_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_204
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_29
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _117_
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_88
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 12512 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_133
timestamp 1586364061
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_137
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_169
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_173
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_181
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_22
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_26
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_8  _100_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_54
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_66
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_4  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_8  _109_
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_110
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 590 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_164
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 16928 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_168
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_175
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_199
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_12
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_48
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_52
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _099_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_60
timestamp 1586364061
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_96
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_103
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_113
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_155
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_192
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_204
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_216
timestamp 1586364061
transform 1 0 20976 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_228
timestamp 1586364061
transform 1 0 22080 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_10
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_21
timestamp 1586364061
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_25
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_37
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_50
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_67
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_6  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_112
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_133
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 20128
box -38 -48 314 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_165
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 866 592
use scs8hd_inv_8  _092_
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_258
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_270
timestamp 1586364061
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_25
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_17
timestamp 1586364061
transform 1 0 2668 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_21
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_33
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_40
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_37
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_52
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_75
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_92
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_85
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_97
timestamp 1586364061
transform 1 0 10028 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 130 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_113
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_113
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_126
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_131
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_152
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_140
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_148
timestamp 1586364061
transform 1 0 14720 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_180
timestamp 1586364061
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_192
timestamp 1586364061
transform 1 0 18768 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_204
timestamp 1586364061
transform 1 0 19872 0 -1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_212
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_20
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_24
timestamp 1586364061
transform 1 0 3312 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_36
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_40
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_52
timestamp 1586364061
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_66
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_84
timestamp 1586364061
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_97
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 406 592
use scs8hd_decap_6  FILLER_35_138
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_146
timestamp 1586364061
transform 1 0 14536 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_163
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_170
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_182
timestamp 1586364061
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_18
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 1142 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_30
timestamp 1586364061
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_37
timestamp 1586364061
transform 1 0 4508 0 -1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_62
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_66
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_72
timestamp 1586364061
transform 1 0 7728 0 -1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_107
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_1  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_8  _098_
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_128
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_258
timestamp 1586364061
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_270
timestamp 1586364061
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_18
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_22
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_29
timestamp 1586364061
transform 1 0 3772 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_33
timestamp 1586364061
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_46
timestamp 1586364061
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_50
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_58
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 774 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 7728 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_70
timestamp 1586364061
transform 1 0 7544 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_inv_8  _110_
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_inv_8  _085_
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_139
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_152
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_157
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_169
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_181
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_192
timestamp 1586364061
transform 1 0 18768 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_204
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_216
timestamp 1586364061
transform 1 0 20976 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_228
timestamp 1586364061
transform 1 0 22080 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 1932 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_11
timestamp 1586364061
transform 1 0 2116 0 -1 23392
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_17
timestamp 1586364061
transform 1 0 2668 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_21
timestamp 1586364061
transform 1 0 3036 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_29
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_36
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_39
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_50
timestamp 1586364061
transform 1 0 5704 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_62
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_38_74
timestamp 1586364061
transform 1 0 7912 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_8  _104_
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_6  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_144
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_148
timestamp 1586364061
transform 1 0 14720 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_162
timestamp 1586364061
transform 1 0 16008 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_258
timestamp 1586364061
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_270
timestamp 1586364061
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_14
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_31
timestamp 1586364061
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_35
timestamp 1586364061
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_48
timestamp 1586364061
transform 1 0 5520 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_60
timestamp 1586364061
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 774 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_76
timestamp 1586364061
transform 1 0 8096 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 130 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 9936 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_87
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_91
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_98
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_104
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_109
timestamp 1586364061
transform 1 0 11132 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_121
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_133
timestamp 1586364061
transform 1 0 13340 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_151
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_168
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_172
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_176
timestamp 1586364061
transform 1 0 17296 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_169
timestamp 1586364061
transform 1 0 16652 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_181
timestamp 1586364061
transform 1 0 17756 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_193
timestamp 1586364061
transform 1 0 18860 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_207
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_205
timestamp 1586364061
transform 1 0 19964 0 -1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_211
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_258
timestamp 1586364061
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_266
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_270
timestamp 1586364061
transform 1 0 25944 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5262 0 5318 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 688 480 808 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 2184 480 2304 6 address[2]
port 2 nsew default input
rlabel metal3 s 27520 824 28000 944 6 address[3]
port 3 nsew default input
rlabel metal2 s 7470 0 7526 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 address[5]
port 5 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[0]
port 6 nsew default input
rlabel metal2 s 846 27520 902 28000 6 chanx_right_in[1]
port 7 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_right_in[2]
port 8 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 chanx_right_in[3]
port 9 nsew default input
rlabel metal3 s 27520 6400 28000 6520 6 chanx_right_in[4]
port 10 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_right_in[5]
port 11 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[6]
port 12 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chanx_right_in[7]
port 13 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_right_in[8]
port 14 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_right_out[0]
port 15 nsew default tristate
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_out[1]
port 16 nsew default tristate
rlabel metal2 s 6090 27520 6146 28000 6 chanx_right_out[2]
port 17 nsew default tristate
rlabel metal3 s 27520 11976 28000 12096 6 chanx_right_out[3]
port 18 nsew default tristate
rlabel metal2 s 9586 0 9642 480 6 chanx_right_out[4]
port 19 nsew default tristate
rlabel metal2 s 11702 0 11758 480 6 chanx_right_out[5]
port 20 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 chanx_right_out[6]
port 21 nsew default tristate
rlabel metal2 s 7838 27520 7894 28000 6 chanx_right_out[7]
port 22 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_right_out[8]
port 23 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chany_top_in[0]
port 24 nsew default input
rlabel metal3 s 0 14696 480 14816 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chany_top_in[3]
port 27 nsew default input
rlabel metal3 s 0 17688 480 17808 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_top_in[6]
port 30 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 11334 27520 11390 28000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 15648 28000 15768 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 17552 28000 17672 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 data_in
port 42 nsew default input
rlabel metal2 s 1030 0 1086 480 6 enable
port 43 nsew default input
rlabel metal3 s 27520 21360 28000 21480 6 right_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 0 25576 480 25696 6 right_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal2 s 18326 27520 18382 28000 6 right_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal2 s 22466 0 22522 480 6 right_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal3 s 27520 19456 28000 19576 6 right_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 0 23944 480 24064 6 right_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal2 s 24674 0 24730 480 6 right_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 right_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal2 s 20074 27520 20130 28000 6 right_top_grid_pin_10_
port 52 nsew default input
rlabel metal2 s 26790 0 26846 480 6 top_left_grid_pin_11_
port 53 nsew default input
rlabel metal2 s 25318 27520 25374 28000 6 top_left_grid_pin_13_
port 54 nsew default input
rlabel metal2 s 27066 27520 27122 28000 6 top_left_grid_pin_15_
port 55 nsew default input
rlabel metal2 s 21822 27520 21878 28000 6 top_left_grid_pin_1_
port 56 nsew default input
rlabel metal3 s 0 27072 480 27192 6 top_left_grid_pin_3_
port 57 nsew default input
rlabel metal3 s 27520 23128 28000 23248 6 top_left_grid_pin_5_
port 58 nsew default input
rlabel metal2 s 23570 27520 23626 28000 6 top_left_grid_pin_7_
port 59 nsew default input
rlabel metal3 s 27520 25032 28000 25152 6 top_left_grid_pin_9_
port 60 nsew default input
rlabel metal3 s 27520 26936 28000 27056 6 top_right_grid_pin_11_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
