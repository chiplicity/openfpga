magic
tech sky130A
magscale 1 2
timestamp 1609017451
<< locali >>
rect 16129 13311 16163 13481
rect 13921 10115 13955 10217
rect 16221 9911 16255 10013
rect 10333 7735 10367 7973
rect 10425 7735 10459 7905
rect 22017 5559 22051 6817
rect 12449 3927 12483 4029
rect 19257 3383 19291 3485
rect 20637 3383 20671 3485
rect 18337 2907 18371 3077
rect 20729 2975 20763 3077
<< viali >>
rect 20453 20009 20487 20043
rect 21097 20009 21131 20043
rect 20269 19873 20303 19907
rect 20913 19873 20947 19907
rect 21005 19465 21039 19499
rect 6837 19261 6871 19295
rect 7389 19261 7423 19295
rect 19717 19261 19751 19295
rect 20269 19261 20303 19295
rect 20821 19261 20855 19295
rect 7021 19125 7055 19159
rect 19901 19125 19935 19159
rect 20453 19125 20487 19159
rect 21097 18921 21131 18955
rect 12357 18853 12391 18887
rect 16129 18853 16163 18887
rect 18521 18853 18555 18887
rect 20177 18853 20211 18887
rect 12081 18785 12115 18819
rect 15853 18785 15887 18819
rect 18245 18785 18279 18819
rect 19901 18785 19935 18819
rect 20913 18785 20947 18819
rect 21005 18377 21039 18411
rect 9689 18241 9723 18275
rect 9413 18173 9447 18207
rect 20821 18173 20855 18207
rect 21097 17833 21131 17867
rect 8309 17697 8343 17731
rect 20913 17697 20947 17731
rect 8585 17629 8619 17663
rect 18797 17289 18831 17323
rect 21005 17289 21039 17323
rect 11529 17153 11563 17187
rect 20177 17153 20211 17187
rect 11253 17085 11287 17119
rect 18613 17085 18647 17119
rect 19901 17085 19935 17119
rect 20821 17085 20855 17119
rect 21097 16745 21131 16779
rect 17969 16677 18003 16711
rect 17693 16609 17727 16643
rect 20913 16609 20947 16643
rect 21005 16201 21039 16235
rect 20177 16065 20211 16099
rect 19901 15997 19935 16031
rect 20821 15997 20855 16031
rect 20453 15657 20487 15691
rect 21097 15657 21131 15691
rect 14657 15589 14691 15623
rect 14381 15521 14415 15555
rect 20269 15521 20303 15555
rect 20913 15521 20947 15555
rect 21005 15113 21039 15147
rect 11897 14977 11931 15011
rect 11621 14909 11655 14943
rect 20821 14909 20855 14943
rect 20545 14569 20579 14603
rect 21097 14569 21131 14603
rect 9965 14501 9999 14535
rect 8769 14433 8803 14467
rect 9689 14433 9723 14467
rect 20913 14433 20947 14467
rect 9045 14365 9079 14399
rect 20729 13889 20763 13923
rect 11161 13821 11195 13855
rect 11437 13821 11471 13855
rect 20361 13821 20395 13855
rect 16129 13481 16163 13515
rect 20453 13481 20487 13515
rect 21097 13481 21131 13515
rect 13553 13345 13587 13379
rect 13829 13345 13863 13379
rect 16488 13413 16522 13447
rect 17969 13413 18003 13447
rect 20269 13345 20303 13379
rect 20913 13345 20947 13379
rect 16129 13277 16163 13311
rect 16221 13277 16255 13311
rect 17601 13141 17635 13175
rect 19993 13141 20027 13175
rect 21281 12937 21315 12971
rect 20545 12801 20579 12835
rect 19625 12733 19659 12767
rect 19901 12733 19935 12767
rect 20361 12733 20395 12767
rect 21097 12733 21131 12767
rect 18061 12597 18095 12631
rect 19349 12597 19383 12631
rect 15301 12393 15335 12427
rect 16865 12393 16899 12427
rect 17233 12393 17267 12427
rect 21097 12393 21131 12427
rect 20361 12325 20395 12359
rect 15669 12257 15703 12291
rect 18144 12257 18178 12291
rect 20085 12257 20119 12291
rect 20913 12257 20947 12291
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 17325 12189 17359 12223
rect 17509 12189 17543 12223
rect 17877 12189 17911 12223
rect 19625 12189 19659 12223
rect 19257 12053 19291 12087
rect 15025 11713 15059 11747
rect 17417 11713 17451 11747
rect 15485 11645 15519 11679
rect 17141 11645 17175 11679
rect 18889 11645 18923 11679
rect 20821 11645 20855 11679
rect 15752 11577 15786 11611
rect 18245 11577 18279 11611
rect 19156 11577 19190 11611
rect 16865 11509 16899 11543
rect 18613 11509 18647 11543
rect 20269 11509 20303 11543
rect 21005 11509 21039 11543
rect 13369 11305 13403 11339
rect 16681 11305 16715 11339
rect 18337 11305 18371 11339
rect 18797 11305 18831 11339
rect 19165 11305 19199 11339
rect 19257 11305 19291 11339
rect 19809 11305 19843 11339
rect 20269 11305 20303 11339
rect 21097 11305 21131 11339
rect 17202 11237 17236 11271
rect 12162 11169 12196 11203
rect 13737 11169 13771 11203
rect 14381 11169 14415 11203
rect 15568 11169 15602 11203
rect 20177 11169 20211 11203
rect 20913 11169 20947 11203
rect 12449 11101 12483 11135
rect 13829 11101 13863 11135
rect 13921 11101 13955 11135
rect 15301 11101 15335 11135
rect 16957 11101 16991 11135
rect 19441 11101 19475 11135
rect 20361 11101 20395 11135
rect 13921 10761 13955 10795
rect 15577 10761 15611 10795
rect 15853 10761 15887 10795
rect 16865 10761 16899 10795
rect 16405 10625 16439 10659
rect 17417 10625 17451 10659
rect 12541 10557 12575 10591
rect 14197 10557 14231 10591
rect 14453 10557 14487 10591
rect 18061 10557 18095 10591
rect 19717 10557 19751 10591
rect 19973 10557 20007 10591
rect 12808 10489 12842 10523
rect 16313 10489 16347 10523
rect 18328 10489 18362 10523
rect 16221 10421 16255 10455
rect 17233 10421 17267 10455
rect 17325 10421 17359 10455
rect 19441 10421 19475 10455
rect 21097 10421 21131 10455
rect 13921 10217 13955 10251
rect 18521 10217 18555 10251
rect 18981 10217 19015 10251
rect 19809 10217 19843 10251
rect 20269 10217 20303 10251
rect 15669 10149 15703 10183
rect 17132 10149 17166 10183
rect 13369 10081 13403 10115
rect 13921 10081 13955 10115
rect 14933 10081 14967 10115
rect 15393 10081 15427 10115
rect 16589 10081 16623 10115
rect 18889 10081 18923 10115
rect 20177 10081 20211 10115
rect 20913 10081 20947 10115
rect 13553 10013 13587 10047
rect 16221 10013 16255 10047
rect 16865 10013 16899 10047
rect 19073 10013 19107 10047
rect 20361 10013 20395 10047
rect 16405 9945 16439 9979
rect 18245 9945 18279 9979
rect 14105 9877 14139 9911
rect 14473 9877 14507 9911
rect 16037 9877 16071 9911
rect 16221 9877 16255 9911
rect 21097 9877 21131 9911
rect 11621 9537 11655 9571
rect 13277 9537 13311 9571
rect 16405 9537 16439 9571
rect 17509 9537 17543 9571
rect 19993 9537 20027 9571
rect 13921 9469 13955 9503
rect 17141 9469 17175 9503
rect 18337 9469 18371 9503
rect 18604 9469 18638 9503
rect 11529 9401 11563 9435
rect 14188 9401 14222 9435
rect 20260 9401 20294 9435
rect 11069 9333 11103 9367
rect 11437 9333 11471 9367
rect 13553 9333 13587 9367
rect 15301 9333 15335 9367
rect 15761 9333 15795 9367
rect 16129 9333 16163 9367
rect 16221 9333 16255 9367
rect 16773 9333 16807 9367
rect 19717 9333 19751 9367
rect 21373 9333 21407 9367
rect 8585 9129 8619 9163
rect 11621 9129 11655 9163
rect 13277 9129 13311 9163
rect 14933 9129 14967 9163
rect 16957 9129 16991 9163
rect 18705 9129 18739 9163
rect 19257 9129 19291 9163
rect 19717 9129 19751 9163
rect 21281 9129 21315 9163
rect 12142 9061 12176 9095
rect 13798 9061 13832 9095
rect 8953 8993 8987 9027
rect 9689 8993 9723 9027
rect 10241 8993 10275 9027
rect 10508 8993 10542 9027
rect 11897 8993 11931 9027
rect 15301 8993 15335 9027
rect 15568 8993 15602 9027
rect 18613 8993 18647 9027
rect 19625 8993 19659 9027
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 13553 8925 13587 8959
rect 17969 8925 18003 8959
rect 18889 8925 18923 8959
rect 19809 8925 19843 8959
rect 16681 8789 16715 8823
rect 17417 8789 17451 8823
rect 18245 8789 18279 8823
rect 20269 8789 20303 8823
rect 20913 8789 20947 8823
rect 9505 8585 9539 8619
rect 11161 8585 11195 8619
rect 11989 8585 12023 8619
rect 18061 8585 18095 8619
rect 20821 8585 20855 8619
rect 21281 8585 21315 8619
rect 14841 8517 14875 8551
rect 11437 8449 11471 8483
rect 18981 8449 19015 8483
rect 19441 8449 19475 8483
rect 8125 8381 8159 8415
rect 9781 8381 9815 8415
rect 10037 8381 10071 8415
rect 13093 8381 13127 8415
rect 15853 8381 15887 8415
rect 16120 8381 16154 8415
rect 18245 8381 18279 8415
rect 19708 8381 19742 8415
rect 8392 8313 8426 8347
rect 13553 8313 13587 8347
rect 17509 8313 17543 8347
rect 12817 8245 12851 8279
rect 17233 8245 17267 8279
rect 18613 8245 18647 8279
rect 10057 8041 10091 8075
rect 10517 8041 10551 8075
rect 11529 8041 11563 8075
rect 14013 8041 14047 8075
rect 14381 8041 14415 8075
rect 15301 8041 15335 8075
rect 18613 8041 18647 8075
rect 21281 8041 21315 8075
rect 10333 7973 10367 8007
rect 10885 7973 10919 8007
rect 10241 7905 10275 7939
rect 9321 7837 9355 7871
rect 9689 7701 9723 7735
rect 10333 7701 10367 7735
rect 10425 7905 10459 7939
rect 11897 7905 11931 7939
rect 13369 7905 13403 7939
rect 15669 7905 15703 7939
rect 15761 7905 15795 7939
rect 16856 7905 16890 7939
rect 20177 7905 20211 7939
rect 20913 7905 20947 7939
rect 10977 7837 11011 7871
rect 11069 7837 11103 7871
rect 11989 7837 12023 7871
rect 12173 7837 12207 7871
rect 13461 7837 13495 7871
rect 13553 7837 13587 7871
rect 14473 7837 14507 7871
rect 14657 7837 14691 7871
rect 15853 7837 15887 7871
rect 16589 7837 16623 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 19349 7837 19383 7871
rect 20269 7837 20303 7871
rect 20453 7837 20487 7871
rect 13001 7769 13035 7803
rect 18245 7769 18279 7803
rect 10425 7701 10459 7735
rect 12633 7701 12667 7735
rect 17969 7701 18003 7735
rect 19809 7701 19843 7735
rect 8861 7497 8895 7531
rect 10609 7497 10643 7531
rect 14105 7497 14139 7531
rect 15853 7497 15887 7531
rect 16865 7497 16899 7531
rect 20361 7497 20395 7531
rect 18613 7429 18647 7463
rect 9413 7361 9447 7395
rect 11161 7361 11195 7395
rect 11713 7361 11747 7395
rect 12449 7361 12483 7395
rect 14657 7361 14691 7395
rect 16497 7361 16531 7395
rect 17417 7361 17451 7395
rect 19809 7361 19843 7395
rect 19993 7361 20027 7395
rect 20913 7361 20947 7395
rect 11069 7293 11103 7327
rect 12705 7293 12739 7327
rect 15117 7293 15151 7327
rect 19717 7293 19751 7327
rect 9229 7225 9263 7259
rect 9873 7225 9907 7259
rect 14473 7225 14507 7259
rect 15393 7225 15427 7259
rect 18061 7225 18095 7259
rect 20821 7225 20855 7259
rect 9321 7157 9355 7191
rect 10977 7157 11011 7191
rect 13829 7157 13863 7191
rect 14565 7157 14599 7191
rect 16221 7157 16255 7191
rect 16313 7157 16347 7191
rect 17233 7157 17267 7191
rect 17325 7157 17359 7191
rect 19073 7157 19107 7191
rect 19349 7157 19383 7191
rect 20729 7157 20763 7191
rect 9321 6953 9355 6987
rect 11069 6953 11103 6987
rect 12725 6953 12759 6987
rect 16681 6953 16715 6987
rect 20453 6953 20487 6987
rect 8208 6817 8242 6851
rect 9945 6817 9979 6851
rect 11601 6817 11635 6851
rect 13369 6817 13403 6851
rect 13636 6817 13670 6851
rect 15301 6817 15335 6851
rect 15568 6817 15602 6851
rect 17213 6817 17247 6851
rect 18797 6817 18831 6851
rect 19064 6817 19098 6851
rect 20913 6817 20947 6851
rect 22017 6817 22051 6851
rect 7941 6749 7975 6783
rect 9689 6749 9723 6783
rect 11345 6749 11379 6783
rect 16957 6749 16991 6783
rect 20177 6681 20211 6715
rect 13093 6613 13127 6647
rect 14749 6613 14783 6647
rect 18337 6613 18371 6647
rect 21097 6613 21131 6647
rect 8861 6409 8895 6443
rect 9137 6409 9171 6443
rect 10609 6409 10643 6443
rect 13093 6409 13127 6443
rect 16037 6409 16071 6443
rect 16313 6409 16347 6443
rect 19441 6409 19475 6443
rect 9689 6273 9723 6307
rect 11161 6273 11195 6307
rect 13737 6273 13771 6307
rect 16865 6273 16899 6307
rect 19809 6273 19843 6307
rect 7481 6205 7515 6239
rect 12633 6205 12667 6239
rect 14657 6205 14691 6239
rect 14924 6205 14958 6239
rect 16681 6205 16715 6239
rect 17509 6205 17543 6239
rect 18061 6205 18095 6239
rect 18317 6205 18351 6239
rect 7748 6137 7782 6171
rect 9505 6137 9539 6171
rect 11069 6137 11103 6171
rect 14105 6137 14139 6171
rect 20076 6137 20110 6171
rect 9597 6069 9631 6103
rect 10241 6069 10275 6103
rect 10977 6069 11011 6103
rect 11713 6069 11747 6103
rect 11989 6069 12023 6103
rect 12449 6069 12483 6103
rect 13461 6069 13495 6103
rect 13553 6069 13587 6103
rect 16773 6069 16807 6103
rect 17325 6069 17359 6103
rect 21189 6069 21223 6103
rect 7665 5865 7699 5899
rect 14013 5865 14047 5899
rect 14473 5865 14507 5899
rect 15301 5865 15335 5899
rect 16405 5865 16439 5899
rect 16773 5865 16807 5899
rect 19257 5865 19291 5899
rect 19809 5865 19843 5899
rect 12624 5797 12658 5831
rect 20269 5797 20303 5831
rect 7389 5729 7423 5763
rect 8033 5729 8067 5763
rect 8677 5729 8711 5763
rect 10149 5729 10183 5763
rect 10416 5729 10450 5763
rect 12357 5729 12391 5763
rect 14381 5729 14415 5763
rect 15669 5729 15703 5763
rect 17509 5729 17543 5763
rect 18245 5729 18279 5763
rect 19165 5729 19199 5763
rect 20177 5729 20211 5763
rect 20913 5729 20947 5763
rect 8125 5661 8159 5695
rect 8217 5661 8251 5695
rect 14657 5661 14691 5695
rect 15761 5661 15795 5695
rect 15945 5661 15979 5695
rect 16865 5661 16899 5695
rect 16957 5661 16991 5695
rect 17785 5661 17819 5695
rect 19349 5661 19383 5695
rect 20361 5661 20395 5695
rect 18797 5593 18831 5627
rect 9137 5525 9171 5559
rect 9689 5525 9723 5559
rect 11529 5525 11563 5559
rect 12081 5525 12115 5559
rect 13737 5525 13771 5559
rect 18429 5525 18463 5559
rect 21097 5525 21131 5559
rect 22017 5525 22051 5559
rect 8493 5321 8527 5355
rect 8769 5321 8803 5355
rect 11437 5321 11471 5355
rect 14933 5321 14967 5355
rect 16405 5321 16439 5355
rect 19993 5321 20027 5355
rect 17693 5253 17727 5287
rect 18889 5253 18923 5287
rect 9321 5185 9355 5219
rect 10057 5185 10091 5219
rect 11713 5185 11747 5219
rect 15577 5185 15611 5219
rect 15945 5185 15979 5219
rect 16957 5185 16991 5219
rect 19441 5185 19475 5219
rect 20545 5185 20579 5219
rect 7113 5117 7147 5151
rect 12541 5117 12575 5151
rect 12808 5117 12842 5151
rect 16865 5117 16899 5151
rect 18337 5117 18371 5151
rect 19257 5117 19291 5151
rect 21005 5117 21039 5151
rect 7380 5049 7414 5083
rect 10324 5049 10358 5083
rect 19349 5049 19383 5083
rect 20453 5049 20487 5083
rect 9137 4981 9171 5015
rect 9229 4981 9263 5015
rect 13921 4981 13955 5015
rect 14197 4981 14231 5015
rect 15301 4981 15335 5015
rect 15393 4981 15427 5015
rect 16773 4981 16807 5015
rect 18521 4981 18555 5015
rect 20361 4981 20395 5015
rect 21189 4981 21223 5015
rect 7205 4777 7239 4811
rect 8217 4777 8251 4811
rect 10609 4777 10643 4811
rect 12725 4777 12759 4811
rect 13093 4777 13127 4811
rect 15485 4777 15519 4811
rect 17325 4777 17359 4811
rect 9781 4709 9815 4743
rect 15853 4709 15887 4743
rect 17868 4709 17902 4743
rect 7573 4641 7607 4675
rect 8585 4641 8619 4675
rect 10241 4641 10275 4675
rect 10977 4641 11011 4675
rect 11805 4641 11839 4675
rect 12449 4641 12483 4675
rect 13185 4641 13219 4675
rect 16221 4641 16255 4675
rect 19901 4641 19935 4675
rect 20913 4641 20947 4675
rect 7665 4573 7699 4607
rect 7757 4573 7791 4607
rect 8677 4573 8711 4607
rect 8861 4573 8895 4607
rect 11069 4573 11103 4607
rect 11253 4573 11287 4607
rect 13369 4573 13403 4607
rect 13921 4573 13955 4607
rect 17601 4573 17635 4607
rect 19993 4573 20027 4607
rect 20085 4573 20119 4607
rect 11621 4505 11655 4539
rect 16865 4505 16899 4539
rect 21097 4505 21131 4539
rect 6929 4437 6963 4471
rect 9321 4437 9355 4471
rect 14197 4437 14231 4471
rect 14749 4437 14783 4471
rect 16589 4437 16623 4471
rect 18981 4437 19015 4471
rect 19533 4437 19567 4471
rect 7205 4233 7239 4267
rect 7573 4233 7607 4267
rect 9229 4233 9263 4267
rect 10425 4233 10459 4267
rect 15669 4233 15703 4267
rect 19901 4233 19935 4267
rect 20177 4233 20211 4267
rect 11529 4165 11563 4199
rect 14749 4165 14783 4199
rect 10977 4097 11011 4131
rect 12081 4097 12115 4131
rect 13093 4097 13127 4131
rect 14013 4097 14047 4131
rect 14105 4097 14139 4131
rect 20729 4097 20763 4131
rect 21373 4097 21407 4131
rect 7849 4029 7883 4063
rect 9781 4029 9815 4063
rect 10149 4029 10183 4063
rect 10885 4029 10919 4063
rect 12449 4029 12483 4063
rect 14565 4029 14599 4063
rect 15117 4029 15151 4063
rect 15945 4029 15979 4063
rect 18521 4029 18555 4063
rect 18788 4029 18822 4063
rect 20545 4029 20579 4063
rect 8116 3961 8150 3995
rect 10793 3961 10827 3995
rect 16212 3961 16246 3995
rect 12449 3893 12483 3927
rect 12541 3893 12575 3927
rect 12909 3893 12943 3927
rect 13001 3893 13035 3927
rect 13553 3893 13587 3927
rect 13921 3893 13955 3927
rect 17325 3893 17359 3927
rect 17601 3893 17635 3927
rect 18061 3893 18095 3927
rect 20637 3893 20671 3927
rect 9045 3689 9079 3723
rect 13829 3689 13863 3723
rect 14197 3689 14231 3723
rect 15853 3689 15887 3723
rect 19809 3689 19843 3723
rect 11621 3621 11655 3655
rect 15393 3621 15427 3655
rect 18889 3621 18923 3655
rect 19533 3621 19567 3655
rect 7665 3553 7699 3587
rect 7932 3553 7966 3587
rect 9965 3553 9999 3587
rect 10232 3553 10266 3587
rect 12716 3553 12750 3587
rect 14565 3553 14599 3587
rect 14657 3553 14691 3587
rect 15669 3553 15703 3587
rect 16589 3553 16623 3587
rect 16681 3553 16715 3587
rect 17693 3553 17727 3587
rect 18797 3553 18831 3587
rect 20177 3553 20211 3587
rect 20269 3553 20303 3587
rect 20913 3553 20947 3587
rect 11989 3485 12023 3519
rect 12449 3485 12483 3519
rect 14749 3485 14783 3519
rect 16865 3485 16899 3519
rect 19073 3485 19107 3519
rect 19257 3485 19291 3519
rect 20453 3485 20487 3519
rect 20637 3485 20671 3519
rect 17877 3417 17911 3451
rect 11345 3349 11379 3383
rect 16221 3349 16255 3383
rect 17325 3349 17359 3383
rect 18429 3349 18463 3383
rect 19257 3349 19291 3383
rect 20637 3349 20671 3383
rect 21097 3349 21131 3383
rect 8861 3145 8895 3179
rect 11253 3145 11287 3179
rect 12541 3145 12575 3179
rect 15117 3145 15151 3179
rect 19441 3145 19475 3179
rect 17601 3077 17635 3111
rect 18061 3077 18095 3111
rect 18337 3077 18371 3111
rect 18429 3077 18463 3111
rect 20729 3077 20763 3111
rect 21005 3077 21039 3111
rect 7481 3009 7515 3043
rect 9137 3009 9171 3043
rect 13001 3009 13035 3043
rect 13185 3009 13219 3043
rect 15393 3009 15427 3043
rect 7748 2941 7782 2975
rect 9873 2941 9907 2975
rect 11805 2941 11839 2975
rect 12909 2941 12943 2975
rect 13737 2941 13771 2975
rect 15660 2941 15694 2975
rect 17141 2941 17175 2975
rect 17417 2941 17451 2975
rect 18889 3009 18923 3043
rect 19073 3009 19107 3043
rect 19901 3009 19935 3043
rect 19993 3009 20027 3043
rect 18797 2941 18831 2975
rect 20729 2941 20763 2975
rect 20821 2941 20855 2975
rect 10140 2873 10174 2907
rect 14004 2873 14038 2907
rect 18337 2873 18371 2907
rect 19809 2873 19843 2907
rect 11989 2805 12023 2839
rect 16773 2805 16807 2839
rect 20453 2805 20487 2839
rect 7941 2601 7975 2635
rect 10149 2601 10183 2635
rect 10517 2601 10551 2635
rect 11529 2601 11563 2635
rect 12173 2601 12207 2635
rect 14013 2601 14047 2635
rect 14381 2601 14415 2635
rect 14749 2601 14783 2635
rect 15485 2601 15519 2635
rect 15945 2601 15979 2635
rect 16497 2601 16531 2635
rect 16957 2601 16991 2635
rect 18429 2601 18463 2635
rect 19625 2601 19659 2635
rect 21281 2601 21315 2635
rect 10885 2533 10919 2567
rect 12900 2533 12934 2567
rect 14841 2533 14875 2567
rect 15853 2533 15887 2567
rect 16865 2533 16899 2567
rect 19073 2533 19107 2567
rect 8309 2465 8343 2499
rect 8401 2465 8435 2499
rect 8953 2465 8987 2499
rect 11989 2465 12023 2499
rect 12633 2465 12667 2499
rect 17693 2465 17727 2499
rect 18797 2465 18831 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 8585 2397 8619 2431
rect 9873 2397 9907 2431
rect 10977 2397 11011 2431
rect 11069 2397 11103 2431
rect 15025 2397 15059 2431
rect 16037 2397 16071 2431
rect 17049 2397 17083 2431
rect 9413 2329 9447 2363
rect 20177 2329 20211 2363
rect 20729 2329 20763 2363
rect 7573 2261 7607 2295
rect 17877 2261 17911 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 20438 20040 20444 20052
rect 20399 20012 20444 20040
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 21082 20040 21088 20052
rect 21043 20012 21088 20040
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 20254 19904 20260 19916
rect 20215 19876 20260 19904
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 20990 19496 20996 19508
rect 20951 19468 20996 19496
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 5718 19252 5724 19304
rect 5776 19292 5782 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 5776 19264 6837 19292
rect 5776 19252 5782 19264
rect 6825 19261 6837 19264
rect 6871 19292 6883 19295
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 6871 19264 7389 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7377 19255 7435 19261
rect 18506 19252 18512 19304
rect 18564 19292 18570 19304
rect 19705 19295 19763 19301
rect 19705 19292 19717 19295
rect 18564 19264 19717 19292
rect 18564 19252 18570 19264
rect 19705 19261 19717 19264
rect 19751 19261 19763 19295
rect 19705 19255 19763 19261
rect 20162 19252 20168 19304
rect 20220 19292 20226 19304
rect 20257 19295 20315 19301
rect 20257 19292 20269 19295
rect 20220 19264 20269 19292
rect 20220 19252 20226 19264
rect 20257 19261 20269 19264
rect 20303 19261 20315 19295
rect 20257 19255 20315 19261
rect 20346 19252 20352 19304
rect 20404 19292 20410 19304
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20404 19264 20821 19292
rect 20404 19252 20410 19264
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 7006 19156 7012 19168
rect 6967 19128 7012 19156
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 19889 19159 19947 19165
rect 19889 19156 19901 19159
rect 19300 19128 19901 19156
rect 19300 19116 19306 19128
rect 19889 19125 19901 19128
rect 19935 19125 19947 19159
rect 19889 19119 19947 19125
rect 20441 19159 20499 19165
rect 20441 19125 20453 19159
rect 20487 19156 20499 19159
rect 20530 19156 20536 19168
rect 20487 19128 20536 19156
rect 20487 19125 20499 19128
rect 20441 19119 20499 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 20254 18952 20260 18964
rect 16132 18924 20260 18952
rect 16132 18893 16160 18924
rect 20254 18912 20260 18924
rect 20312 18912 20318 18964
rect 21082 18952 21088 18964
rect 21043 18924 21088 18952
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 12345 18887 12403 18893
rect 12345 18853 12357 18887
rect 12391 18884 12403 18887
rect 16117 18887 16175 18893
rect 12391 18856 15976 18884
rect 12391 18853 12403 18856
rect 12345 18847 12403 18853
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 12069 18819 12127 18825
rect 12069 18816 12081 18819
rect 11756 18788 12081 18816
rect 11756 18776 11762 18788
rect 12069 18785 12081 18788
rect 12115 18785 12127 18819
rect 15838 18816 15844 18828
rect 15799 18788 15844 18816
rect 12069 18779 12127 18785
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 15948 18816 15976 18856
rect 16117 18853 16129 18887
rect 16163 18853 16175 18887
rect 18506 18884 18512 18896
rect 16117 18847 16175 18853
rect 16224 18856 18368 18884
rect 18467 18856 18512 18884
rect 16224 18816 16252 18856
rect 15948 18788 16252 18816
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 18233 18819 18291 18825
rect 18233 18816 18245 18819
rect 16908 18788 18245 18816
rect 16908 18776 16914 18788
rect 18233 18785 18245 18788
rect 18279 18785 18291 18819
rect 18340 18816 18368 18856
rect 18506 18844 18512 18856
rect 18564 18844 18570 18896
rect 20162 18884 20168 18896
rect 18616 18856 20024 18884
rect 20123 18856 20168 18884
rect 18616 18816 18644 18856
rect 19886 18816 19892 18828
rect 18340 18788 18644 18816
rect 19847 18788 19892 18816
rect 18233 18779 18291 18785
rect 19886 18776 19892 18788
rect 19944 18776 19950 18828
rect 19996 18816 20024 18856
rect 20162 18844 20168 18856
rect 20220 18844 20226 18896
rect 20806 18884 20812 18896
rect 20272 18856 20812 18884
rect 20272 18816 20300 18856
rect 20806 18844 20812 18856
rect 20864 18844 20870 18896
rect 19996 18788 20300 18816
rect 20714 18776 20720 18828
rect 20772 18816 20778 18828
rect 20901 18819 20959 18825
rect 20901 18816 20913 18819
rect 20772 18788 20913 18816
rect 20772 18776 20778 18788
rect 20901 18785 20913 18788
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 20990 18408 20996 18420
rect 20951 18380 20996 18408
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 20346 18340 20352 18352
rect 9692 18312 20352 18340
rect 9692 18281 9720 18312
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 8846 18164 8852 18216
rect 8904 18204 8910 18216
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 8904 18176 9413 18204
rect 8904 18164 8910 18176
rect 9401 18173 9413 18176
rect 9447 18173 9459 18207
rect 20806 18204 20812 18216
rect 20767 18176 20812 18204
rect 9401 18167 9459 18173
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 21082 17864 21088 17876
rect 21043 17836 21088 17864
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17728 8355 17731
rect 8386 17728 8392 17740
rect 8343 17700 8392 17728
rect 8343 17697 8355 17700
rect 8297 17691 8355 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 20162 17688 20168 17740
rect 20220 17728 20226 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20220 17700 20913 17728
rect 20220 17688 20226 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 20714 17660 20720 17672
rect 8619 17632 20720 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 18782 17320 18788 17332
rect 18743 17292 18788 17320
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 20990 17320 20996 17332
rect 20951 17292 20996 17320
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 20162 17184 20168 17196
rect 11563 17156 20024 17184
rect 20123 17156 20168 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 11238 17116 11244 17128
rect 11199 17088 11244 17116
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 18012 17088 18613 17116
rect 18012 17076 18018 17088
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 19889 17119 19947 17125
rect 19889 17085 19901 17119
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 13078 17008 13084 17060
rect 13136 17048 13142 17060
rect 19904 17048 19932 17079
rect 13136 17020 19932 17048
rect 19996 17048 20024 17156
rect 20162 17144 20168 17156
rect 20220 17144 20226 17196
rect 20254 17076 20260 17128
rect 20312 17116 20318 17128
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 20312 17088 20821 17116
rect 20312 17076 20318 17088
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 20714 17048 20720 17060
rect 19996 17020 20720 17048
rect 13136 17008 13142 17020
rect 20714 17008 20720 17020
rect 20772 17008 20778 17060
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 21082 16776 21088 16788
rect 21043 16748 21088 16776
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 17954 16708 17960 16720
rect 17915 16680 17960 16708
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 18104 16680 20944 16708
rect 18104 16668 18110 16680
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16640 17739 16643
rect 18782 16640 18788 16652
rect 17727 16612 18788 16640
rect 17727 16609 17739 16612
rect 17681 16603 17739 16609
rect 18782 16600 18788 16612
rect 18840 16600 18846 16652
rect 20916 16649 20944 16680
rect 20901 16643 20959 16649
rect 20901 16609 20913 16643
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16096 20223 16099
rect 20254 16096 20260 16108
rect 20211 16068 20260 16096
rect 20211 16065 20223 16068
rect 20165 16059 20223 16065
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 19794 15988 19800 16040
rect 19852 16028 19858 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19852 16000 19901 16028
rect 19852 15988 19858 16000
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 20806 16028 20812 16040
rect 20767 16000 20812 16028
rect 19889 15991 19947 15997
rect 20806 15988 20812 16000
rect 20864 15988 20870 16040
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 21082 15688 21088 15700
rect 21043 15660 21088 15688
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 14645 15623 14703 15629
rect 14645 15589 14657 15623
rect 14691 15620 14703 15623
rect 18046 15620 18052 15632
rect 14691 15592 18052 15620
rect 14691 15589 14703 15592
rect 14645 15583 14703 15589
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 13998 15512 14004 15564
rect 14056 15552 14062 15564
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 14056 15524 14381 15552
rect 14056 15512 14062 15524
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 15252 15524 20269 15552
rect 15252 15512 15258 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20772 15524 20913 15552
rect 20772 15512 20778 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 20990 15144 20996 15156
rect 20951 15116 20996 15144
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 15194 15008 15200 15020
rect 11931 14980 15200 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 11609 14943 11667 14949
rect 11609 14940 11621 14943
rect 11112 14912 11621 14940
rect 11112 14900 11118 14912
rect 11609 14909 11621 14912
rect 11655 14909 11667 14943
rect 11609 14903 11667 14909
rect 18690 14900 18696 14952
rect 18748 14940 18754 14952
rect 20809 14943 20867 14949
rect 20809 14940 20821 14943
rect 18748 14912 20821 14940
rect 18748 14900 18754 14912
rect 20809 14909 20821 14912
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 20533 14603 20591 14609
rect 20533 14569 20545 14603
rect 20579 14600 20591 14603
rect 20622 14600 20628 14612
rect 20579 14572 20628 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 9953 14535 10011 14541
rect 9953 14501 9965 14535
rect 9999 14532 10011 14535
rect 20806 14532 20812 14544
rect 9999 14504 20812 14532
rect 9999 14501 10011 14504
rect 9953 14495 10011 14501
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 8570 14424 8576 14476
rect 8628 14464 8634 14476
rect 8757 14467 8815 14473
rect 8757 14464 8769 14467
rect 8628 14436 8769 14464
rect 8628 14424 8634 14436
rect 8757 14433 8769 14436
rect 8803 14433 8815 14467
rect 9674 14464 9680 14476
rect 9635 14436 9680 14464
rect 8757 14427 8815 14433
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 18782 14424 18788 14476
rect 18840 14464 18846 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 18840 14436 20913 14464
rect 18840 14424 18846 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 9033 14399 9091 14405
rect 9033 14365 9045 14399
rect 9079 14396 9091 14399
rect 20714 14396 20720 14408
rect 9079 14368 20720 14396
rect 9079 14365 9091 14368
rect 9033 14359 9091 14365
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 20714 13920 20720 13932
rect 20675 13892 20720 13920
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 11020 13824 11161 13852
rect 11020 13812 11026 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11149 13815 11207 13821
rect 11425 13855 11483 13861
rect 11425 13821 11437 13855
rect 11471 13852 11483 13855
rect 18690 13852 18696 13864
rect 11471 13824 18696 13852
rect 11471 13821 11483 13824
rect 11425 13815 11483 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20622 13852 20628 13864
rect 20395 13824 20628 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 17862 13512 17868 13524
rect 16163 13484 17868 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 20438 13512 20444 13524
rect 20399 13484 20444 13512
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 21082 13512 21088 13524
rect 21043 13484 21088 13512
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 16476 13447 16534 13453
rect 16476 13413 16488 13447
rect 16522 13444 16534 13447
rect 16574 13444 16580 13456
rect 16522 13416 16580 13444
rect 16522 13413 16534 13416
rect 16476 13407 16534 13413
rect 16574 13404 16580 13416
rect 16632 13444 16638 13456
rect 17957 13447 18015 13453
rect 17957 13444 17969 13447
rect 16632 13416 17969 13444
rect 16632 13404 16638 13416
rect 17957 13413 17969 13416
rect 18003 13413 18015 13447
rect 17957 13407 18015 13413
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13044 13348 13553 13376
rect 13044 13336 13050 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13376 13875 13379
rect 18782 13376 18788 13388
rect 13863 13348 18788 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13376 20315 13379
rect 20530 13376 20536 13388
rect 20303 13348 20536 13376
rect 20303 13345 20315 13348
rect 20257 13339 20315 13345
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 20901 13379 20959 13385
rect 20901 13345 20913 13379
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 16163 13280 16221 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 19978 13268 19984 13320
rect 20036 13308 20042 13320
rect 20916 13308 20944 13339
rect 20036 13280 20944 13308
rect 20036 13268 20042 13280
rect 16482 13132 16488 13184
rect 16540 13172 16546 13184
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 16540 13144 17601 13172
rect 16540 13132 16546 13144
rect 17589 13141 17601 13144
rect 17635 13141 17647 13175
rect 17589 13135 17647 13141
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13172 20039 13175
rect 20254 13172 20260 13184
rect 20027 13144 20260 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 20530 12832 20536 12844
rect 14332 12804 20392 12832
rect 20491 12804 20536 12832
rect 14332 12792 14338 12804
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19576 12736 19625 12764
rect 19576 12724 19582 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 19978 12764 19984 12776
rect 19935 12736 19984 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 20364 12773 20392 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 21085 12767 21143 12773
rect 21085 12764 21097 12767
rect 20496 12736 21097 12764
rect 20496 12724 20502 12736
rect 21085 12733 21097 12736
rect 21131 12733 21143 12767
rect 21085 12727 21143 12733
rect 18046 12628 18052 12640
rect 18007 12600 18052 12628
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 20622 12628 20628 12640
rect 19383 12600 20628 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15838 12424 15844 12436
rect 15335 12396 15844 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 16850 12424 16856 12436
rect 16811 12396 16856 12424
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 18046 12424 18052 12436
rect 17267 12396 18052 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 21082 12424 21088 12436
rect 21043 12396 21088 12424
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 13170 12316 13176 12368
rect 13228 12356 13234 12368
rect 20162 12356 20168 12368
rect 13228 12328 20168 12356
rect 13228 12316 13234 12328
rect 20162 12316 20168 12328
rect 20220 12316 20226 12368
rect 20349 12359 20407 12365
rect 20349 12325 20361 12359
rect 20395 12356 20407 12359
rect 20438 12356 20444 12368
rect 20395 12328 20444 12356
rect 20395 12325 20407 12328
rect 20349 12319 20407 12325
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 18138 12297 18144 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15068 12260 15669 12288
rect 15068 12248 15074 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 18132 12288 18144 12297
rect 15657 12251 15715 12257
rect 17512 12260 18144 12288
rect 15746 12220 15752 12232
rect 15707 12192 15752 12220
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15930 12220 15936 12232
rect 15891 12192 15936 12220
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17512 12229 17540 12260
rect 18132 12251 18144 12260
rect 18138 12248 18144 12251
rect 18196 12248 18202 12300
rect 20070 12288 20076 12300
rect 20031 12260 20076 12288
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12189 17555 12223
rect 17862 12220 17868 12232
rect 17823 12192 17868 12220
rect 17497 12183 17555 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19208 12192 19625 12220
rect 19208 12180 19214 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 19886 12152 19892 12164
rect 18800 12124 19892 12152
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 18800 12084 18828 12124
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 19242 12084 19248 12096
rect 13412 12056 18828 12084
rect 19203 12056 19248 12084
rect 13412 12044 13418 12056
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 12250 11840 12256 11892
rect 12308 11880 12314 11892
rect 17402 11880 17408 11892
rect 12308 11852 17408 11880
rect 12308 11840 12314 11852
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 20898 11880 20904 11892
rect 18892 11852 20904 11880
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 11790 11744 11796 11756
rect 11020 11716 11796 11744
rect 11020 11704 11026 11716
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 15010 11744 15016 11756
rect 14971 11716 15016 11744
rect 15010 11704 15016 11716
rect 15068 11704 15074 11756
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11744 17463 11747
rect 18892 11744 18920 11852
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 17451 11716 18920 11744
rect 17451 11713 17463 11716
rect 17405 11707 17463 11713
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 15344 11648 15485 11676
rect 15344 11636 15350 11648
rect 15473 11645 15485 11648
rect 15519 11645 15531 11679
rect 15473 11639 15531 11645
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 16816 11648 17141 11676
rect 16816 11636 16822 11648
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 17920 11648 18889 11676
rect 17920 11636 17926 11648
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 19076 11648 20484 11676
rect 15740 11611 15798 11617
rect 15740 11577 15752 11611
rect 15786 11608 15798 11611
rect 15930 11608 15936 11620
rect 15786 11580 15936 11608
rect 15786 11577 15798 11580
rect 15740 11571 15798 11577
rect 15930 11568 15936 11580
rect 15988 11608 15994 11620
rect 16666 11608 16672 11620
rect 15988 11580 16672 11608
rect 15988 11568 15994 11580
rect 16666 11568 16672 11580
rect 16724 11568 16730 11620
rect 18233 11611 18291 11617
rect 18233 11577 18245 11611
rect 18279 11608 18291 11611
rect 19076 11608 19104 11648
rect 18279 11580 19104 11608
rect 19144 11611 19202 11617
rect 18279 11577 18291 11580
rect 18233 11571 18291 11577
rect 19144 11577 19156 11611
rect 19190 11608 19202 11611
rect 19242 11608 19248 11620
rect 19190 11580 19248 11608
rect 19190 11577 19202 11580
rect 19144 11571 19202 11577
rect 19242 11568 19248 11580
rect 19300 11608 19306 11620
rect 20346 11608 20352 11620
rect 19300 11580 20352 11608
rect 19300 11568 19306 11580
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 20456 11608 20484 11648
rect 20622 11636 20628 11688
rect 20680 11676 20686 11688
rect 20809 11679 20867 11685
rect 20809 11676 20821 11679
rect 20680 11648 20821 11676
rect 20680 11636 20686 11648
rect 20809 11645 20821 11648
rect 20855 11645 20867 11679
rect 20809 11639 20867 11645
rect 20898 11608 20904 11620
rect 20456 11580 20904 11608
rect 20898 11568 20904 11580
rect 20956 11568 20962 11620
rect 16850 11540 16856 11552
rect 16811 11512 16856 11540
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 19334 11540 19340 11552
rect 18647 11512 19340 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 20257 11543 20315 11549
rect 20257 11540 20269 11543
rect 19484 11512 20269 11540
rect 19484 11500 19490 11512
rect 20257 11509 20269 11512
rect 20303 11509 20315 11543
rect 20257 11503 20315 11509
rect 20993 11543 21051 11549
rect 20993 11509 21005 11543
rect 21039 11540 21051 11543
rect 22094 11540 22100 11552
rect 21039 11512 22100 11540
rect 21039 11509 21051 11512
rect 20993 11503 21051 11509
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 13170 11336 13176 11348
rect 4120 11308 13176 11336
rect 4120 11296 4126 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13354 11336 13360 11348
rect 13315 11308 13360 11336
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 16666 11336 16672 11348
rect 16627 11308 16672 11336
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 18196 11308 18337 11336
rect 18196 11296 18202 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18782 11336 18788 11348
rect 18743 11308 18788 11336
rect 18325 11299 18383 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 19150 11336 19156 11348
rect 19111 11308 19156 11336
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 19245 11339 19303 11345
rect 19245 11305 19257 11339
rect 19291 11336 19303 11339
rect 19797 11339 19855 11345
rect 19797 11336 19809 11339
rect 19291 11308 19809 11336
rect 19291 11305 19303 11308
rect 19245 11299 19303 11305
rect 19797 11305 19809 11308
rect 19843 11305 19855 11339
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 19797 11299 19855 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11305 21143 11339
rect 21085 11299 21143 11305
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 17190 11271 17248 11277
rect 17190 11268 17202 11271
rect 16908 11240 17202 11268
rect 16908 11228 16914 11240
rect 17190 11237 17202 11240
rect 17236 11237 17248 11271
rect 17190 11231 17248 11237
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 21100 11268 21128 11299
rect 17460 11240 21128 11268
rect 17460 11228 17466 11240
rect 12158 11209 12164 11212
rect 12150 11203 12164 11209
rect 12150 11200 12162 11203
rect 12119 11172 12162 11200
rect 12150 11169 12162 11172
rect 12150 11163 12164 11169
rect 12158 11160 12164 11163
rect 12216 11160 12222 11212
rect 15562 11209 15568 11212
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11200 13783 11203
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 13771 11172 14381 11200
rect 13771 11169 13783 11172
rect 13725 11163 13783 11169
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 15556 11163 15568 11209
rect 15620 11200 15626 11212
rect 15620 11172 15656 11200
rect 15562 11160 15568 11163
rect 15620 11160 15626 11172
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19886 11200 19892 11212
rect 19392 11172 19892 11200
rect 19392 11160 19398 11172
rect 19886 11160 19892 11172
rect 19944 11200 19950 11212
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 19944 11172 20177 11200
rect 19944 11160 19950 11172
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20898 11200 20904 11212
rect 20859 11172 20904 11200
rect 20165 11163 20223 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 12618 11132 12624 11144
rect 12483 11104 12624 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13814 11132 13820 11144
rect 13775 11104 13820 11132
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 15286 11132 15292 11144
rect 13964 11104 14009 11132
rect 15199 11104 15292 11132
rect 13964 11092 13970 11104
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 16942 11132 16948 11144
rect 16903 11104 16948 11132
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 19426 11132 19432 11144
rect 19387 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20404 11104 20449 11132
rect 20404 11092 20410 11104
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 15304 10996 15332 11092
rect 14240 10968 15332 10996
rect 14240 10956 14246 10968
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 13906 10792 13912 10804
rect 13867 10764 13912 10792
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 15562 10792 15568 10804
rect 15523 10764 15568 10792
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 15746 10752 15752 10804
rect 15804 10792 15810 10804
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15804 10764 15853 10792
rect 15804 10752 15810 10764
rect 15841 10761 15853 10764
rect 15887 10761 15899 10795
rect 15841 10755 15899 10761
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 17310 10792 17316 10804
rect 16899 10764 17316 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 13924 10656 13952 10752
rect 15580 10656 15608 10752
rect 16393 10659 16451 10665
rect 16393 10656 16405 10659
rect 13924 10628 14320 10656
rect 15580 10628 16405 10656
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12492 10560 12541 10588
rect 12492 10548 12498 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 14182 10588 14188 10600
rect 14143 10560 14188 10588
rect 12529 10551 12587 10557
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 14292 10588 14320 10628
rect 16393 10625 16405 10628
rect 16439 10625 16451 10659
rect 16393 10619 16451 10625
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 16908 10628 17417 10656
rect 16908 10616 16914 10628
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19484 10628 19840 10656
rect 19484 10616 19490 10628
rect 14441 10591 14499 10597
rect 14441 10588 14453 10591
rect 14292 10560 14453 10588
rect 14441 10557 14453 10560
rect 14487 10557 14499 10591
rect 14441 10551 14499 10557
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17862 10588 17868 10600
rect 17000 10560 17868 10588
rect 17000 10548 17006 10560
rect 17862 10548 17868 10560
rect 17920 10588 17926 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17920 10560 18061 10588
rect 17920 10548 17926 10560
rect 18049 10557 18061 10560
rect 18095 10588 18107 10591
rect 19705 10591 19763 10597
rect 19705 10588 19717 10591
rect 18095 10560 19717 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 19705 10557 19717 10560
rect 19751 10557 19763 10591
rect 19812 10588 19840 10628
rect 19961 10591 20019 10597
rect 19961 10588 19973 10591
rect 19812 10560 19973 10588
rect 19705 10551 19763 10557
rect 19961 10557 19973 10560
rect 20007 10557 20019 10591
rect 19961 10551 20019 10557
rect 12796 10523 12854 10529
rect 12796 10489 12808 10523
rect 12842 10520 12854 10523
rect 13906 10520 13912 10532
rect 12842 10492 13912 10520
rect 12842 10489 12854 10492
rect 12796 10483 12854 10489
rect 13906 10480 13912 10492
rect 13964 10480 13970 10532
rect 15746 10480 15752 10532
rect 15804 10520 15810 10532
rect 18322 10529 18328 10532
rect 16301 10523 16359 10529
rect 16301 10520 16313 10523
rect 15804 10492 16313 10520
rect 15804 10480 15810 10492
rect 16301 10489 16313 10492
rect 16347 10489 16359 10523
rect 18316 10520 18328 10529
rect 18283 10492 18328 10520
rect 16301 10483 16359 10489
rect 18316 10483 18328 10492
rect 18322 10480 18328 10483
rect 18380 10480 18386 10532
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 17218 10452 17224 10464
rect 17179 10424 17224 10452
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 17313 10455 17371 10461
rect 17313 10421 17325 10455
rect 17359 10452 17371 10455
rect 18046 10452 18052 10464
rect 17359 10424 18052 10452
rect 17359 10421 17371 10424
rect 17313 10415 17371 10421
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 19426 10452 19432 10464
rect 19387 10424 19432 10452
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 21082 10452 21088 10464
rect 21043 10424 21088 10452
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 13909 10251 13967 10257
rect 13909 10217 13921 10251
rect 13955 10248 13967 10251
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 13955 10220 18521 10248
rect 13955 10217 13967 10220
rect 13909 10211 13967 10217
rect 18509 10217 18521 10220
rect 18555 10217 18567 10251
rect 18509 10211 18567 10217
rect 18969 10251 19027 10257
rect 18969 10217 18981 10251
rect 19015 10248 19027 10251
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19015 10220 19809 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 20254 10248 20260 10260
rect 20215 10220 20260 10248
rect 19797 10211 19855 10217
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 15657 10183 15715 10189
rect 15657 10180 15669 10183
rect 9640 10152 15669 10180
rect 9640 10140 9646 10152
rect 15657 10149 15669 10152
rect 15703 10180 15715 10183
rect 16206 10180 16212 10192
rect 15703 10152 16212 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 17120 10183 17178 10189
rect 16408 10152 17080 10180
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10112 13415 10115
rect 13909 10115 13967 10121
rect 13909 10112 13921 10115
rect 13403 10084 13921 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 13909 10081 13921 10084
rect 13955 10081 13967 10115
rect 13909 10075 13967 10081
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10112 14979 10115
rect 15381 10115 15439 10121
rect 15381 10112 15393 10115
rect 14967 10084 15393 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15381 10081 15393 10084
rect 15427 10112 15439 10115
rect 16408 10112 16436 10152
rect 16574 10112 16580 10124
rect 15427 10084 16436 10112
rect 16535 10084 16580 10112
rect 15427 10081 15439 10084
rect 15381 10075 15439 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 16942 10112 16948 10124
rect 16868 10084 16948 10112
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 16868 10053 16896 10084
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 17052 10112 17080 10152
rect 17120 10149 17132 10183
rect 17166 10180 17178 10183
rect 21082 10180 21088 10192
rect 17166 10152 21088 10180
rect 17166 10149 17178 10152
rect 17120 10143 17178 10149
rect 18046 10112 18052 10124
rect 17052 10084 18052 10112
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 18196 10084 18889 10112
rect 18196 10072 18202 10084
rect 18877 10081 18889 10084
rect 18923 10081 18935 10115
rect 18877 10075 18935 10081
rect 19886 10072 19892 10124
rect 19944 10112 19950 10124
rect 20165 10115 20223 10121
rect 20165 10112 20177 10115
rect 19944 10084 20177 10112
rect 19944 10072 19950 10084
rect 20165 10081 20177 10084
rect 20211 10081 20223 10115
rect 20272 10112 20300 10152
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 20898 10112 20904 10124
rect 20272 10084 20392 10112
rect 20859 10084 20904 10112
rect 20165 10075 20223 10081
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 12216 10016 13553 10044
rect 12216 10004 12222 10016
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 13541 10007 13599 10013
rect 13648 10016 16221 10044
rect 13354 9936 13360 9988
rect 13412 9976 13418 9988
rect 13648 9976 13676 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10013 16911 10047
rect 18322 10044 18328 10056
rect 18235 10016 18328 10044
rect 16853 10007 16911 10013
rect 13412 9948 13676 9976
rect 13412 9936 13418 9948
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 16393 9979 16451 9985
rect 16393 9976 16405 9979
rect 14240 9948 16405 9976
rect 14240 9936 14246 9948
rect 16393 9945 16405 9948
rect 16439 9976 16451 9979
rect 16868 9976 16896 10007
rect 18248 9985 18276 10016
rect 18322 10004 18328 10016
rect 18380 10044 18386 10056
rect 20364 10053 20392 10084
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 19061 10047 19119 10053
rect 19061 10044 19073 10047
rect 18380 10016 19073 10044
rect 18380 10004 18386 10016
rect 19061 10013 19073 10016
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 20349 10047 20407 10053
rect 20349 10013 20361 10047
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 16439 9948 16896 9976
rect 18233 9979 18291 9985
rect 16439 9945 16451 9948
rect 16393 9939 16451 9945
rect 18233 9945 18245 9979
rect 18279 9945 18291 9979
rect 18233 9939 18291 9945
rect 658 9868 664 9920
rect 716 9908 722 9920
rect 9582 9908 9588 9920
rect 716 9880 9588 9908
rect 716 9868 722 9880
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 14090 9908 14096 9920
rect 14051 9880 14096 9908
rect 14090 9868 14096 9880
rect 14148 9908 14154 9920
rect 14461 9911 14519 9917
rect 14461 9908 14473 9911
rect 14148 9880 14473 9908
rect 14148 9868 14154 9880
rect 14461 9877 14473 9880
rect 14507 9877 14519 9911
rect 14461 9871 14519 9877
rect 15746 9868 15752 9920
rect 15804 9908 15810 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15804 9880 16037 9908
rect 15804 9868 15810 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 16025 9871 16083 9877
rect 16209 9911 16267 9917
rect 16209 9877 16221 9911
rect 16255 9908 16267 9911
rect 21085 9911 21143 9917
rect 21085 9908 21097 9911
rect 16255 9880 21097 9908
rect 16255 9877 16267 9880
rect 16209 9871 16267 9877
rect 21085 9877 21097 9880
rect 21131 9877 21143 9911
rect 21085 9871 21143 9877
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 14182 9704 14188 9716
rect 13924 9676 14188 9704
rect 11606 9568 11612 9580
rect 11567 9540 11612 9568
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 13262 9568 13268 9580
rect 13223 9540 13268 9568
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 13924 9509 13952 9676
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 18340 9676 19380 9704
rect 17862 9596 17868 9648
rect 17920 9636 17926 9648
rect 18340 9636 18368 9676
rect 17920 9608 18368 9636
rect 17920 9596 17926 9608
rect 16393 9571 16451 9577
rect 16393 9537 16405 9571
rect 16439 9568 16451 9571
rect 16666 9568 16672 9580
rect 16439 9540 16672 9568
rect 16439 9537 16451 9540
rect 16393 9531 16451 9537
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 18138 9568 18144 9580
rect 17543 9540 18144 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13688 9472 13921 9500
rect 13688 9460 13694 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 15746 9460 15752 9512
rect 15804 9500 15810 9512
rect 18340 9509 18368 9608
rect 19352 9568 19380 9676
rect 19981 9571 20039 9577
rect 19981 9568 19993 9571
rect 19352 9540 19993 9568
rect 19981 9537 19993 9540
rect 20027 9537 20039 9571
rect 19981 9531 20039 9537
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 15804 9472 17141 9500
rect 15804 9460 15810 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 18325 9503 18383 9509
rect 18325 9469 18337 9503
rect 18371 9500 18383 9503
rect 18414 9500 18420 9512
rect 18371 9472 18420 9500
rect 18371 9469 18383 9472
rect 18325 9463 18383 9469
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 18592 9503 18650 9509
rect 18592 9469 18604 9503
rect 18638 9500 18650 9503
rect 19426 9500 19432 9512
rect 18638 9472 19432 9500
rect 18638 9469 18650 9472
rect 18592 9463 18650 9469
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 10502 9392 10508 9444
rect 10560 9432 10566 9444
rect 11517 9435 11575 9441
rect 11517 9432 11529 9435
rect 10560 9404 11529 9432
rect 10560 9392 10566 9404
rect 11517 9401 11529 9404
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 14176 9435 14234 9441
rect 14176 9401 14188 9435
rect 14222 9432 14234 9435
rect 14734 9432 14740 9444
rect 14222 9404 14740 9432
rect 14222 9401 14234 9404
rect 14176 9395 14234 9401
rect 14734 9392 14740 9404
rect 14792 9392 14798 9444
rect 19794 9432 19800 9444
rect 15764 9404 19800 9432
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 11020 9336 11069 9364
rect 11020 9324 11026 9336
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 11057 9327 11115 9333
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11425 9367 11483 9373
rect 11425 9364 11437 9367
rect 11296 9336 11437 9364
rect 11296 9324 11302 9336
rect 11425 9333 11437 9336
rect 11471 9333 11483 9367
rect 11425 9327 11483 9333
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13320 9336 13553 9364
rect 13320 9324 13326 9336
rect 13541 9333 13553 9336
rect 13587 9333 13599 9367
rect 13541 9327 13599 9333
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15378 9364 15384 9376
rect 15335 9336 15384 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15764 9373 15792 9404
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 20248 9435 20306 9441
rect 20248 9401 20260 9435
rect 20294 9432 20306 9435
rect 20622 9432 20628 9444
rect 20294 9404 20628 9432
rect 20294 9401 20306 9404
rect 20248 9395 20306 9401
rect 20622 9392 20628 9404
rect 20680 9392 20686 9444
rect 15749 9367 15807 9373
rect 15749 9333 15761 9367
rect 15795 9333 15807 9367
rect 16114 9364 16120 9376
rect 16075 9336 16120 9364
rect 15749 9327 15807 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16206 9324 16212 9376
rect 16264 9364 16270 9376
rect 16264 9336 16309 9364
rect 16264 9324 16270 9336
rect 16390 9324 16396 9376
rect 16448 9364 16454 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 16448 9336 16773 9364
rect 16448 9324 16454 9336
rect 16761 9333 16773 9336
rect 16807 9364 16819 9367
rect 17218 9364 17224 9376
rect 16807 9336 17224 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 19702 9364 19708 9376
rect 19663 9336 19708 9364
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 20162 9364 20168 9376
rect 20036 9336 20168 9364
rect 20036 9324 20042 9336
rect 20162 9324 20168 9336
rect 20220 9364 20226 9376
rect 21361 9367 21419 9373
rect 21361 9364 21373 9367
rect 20220 9336 21373 9364
rect 20220 9324 20226 9336
rect 21361 9333 21373 9336
rect 21407 9333 21419 9367
rect 21361 9327 21419 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 9674 9160 9680 9172
rect 8619 9132 9680 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 11606 9160 11612 9172
rect 11567 9132 11612 9160
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 13265 9163 13323 9169
rect 13265 9129 13277 9163
rect 13311 9129 13323 9163
rect 13265 9123 13323 9129
rect 11624 9092 11652 9120
rect 12130 9095 12188 9101
rect 12130 9092 12142 9095
rect 10244 9064 11100 9092
rect 11624 9064 12142 9092
rect 8941 9027 8999 9033
rect 8941 8993 8953 9027
rect 8987 9024 8999 9027
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 8987 8996 9689 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10244 9033 10272 9064
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 10100 8996 10241 9024
rect 10100 8984 10106 8996
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 10496 9027 10554 9033
rect 10496 8993 10508 9027
rect 10542 9024 10554 9027
rect 10962 9024 10968 9036
rect 10542 8996 10968 9024
rect 10542 8993 10554 8996
rect 10496 8987 10554 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11072 9024 11100 9064
rect 12130 9061 12142 9064
rect 12176 9061 12188 9095
rect 13280 9092 13308 9123
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 14921 9163 14979 9169
rect 14921 9160 14933 9163
rect 14792 9132 14933 9160
rect 14792 9120 14798 9132
rect 14921 9129 14933 9132
rect 14967 9129 14979 9163
rect 14921 9123 14979 9129
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16172 9132 16957 9160
rect 16172 9120 16178 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 18693 9163 18751 9169
rect 18693 9129 18705 9163
rect 18739 9160 18751 9163
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 18739 9132 19257 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 19705 9163 19763 9169
rect 19705 9129 19717 9163
rect 19751 9160 19763 9163
rect 20530 9160 20536 9172
rect 19751 9132 20536 9160
rect 19751 9129 19763 9132
rect 19705 9123 19763 9129
rect 20530 9120 20536 9132
rect 20588 9160 20594 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 20588 9132 21281 9160
rect 20588 9120 20594 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 13538 9092 13544 9104
rect 13280 9064 13544 9092
rect 12130 9055 12188 9061
rect 13538 9052 13544 9064
rect 13596 9092 13602 9104
rect 13786 9095 13844 9101
rect 13786 9092 13798 9095
rect 13596 9064 13798 9092
rect 13596 9052 13602 9064
rect 13786 9061 13798 9064
rect 13832 9061 13844 9095
rect 13786 9055 13844 9061
rect 19426 9052 19432 9104
rect 19484 9092 19490 9104
rect 19484 9064 20024 9092
rect 19484 9052 19490 9064
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 11072 8996 11897 9024
rect 11885 8993 11897 8996
rect 11931 9024 11943 9027
rect 12434 9024 12440 9036
rect 11931 8996 12440 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 12434 8984 12440 8996
rect 12492 8984 12498 9036
rect 13630 9024 13636 9036
rect 13543 8996 13636 9024
rect 9030 8956 9036 8968
rect 8991 8928 9036 8956
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9490 8956 9496 8968
rect 9263 8928 9496 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 13556 8965 13584 8996
rect 13630 8984 13636 8996
rect 13688 9024 13694 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 13688 8996 15301 9024
rect 13688 8984 13694 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15378 8984 15384 9036
rect 15436 9024 15442 9036
rect 15556 9027 15614 9033
rect 15556 9024 15568 9027
rect 15436 8996 15568 9024
rect 15436 8984 15442 8996
rect 15556 8993 15568 8996
rect 15602 9024 15614 9027
rect 15838 9024 15844 9036
rect 15602 8996 15844 9024
rect 15602 8993 15614 8996
rect 15556 8987 15614 8993
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 16114 8984 16120 9036
rect 16172 9024 16178 9036
rect 16850 9024 16856 9036
rect 16172 8996 16856 9024
rect 16172 8984 16178 8996
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 18966 9024 18972 9036
rect 18647 8996 18972 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 18966 8984 18972 8996
rect 19024 8984 19030 9036
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 9024 19671 9027
rect 19886 9024 19892 9036
rect 19659 8996 19892 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18782 8956 18788 8968
rect 18003 8928 18788 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8956 18935 8959
rect 19702 8956 19708 8968
rect 18923 8928 19708 8956
rect 18923 8925 18935 8928
rect 18877 8919 18935 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8956 19855 8959
rect 19996 8956 20024 9064
rect 19843 8928 20024 8956
rect 19843 8925 19855 8928
rect 19797 8919 19855 8925
rect 20714 8888 20720 8900
rect 16224 8860 18368 8888
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 11790 8820 11796 8832
rect 10468 8792 11796 8820
rect 10468 8780 10474 8792
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 14182 8780 14188 8832
rect 14240 8820 14246 8832
rect 16224 8820 16252 8860
rect 16666 8820 16672 8832
rect 14240 8792 16252 8820
rect 16627 8792 16672 8820
rect 14240 8780 14246 8792
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 16908 8792 17417 8820
rect 16908 8780 16914 8792
rect 17405 8789 17417 8792
rect 17451 8789 17463 8823
rect 17405 8783 17463 8789
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 18233 8823 18291 8829
rect 18233 8820 18245 8823
rect 18012 8792 18245 8820
rect 18012 8780 18018 8792
rect 18233 8789 18245 8792
rect 18279 8789 18291 8823
rect 18340 8820 18368 8860
rect 19812 8860 20720 8888
rect 19812 8820 19840 8860
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 18340 8792 19840 8820
rect 18233 8783 18291 8789
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 20257 8823 20315 8829
rect 20257 8820 20269 8823
rect 19944 8792 20269 8820
rect 19944 8780 19950 8792
rect 20257 8789 20269 8792
rect 20303 8820 20315 8823
rect 20901 8823 20959 8829
rect 20901 8820 20913 8823
rect 20303 8792 20913 8820
rect 20303 8789 20315 8792
rect 20257 8783 20315 8789
rect 20901 8789 20913 8792
rect 20947 8789 20959 8823
rect 20901 8783 20959 8789
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 11020 8588 11161 8616
rect 11020 8576 11026 8588
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 11149 8579 11207 8585
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 11977 8619 12035 8625
rect 11977 8616 11989 8619
rect 11848 8588 11989 8616
rect 11848 8576 11854 8588
rect 11977 8585 11989 8588
rect 12023 8616 12035 8619
rect 16114 8616 16120 8628
rect 12023 8588 16120 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 17494 8616 17500 8628
rect 16632 8588 17500 8616
rect 16632 8576 16638 8588
rect 17494 8576 17500 8588
rect 17552 8616 17558 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17552 8588 18061 8616
rect 17552 8576 17558 8588
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 18049 8579 18107 8585
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 20809 8619 20867 8625
rect 20809 8616 20821 8619
rect 20680 8588 20821 8616
rect 20680 8576 20686 8588
rect 20809 8585 20821 8588
rect 20855 8585 20867 8619
rect 20809 8579 20867 8585
rect 20898 8576 20904 8628
rect 20956 8616 20962 8628
rect 21269 8619 21327 8625
rect 21269 8616 21281 8619
rect 20956 8588 21281 8616
rect 20956 8576 20962 8588
rect 21269 8585 21281 8588
rect 21315 8585 21327 8619
rect 21269 8579 21327 8585
rect 9508 8480 9536 8576
rect 13630 8508 13636 8560
rect 13688 8548 13694 8560
rect 14829 8551 14887 8557
rect 14829 8548 14841 8551
rect 13688 8520 14841 8548
rect 13688 8508 13694 8520
rect 14829 8517 14841 8520
rect 14875 8517 14887 8551
rect 14829 8511 14887 8517
rect 9508 8452 9904 8480
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8412 8171 8415
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 8159 8384 9781 8412
rect 8159 8381 8171 8384
rect 8113 8375 8171 8381
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 9876 8412 9904 8452
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11425 8483 11483 8489
rect 11425 8480 11437 8483
rect 11296 8452 11437 8480
rect 11296 8440 11302 8452
rect 11425 8449 11437 8452
rect 11471 8449 11483 8483
rect 11425 8443 11483 8449
rect 10025 8415 10083 8421
rect 10025 8412 10037 8415
rect 9876 8384 10037 8412
rect 9769 8375 9827 8381
rect 10025 8381 10037 8384
rect 10071 8381 10083 8415
rect 10025 8375 10083 8381
rect 13081 8415 13139 8421
rect 13081 8381 13093 8415
rect 13127 8412 13139 8415
rect 14366 8412 14372 8424
rect 13127 8384 14372 8412
rect 13127 8381 13139 8384
rect 13081 8375 13139 8381
rect 8380 8347 8438 8353
rect 8380 8313 8392 8347
rect 8426 8344 8438 8347
rect 9214 8344 9220 8356
rect 8426 8316 9220 8344
rect 8426 8313 8438 8316
rect 8380 8307 8438 8313
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 9784 8276 9812 8375
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 13541 8347 13599 8353
rect 13541 8313 13553 8347
rect 13587 8344 13599 8347
rect 14182 8344 14188 8356
rect 13587 8316 14188 8344
rect 13587 8313 13599 8316
rect 13541 8307 13599 8313
rect 14182 8304 14188 8316
rect 14240 8304 14246 8356
rect 14844 8344 14872 8511
rect 18598 8508 18604 8560
rect 18656 8548 18662 8560
rect 18656 8520 19472 8548
rect 18656 8508 18662 8520
rect 18966 8480 18972 8492
rect 18927 8452 18972 8480
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19444 8489 19472 8520
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 15841 8415 15899 8421
rect 15841 8381 15853 8415
rect 15887 8412 15899 8415
rect 16108 8415 16166 8421
rect 15887 8384 16068 8412
rect 15887 8381 15899 8384
rect 15841 8375 15899 8381
rect 16040 8356 16068 8384
rect 16108 8381 16120 8415
rect 16154 8412 16166 8415
rect 16666 8412 16672 8424
rect 16154 8384 16672 8412
rect 16154 8381 16166 8384
rect 16108 8375 16166 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 19702 8421 19708 8424
rect 18233 8415 18291 8421
rect 18233 8412 18245 8415
rect 16776 8384 18245 8412
rect 14844 8316 15976 8344
rect 10042 8276 10048 8288
rect 9784 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 12802 8276 12808 8288
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 15948 8276 15976 8316
rect 16022 8304 16028 8356
rect 16080 8304 16086 8356
rect 16776 8344 16804 8384
rect 18233 8381 18245 8384
rect 18279 8381 18291 8415
rect 19696 8412 19708 8421
rect 19663 8384 19708 8412
rect 18233 8375 18291 8381
rect 19696 8375 19708 8384
rect 19702 8372 19708 8375
rect 19760 8372 19766 8424
rect 16132 8316 16804 8344
rect 17497 8347 17555 8353
rect 16132 8276 16160 8316
rect 17497 8313 17509 8347
rect 17543 8344 17555 8347
rect 18506 8344 18512 8356
rect 17543 8316 18512 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 17218 8276 17224 8288
rect 15948 8248 16160 8276
rect 17179 8248 17224 8276
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 18598 8276 18604 8288
rect 18559 8248 18604 8276
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10502 8072 10508 8084
rect 10463 8044 10508 8072
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 11698 8072 11704 8084
rect 11563 8044 11704 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 13998 8072 14004 8084
rect 13959 8044 14004 8072
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 14366 8072 14372 8084
rect 14327 8044 14372 8072
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 16206 8072 16212 8084
rect 15335 8044 16212 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 18564 8044 18613 8072
rect 18564 8032 18570 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 20312 8044 21281 8072
rect 20312 8032 20318 8044
rect 21269 8041 21281 8044
rect 21315 8041 21327 8075
rect 21269 8035 21327 8041
rect 10321 8007 10379 8013
rect 10321 7973 10333 8007
rect 10367 8004 10379 8007
rect 10873 8007 10931 8013
rect 10873 8004 10885 8007
rect 10367 7976 10885 8004
rect 10367 7973 10379 7976
rect 10321 7967 10379 7973
rect 10873 7973 10885 7976
rect 10919 7973 10931 8007
rect 10873 7967 10931 7973
rect 10962 7964 10968 8016
rect 11020 7964 11026 8016
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7936 10287 7939
rect 10413 7939 10471 7945
rect 10413 7936 10425 7939
rect 10275 7908 10425 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10413 7905 10425 7908
rect 10459 7905 10471 7939
rect 10980 7936 11008 7964
rect 10980 7908 11100 7936
rect 10413 7899 10471 7905
rect 11072 7877 11100 7908
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11756 7908 11897 7936
rect 11756 7896 11762 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 12860 7908 13369 7936
rect 12860 7896 12866 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 13357 7899 13415 7905
rect 15212 7908 15669 7936
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 9355 7840 10977 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11974 7868 11980 7880
rect 11935 7840 11980 7868
rect 11057 7831 11115 7837
rect 10980 7800 11008 7831
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7868 12219 7871
rect 12526 7868 12532 7880
rect 12207 7840 12532 7868
rect 12207 7837 12219 7840
rect 12161 7831 12219 7837
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 13320 7840 13461 7868
rect 13320 7828 13326 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 14461 7871 14519 7877
rect 13596 7840 13641 7868
rect 13596 7828 13602 7840
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 14734 7868 14740 7880
rect 14691 7840 14740 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 11238 7800 11244 7812
rect 10980 7772 11244 7800
rect 11238 7760 11244 7772
rect 11296 7800 11302 7812
rect 11790 7800 11796 7812
rect 11296 7772 11796 7800
rect 11296 7760 11302 7772
rect 11790 7760 11796 7772
rect 11848 7760 11854 7812
rect 12989 7803 13047 7809
rect 12989 7769 13001 7803
rect 13035 7800 13047 7803
rect 14476 7800 14504 7831
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 13035 7772 14504 7800
rect 13035 7769 13047 7772
rect 12989 7763 13047 7769
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 8996 7704 9689 7732
rect 8996 7692 9002 7704
rect 9677 7701 9689 7704
rect 9723 7732 9735 7735
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 9723 7704 10333 7732
rect 9723 7701 9735 7704
rect 9677 7695 9735 7701
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 10413 7735 10471 7741
rect 10413 7701 10425 7735
rect 10459 7732 10471 7735
rect 12066 7732 12072 7744
rect 10459 7704 12072 7732
rect 10459 7701 10471 7704
rect 10413 7695 10471 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 12621 7735 12679 7741
rect 12621 7732 12633 7735
rect 12400 7704 12633 7732
rect 12400 7692 12406 7704
rect 12621 7701 12633 7704
rect 12667 7732 12679 7735
rect 15212 7732 15240 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16844 7939 16902 7945
rect 15804 7908 15849 7936
rect 15804 7896 15810 7908
rect 16844 7905 16856 7939
rect 16890 7936 16902 7939
rect 17218 7936 17224 7948
rect 16890 7908 17224 7936
rect 16890 7905 16902 7908
rect 16844 7899 16902 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 20165 7939 20223 7945
rect 20165 7936 20177 7939
rect 19944 7908 20177 7936
rect 19944 7896 19950 7908
rect 20165 7905 20177 7908
rect 20211 7936 20223 7939
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 20211 7908 20913 7936
rect 20211 7905 20223 7908
rect 20165 7899 20223 7905
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 15838 7868 15844 7880
rect 15799 7840 15844 7868
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 16574 7868 16580 7880
rect 16080 7840 16580 7868
rect 16080 7828 16086 7840
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 19337 7871 19395 7877
rect 18831 7840 19012 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 18233 7803 18291 7809
rect 18233 7769 18245 7803
rect 18279 7800 18291 7803
rect 18874 7800 18880 7812
rect 18279 7772 18880 7800
rect 18279 7769 18291 7772
rect 18233 7763 18291 7769
rect 18874 7760 18880 7772
rect 18932 7760 18938 7812
rect 12667 7704 15240 7732
rect 12667 7701 12679 7704
rect 12621 7695 12679 7701
rect 17862 7692 17868 7744
rect 17920 7732 17926 7744
rect 17957 7735 18015 7741
rect 17957 7732 17969 7735
rect 17920 7704 17969 7732
rect 17920 7692 17926 7704
rect 17957 7701 17969 7704
rect 18003 7732 18015 7735
rect 18984 7732 19012 7840
rect 19337 7837 19349 7871
rect 19383 7868 19395 7871
rect 19702 7868 19708 7880
rect 19383 7840 19708 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 20254 7868 20260 7880
rect 20215 7840 20260 7868
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7868 20499 7871
rect 20622 7868 20628 7880
rect 20487 7840 20628 7868
rect 20487 7837 20499 7840
rect 20441 7831 20499 7837
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 19794 7732 19800 7744
rect 18003 7704 19012 7732
rect 19755 7704 19800 7732
rect 18003 7701 18015 7704
rect 17957 7695 18015 7701
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 8846 7528 8852 7540
rect 8807 7500 8852 7528
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 10597 7531 10655 7537
rect 10597 7497 10609 7531
rect 10643 7528 10655 7531
rect 11974 7528 11980 7540
rect 10643 7500 11980 7528
rect 10643 7497 10655 7500
rect 10597 7491 10655 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 13872 7500 14105 7528
rect 13872 7488 13878 7500
rect 14093 7497 14105 7500
rect 14139 7497 14151 7531
rect 14093 7491 14151 7497
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 16758 7528 16764 7540
rect 15887 7500 16764 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 16853 7531 16911 7537
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 18690 7528 18696 7540
rect 16899 7500 18696 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 20070 7488 20076 7540
rect 20128 7528 20134 7540
rect 20349 7531 20407 7537
rect 20349 7528 20361 7531
rect 20128 7500 20361 7528
rect 20128 7488 20134 7500
rect 20349 7497 20361 7500
rect 20395 7497 20407 7531
rect 20349 7491 20407 7497
rect 18601 7463 18659 7469
rect 18601 7429 18613 7463
rect 18647 7460 18659 7463
rect 20254 7460 20260 7472
rect 18647 7432 20260 7460
rect 18647 7429 18659 7432
rect 18601 7423 18659 7429
rect 20254 7420 20260 7432
rect 20312 7420 20318 7472
rect 9398 7392 9404 7404
rect 9359 7364 9404 7392
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 11146 7392 11152 7404
rect 11107 7364 11152 7392
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11698 7392 11704 7404
rect 11659 7364 11704 7392
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12434 7392 12440 7404
rect 12395 7364 12440 7392
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 13964 7364 14657 7392
rect 13964 7352 13970 7364
rect 14645 7361 14657 7364
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 16666 7392 16672 7404
rect 16531 7364 16672 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17276 7364 17417 7392
rect 17276 7352 17282 7364
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 19794 7392 19800 7404
rect 19755 7364 19800 7392
rect 17405 7355 17463 7361
rect 19794 7352 19800 7364
rect 19852 7352 19858 7404
rect 19978 7392 19984 7404
rect 19939 7364 19984 7392
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20901 7395 20959 7401
rect 20901 7392 20913 7395
rect 20220 7364 20913 7392
rect 20220 7352 20226 7364
rect 20901 7361 20913 7364
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7324 11115 7327
rect 11238 7324 11244 7336
rect 11103 7296 11244 7324
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 12452 7324 12480 7352
rect 11388 7296 12480 7324
rect 11388 7284 11394 7296
rect 12526 7284 12532 7336
rect 12584 7324 12590 7336
rect 12693 7327 12751 7333
rect 12693 7324 12705 7327
rect 12584 7296 12705 7324
rect 12584 7284 12590 7296
rect 12693 7293 12705 7296
rect 12739 7293 12751 7327
rect 12693 7287 12751 7293
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 17954 7324 17960 7336
rect 15151 7296 17960 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 19702 7324 19708 7336
rect 19663 7296 19708 7324
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 9217 7259 9275 7265
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 9861 7259 9919 7265
rect 9861 7256 9873 7259
rect 9263 7228 9873 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 9861 7225 9873 7228
rect 9907 7225 9919 7259
rect 14458 7256 14464 7268
rect 14419 7228 14464 7256
rect 9861 7219 9919 7225
rect 14458 7216 14464 7228
rect 14516 7216 14522 7268
rect 14642 7216 14648 7268
rect 14700 7256 14706 7268
rect 15381 7259 15439 7265
rect 15381 7256 15393 7259
rect 14700 7228 15393 7256
rect 14700 7216 14706 7228
rect 15381 7225 15393 7228
rect 15427 7225 15439 7259
rect 18049 7259 18107 7265
rect 18049 7256 18061 7259
rect 15381 7219 15439 7225
rect 17236 7228 18061 7256
rect 17236 7200 17264 7228
rect 18049 7225 18061 7228
rect 18095 7225 18107 7259
rect 18049 7219 18107 7225
rect 19518 7216 19524 7268
rect 19576 7256 19582 7268
rect 20809 7259 20867 7265
rect 20809 7256 20821 7259
rect 19576 7228 20821 7256
rect 19576 7216 19582 7228
rect 20809 7225 20821 7228
rect 20855 7225 20867 7259
rect 20809 7219 20867 7225
rect 9306 7188 9312 7200
rect 9267 7160 9312 7188
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 10928 7160 10977 7188
rect 10928 7148 10934 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 13906 7188 13912 7200
rect 13863 7160 13912 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14550 7188 14556 7200
rect 14511 7160 14556 7188
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 16206 7188 16212 7200
rect 16167 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 17218 7188 17224 7200
rect 16356 7160 16401 7188
rect 17179 7160 17224 7188
rect 16356 7148 16362 7160
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 17313 7191 17371 7197
rect 17313 7157 17325 7191
rect 17359 7188 17371 7191
rect 18138 7188 18144 7200
rect 17359 7160 18144 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 18138 7148 18144 7160
rect 18196 7188 18202 7200
rect 18874 7188 18880 7200
rect 18196 7160 18880 7188
rect 18196 7148 18202 7160
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 19061 7191 19119 7197
rect 19061 7157 19073 7191
rect 19107 7188 19119 7191
rect 19150 7188 19156 7200
rect 19107 7160 19156 7188
rect 19107 7157 19119 7160
rect 19061 7151 19119 7157
rect 19150 7148 19156 7160
rect 19208 7148 19214 7200
rect 19337 7191 19395 7197
rect 19337 7157 19349 7191
rect 19383 7188 19395 7191
rect 20070 7188 20076 7200
rect 19383 7160 20076 7188
rect 19383 7157 19395 7160
rect 19337 7151 19395 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20714 7188 20720 7200
rect 20675 7160 20720 7188
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 9309 6987 9367 6993
rect 9309 6953 9321 6987
rect 9355 6984 9367 6987
rect 9398 6984 9404 6996
rect 9355 6956 9404 6984
rect 9355 6953 9367 6956
rect 9309 6947 9367 6953
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 11057 6987 11115 6993
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11146 6984 11152 6996
rect 11103 6956 11152 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 12713 6987 12771 6993
rect 12713 6984 12725 6987
rect 12584 6956 12725 6984
rect 12584 6944 12590 6956
rect 12713 6953 12725 6956
rect 12759 6953 12771 6987
rect 16666 6984 16672 6996
rect 16627 6956 16672 6984
rect 12713 6947 12771 6953
rect 16666 6944 16672 6956
rect 16724 6944 16730 6996
rect 19978 6944 19984 6996
rect 20036 6984 20042 6996
rect 20441 6987 20499 6993
rect 20441 6984 20453 6987
rect 20036 6956 20453 6984
rect 20036 6944 20042 6956
rect 20441 6953 20453 6956
rect 20487 6953 20499 6987
rect 20441 6947 20499 6953
rect 8196 6851 8254 6857
rect 8196 6817 8208 6851
rect 8242 6848 8254 6851
rect 8754 6848 8760 6860
rect 8242 6820 8760 6848
rect 8242 6817 8254 6820
rect 8196 6811 8254 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 9416 6848 9444 6944
rect 9933 6851 9991 6857
rect 9933 6848 9945 6851
rect 9416 6820 9945 6848
rect 9933 6817 9945 6820
rect 9979 6817 9991 6851
rect 11164 6848 11192 6944
rect 15488 6888 16160 6916
rect 11589 6851 11647 6857
rect 11589 6848 11601 6851
rect 11164 6820 11601 6848
rect 9933 6811 9991 6817
rect 11589 6817 11601 6820
rect 11635 6817 11647 6851
rect 11589 6811 11647 6817
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 12492 6820 13369 6848
rect 12492 6808 12498 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 13624 6851 13682 6857
rect 13624 6817 13636 6851
rect 13670 6848 13682 6851
rect 15289 6851 15347 6857
rect 13670 6820 15240 6848
rect 13670 6817 13682 6820
rect 13624 6811 13682 6817
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 11330 6780 11336 6792
rect 11291 6752 11336 6780
rect 9677 6743 9735 6749
rect 7944 6644 7972 6743
rect 9692 6644 9720 6743
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11348 6644 11376 6740
rect 7944 6616 11376 6644
rect 13081 6647 13139 6653
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 13262 6644 13268 6656
rect 13127 6616 13268 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 13262 6604 13268 6616
rect 13320 6644 13326 6656
rect 14550 6644 14556 6656
rect 13320 6616 14556 6644
rect 13320 6604 13326 6616
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 14734 6644 14740 6656
rect 14695 6616 14740 6644
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 15212 6644 15240 6820
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 15488 6848 15516 6888
rect 15335 6820 15516 6848
rect 15556 6851 15614 6857
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15556 6817 15568 6851
rect 15602 6848 15614 6851
rect 16022 6848 16028 6860
rect 15602 6820 16028 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16132 6848 16160 6888
rect 16574 6848 16580 6860
rect 16132 6820 16580 6848
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16684 6848 16712 6944
rect 19150 6876 19156 6928
rect 19208 6916 19214 6928
rect 19208 6888 19288 6916
rect 19208 6876 19214 6888
rect 17201 6851 17259 6857
rect 17201 6848 17213 6851
rect 16684 6820 17213 6848
rect 17201 6817 17213 6820
rect 17247 6817 17259 6851
rect 17201 6811 17259 6817
rect 17586 6808 17592 6860
rect 17644 6848 17650 6860
rect 19058 6857 19064 6860
rect 18785 6851 18843 6857
rect 18785 6848 18797 6851
rect 17644 6820 18797 6848
rect 17644 6808 17650 6820
rect 18785 6817 18797 6820
rect 18831 6817 18843 6851
rect 18785 6811 18843 6817
rect 19052 6811 19064 6857
rect 19116 6848 19122 6860
rect 19260 6848 19288 6888
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 19116 6820 19152 6848
rect 19260 6820 20913 6848
rect 19058 6808 19064 6811
rect 19116 6808 19122 6820
rect 20901 6817 20913 6820
rect 20947 6848 20959 6851
rect 22005 6851 22063 6857
rect 22005 6848 22017 6851
rect 20947 6820 22017 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 22005 6817 22017 6820
rect 22051 6817 22063 6851
rect 22005 6811 22063 6817
rect 16592 6780 16620 6808
rect 16942 6780 16948 6792
rect 16592 6752 16948 6780
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 20162 6712 20168 6724
rect 20123 6684 20168 6712
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 17862 6644 17868 6656
rect 15212 6616 17868 6644
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 18196 6616 18337 6644
rect 18196 6604 18202 6616
rect 18325 6613 18337 6616
rect 18371 6613 18383 6647
rect 18325 6607 18383 6613
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 20680 6616 21097 6644
rect 20680 6604 20686 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8812 6412 8861 6440
rect 8812 6400 8818 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9306 6440 9312 6452
rect 9171 6412 9312 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 8864 6304 8892 6403
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 10594 6440 10600 6452
rect 10555 6412 10600 6440
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 13078 6440 13084 6452
rect 13039 6412 13084 6440
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 16022 6440 16028 6452
rect 15983 6412 16028 6440
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 16298 6440 16304 6452
rect 16259 6412 16304 6440
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 18064 6412 19012 6440
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 8864 6276 9689 6304
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 11146 6304 11152 6316
rect 11107 6276 11152 6304
rect 9677 6267 9735 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 13722 6304 13728 6316
rect 13683 6276 13728 6304
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 16022 6264 16028 6316
rect 16080 6304 16086 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16080 6276 16865 6304
rect 16080 6264 16086 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6236 7527 6239
rect 8202 6236 8208 6248
rect 7515 6208 8208 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6236 12679 6239
rect 13630 6236 13636 6248
rect 12667 6208 13636 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 14912 6239 14970 6245
rect 14912 6205 14924 6239
rect 14958 6236 14970 6239
rect 16482 6236 16488 6248
rect 14958 6208 16488 6236
rect 14958 6205 14970 6208
rect 14912 6199 14970 6205
rect 7736 6171 7794 6177
rect 7736 6137 7748 6171
rect 7782 6168 7794 6171
rect 8294 6168 8300 6180
rect 7782 6140 8300 6168
rect 7782 6137 7794 6140
rect 7736 6131 7794 6137
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 9490 6168 9496 6180
rect 9451 6140 9496 6168
rect 9490 6128 9496 6140
rect 9548 6128 9554 6180
rect 10686 6128 10692 6180
rect 10744 6168 10750 6180
rect 11057 6171 11115 6177
rect 11057 6168 11069 6171
rect 10744 6140 11069 6168
rect 10744 6128 10750 6140
rect 11057 6137 11069 6140
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 14093 6171 14151 6177
rect 14093 6168 14105 6171
rect 13964 6140 14105 6168
rect 13964 6128 13970 6140
rect 14093 6137 14105 6140
rect 14139 6168 14151 6171
rect 14458 6168 14464 6180
rect 14139 6140 14464 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 14660 6168 14688 6199
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 16666 6236 16672 6248
rect 16627 6208 16672 6236
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 17494 6236 17500 6248
rect 17455 6208 17500 6236
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 18064 6245 18092 6412
rect 18984 6372 19012 6412
rect 19058 6400 19064 6452
rect 19116 6440 19122 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19116 6412 19441 6440
rect 19116 6400 19122 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 18984 6344 19840 6372
rect 19812 6313 19840 6344
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17604 6208 18061 6236
rect 14660 6140 16988 6168
rect 16960 6112 16988 6140
rect 17604 6112 17632 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18138 6196 18144 6248
rect 18196 6236 18202 6248
rect 18305 6239 18363 6245
rect 18305 6236 18317 6239
rect 18196 6208 18317 6236
rect 18196 6196 18202 6208
rect 18305 6205 18317 6208
rect 18351 6236 18363 6239
rect 18351 6208 19748 6236
rect 18351 6205 18363 6208
rect 18305 6199 18363 6205
rect 9582 6100 9588 6112
rect 9543 6072 9588 6100
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 9732 6072 10241 6100
rect 9732 6060 9738 6072
rect 10229 6069 10241 6072
rect 10275 6100 10287 6103
rect 10870 6100 10876 6112
rect 10275 6072 10876 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 10965 6103 11023 6109
rect 10965 6069 10977 6103
rect 11011 6100 11023 6103
rect 11238 6100 11244 6112
rect 11011 6072 11244 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11698 6100 11704 6112
rect 11659 6072 11704 6100
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 11977 6103 12035 6109
rect 11977 6100 11989 6103
rect 11848 6072 11989 6100
rect 11848 6060 11854 6072
rect 11977 6069 11989 6072
rect 12023 6069 12035 6103
rect 11977 6063 12035 6069
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 12124 6072 12449 6100
rect 12124 6060 12130 6072
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 12768 6072 13461 6100
rect 12768 6060 12774 6072
rect 13449 6069 13461 6072
rect 13495 6069 13507 6103
rect 13449 6063 13507 6069
rect 13541 6103 13599 6109
rect 13541 6069 13553 6103
rect 13587 6100 13599 6103
rect 13998 6100 14004 6112
rect 13587 6072 14004 6100
rect 13587 6069 13599 6072
rect 13541 6063 13599 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 16758 6100 16764 6112
rect 16719 6072 16764 6100
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 17313 6103 17371 6109
rect 17313 6100 17325 6103
rect 17000 6072 17325 6100
rect 17000 6060 17006 6072
rect 17313 6069 17325 6072
rect 17359 6100 17371 6103
rect 17586 6100 17592 6112
rect 17359 6072 17592 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 19720 6100 19748 6208
rect 20064 6171 20122 6177
rect 20064 6137 20076 6171
rect 20110 6168 20122 6171
rect 20162 6168 20168 6180
rect 20110 6140 20168 6168
rect 20110 6137 20122 6140
rect 20064 6131 20122 6137
rect 20162 6128 20168 6140
rect 20220 6128 20226 6180
rect 20346 6100 20352 6112
rect 19720 6072 20352 6100
rect 20346 6060 20352 6072
rect 20404 6060 20410 6112
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 21177 6103 21235 6109
rect 21177 6100 21189 6103
rect 20496 6072 21189 6100
rect 20496 6060 20502 6072
rect 21177 6069 21189 6072
rect 21223 6069 21235 6103
rect 21177 6063 21235 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 8386 5896 8392 5908
rect 7699 5868 8392 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 13998 5896 14004 5908
rect 13959 5868 14004 5896
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 14424 5868 14473 5896
rect 14424 5856 14430 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5896 15347 5899
rect 16206 5896 16212 5908
rect 15335 5868 16212 5896
rect 15335 5865 15347 5868
rect 15289 5859 15347 5865
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 16393 5899 16451 5905
rect 16393 5865 16405 5899
rect 16439 5896 16451 5899
rect 16666 5896 16672 5908
rect 16439 5868 16672 5896
rect 16439 5865 16451 5868
rect 16393 5859 16451 5865
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 16761 5899 16819 5905
rect 16761 5865 16773 5899
rect 16807 5896 16819 5899
rect 17862 5896 17868 5908
rect 16807 5868 17868 5896
rect 16807 5865 16819 5868
rect 16761 5859 16819 5865
rect 9950 5828 9956 5840
rect 7944 5800 9956 5828
rect 7377 5763 7435 5769
rect 7377 5729 7389 5763
rect 7423 5760 7435 5763
rect 7558 5760 7564 5772
rect 7423 5732 7564 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 7558 5720 7564 5732
rect 7616 5760 7622 5772
rect 7944 5760 7972 5800
rect 9950 5788 9956 5800
rect 10008 5788 10014 5840
rect 12612 5831 12670 5837
rect 10152 5800 12388 5828
rect 7616 5732 7972 5760
rect 8021 5763 8079 5769
rect 7616 5720 7622 5732
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8665 5763 8723 5769
rect 8665 5760 8677 5763
rect 8067 5732 8677 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8665 5729 8677 5732
rect 8711 5729 8723 5763
rect 8665 5723 8723 5729
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10152 5769 10180 5800
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 10100 5732 10149 5760
rect 10100 5720 10106 5732
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10404 5763 10462 5769
rect 10404 5729 10416 5763
rect 10450 5760 10462 5763
rect 11146 5760 11152 5772
rect 10450 5732 11152 5760
rect 10450 5729 10462 5732
rect 10404 5723 10462 5729
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 12360 5769 12388 5800
rect 12612 5797 12624 5831
rect 12658 5828 12670 5831
rect 13354 5828 13360 5840
rect 12658 5800 13360 5828
rect 12658 5797 12670 5800
rect 12612 5791 12670 5797
rect 13354 5788 13360 5800
rect 13412 5828 13418 5840
rect 13412 5800 14688 5828
rect 13412 5788 13418 5800
rect 12345 5763 12403 5769
rect 12345 5729 12357 5763
rect 12391 5760 12403 5763
rect 12434 5760 12440 5772
rect 12391 5732 12440 5760
rect 12391 5729 12403 5732
rect 12345 5723 12403 5729
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 14090 5720 14096 5772
rect 14148 5760 14154 5772
rect 14369 5763 14427 5769
rect 14369 5760 14381 5763
rect 14148 5732 14381 5760
rect 14148 5720 14154 5732
rect 14369 5729 14381 5732
rect 14415 5729 14427 5763
rect 14369 5723 14427 5729
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7248 5664 8125 5692
rect 7248 5652 7254 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8294 5692 8300 5704
rect 8251 5664 8300 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 14384 5624 14412 5723
rect 14660 5701 14688 5800
rect 15746 5788 15752 5840
rect 15804 5828 15810 5840
rect 16776 5828 16804 5859
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 19245 5899 19303 5905
rect 19245 5865 19257 5899
rect 19291 5896 19303 5899
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 19291 5868 19809 5896
rect 19291 5865 19303 5868
rect 19245 5859 19303 5865
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 19797 5859 19855 5865
rect 15804 5800 16804 5828
rect 15804 5788 15810 5800
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5692 14703 5695
rect 14734 5692 14740 5704
rect 14691 5664 14740 5692
rect 14691 5661 14703 5664
rect 14645 5655 14703 5661
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 15470 5624 15476 5636
rect 13280 5596 13860 5624
rect 14384 5596 15476 5624
rect 9122 5556 9128 5568
rect 9083 5528 9128 5556
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9677 5559 9735 5565
rect 9677 5556 9689 5559
rect 9548 5528 9689 5556
rect 9548 5516 9554 5528
rect 9677 5525 9689 5528
rect 9723 5525 9735 5559
rect 9677 5519 9735 5525
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 11112 5528 11529 5556
rect 11112 5516 11118 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 12066 5556 12072 5568
rect 11979 5528 12072 5556
rect 11517 5519 11575 5525
rect 12066 5516 12072 5528
rect 12124 5556 12130 5568
rect 13280 5556 13308 5596
rect 13722 5556 13728 5568
rect 12124 5528 13308 5556
rect 13683 5528 13728 5556
rect 12124 5516 12130 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 13832 5556 13860 5596
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 15856 5556 15884 5800
rect 17770 5788 17776 5840
rect 17828 5828 17834 5840
rect 20257 5831 20315 5837
rect 20257 5828 20269 5831
rect 17828 5800 20269 5828
rect 17828 5788 17834 5800
rect 20257 5797 20269 5800
rect 20303 5797 20315 5831
rect 20257 5791 20315 5797
rect 17497 5763 17555 5769
rect 17497 5729 17509 5763
rect 17543 5760 17555 5763
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 17543 5732 18245 5760
rect 17543 5729 17555 5732
rect 17497 5723 17555 5729
rect 18233 5729 18245 5732
rect 18279 5760 18291 5763
rect 18690 5760 18696 5772
rect 18279 5732 18696 5760
rect 18279 5729 18291 5732
rect 18233 5723 18291 5729
rect 18690 5720 18696 5732
rect 18748 5720 18754 5772
rect 19153 5763 19211 5769
rect 19153 5729 19165 5763
rect 19199 5760 19211 5763
rect 19978 5760 19984 5772
rect 19199 5732 19984 5760
rect 19199 5729 19211 5732
rect 19153 5723 19211 5729
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 20165 5763 20223 5769
rect 20165 5729 20177 5763
rect 20211 5760 20223 5763
rect 20898 5760 20904 5772
rect 20211 5732 20576 5760
rect 20859 5732 20904 5760
rect 20211 5729 20223 5732
rect 20165 5723 20223 5729
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 16022 5692 16028 5704
rect 15979 5664 16028 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16850 5692 16856 5704
rect 16811 5664 16856 5692
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5661 17003 5695
rect 16945 5655 17003 5661
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5692 17831 5695
rect 18966 5692 18972 5704
rect 17819 5664 18972 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 16960 5624 16988 5655
rect 18966 5652 18972 5664
rect 19024 5652 19030 5704
rect 19058 5652 19064 5704
rect 19116 5692 19122 5704
rect 19337 5695 19395 5701
rect 19337 5692 19349 5695
rect 19116 5664 19349 5692
rect 19116 5652 19122 5664
rect 19337 5661 19349 5664
rect 19383 5661 19395 5695
rect 19337 5655 19395 5661
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20548 5692 20576 5732
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21634 5692 21640 5704
rect 20404 5664 20449 5692
rect 20548 5664 21640 5692
rect 20404 5652 20410 5664
rect 21634 5652 21640 5664
rect 21692 5652 21698 5704
rect 16540 5596 16988 5624
rect 18785 5627 18843 5633
rect 16540 5584 16546 5596
rect 18785 5593 18797 5627
rect 18831 5624 18843 5627
rect 19518 5624 19524 5636
rect 18831 5596 19524 5624
rect 18831 5593 18843 5596
rect 18785 5587 18843 5593
rect 19518 5584 19524 5596
rect 19576 5584 19582 5636
rect 21542 5624 21548 5636
rect 20916 5596 21548 5624
rect 13832 5528 15884 5556
rect 18417 5559 18475 5565
rect 18417 5525 18429 5559
rect 18463 5556 18475 5559
rect 20916 5556 20944 5596
rect 21542 5584 21548 5596
rect 21600 5584 21606 5636
rect 21082 5556 21088 5568
rect 18463 5528 20944 5556
rect 21043 5528 21088 5556
rect 18463 5525 18475 5528
rect 18417 5519 18475 5525
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 22002 5556 22008 5568
rect 21963 5528 22008 5556
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8352 5324 8493 5352
rect 8352 5312 8358 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9030 5352 9036 5364
rect 8803 5324 9036 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11425 5355 11483 5361
rect 11425 5352 11437 5355
rect 11204 5324 11437 5352
rect 11204 5312 11210 5324
rect 11425 5321 11437 5324
rect 11471 5321 11483 5355
rect 11425 5315 11483 5321
rect 14921 5355 14979 5361
rect 14921 5321 14933 5355
rect 14967 5352 14979 5355
rect 15746 5352 15752 5364
rect 14967 5324 15752 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16393 5355 16451 5361
rect 16393 5321 16405 5355
rect 16439 5352 16451 5355
rect 16758 5352 16764 5364
rect 16439 5324 16764 5352
rect 16439 5321 16451 5324
rect 16393 5315 16451 5321
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 16850 5312 16856 5364
rect 16908 5352 16914 5364
rect 19150 5352 19156 5364
rect 16908 5324 19156 5352
rect 16908 5312 16914 5324
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 19978 5352 19984 5364
rect 19939 5324 19984 5352
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 17681 5287 17739 5293
rect 15580 5256 16528 5284
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 9272 5188 9321 5216
rect 9272 5176 9278 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 10042 5216 10048 5228
rect 10003 5188 10048 5216
rect 9309 5179 9367 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 15580 5225 15608 5256
rect 16500 5228 16528 5256
rect 17681 5253 17693 5287
rect 17727 5284 17739 5287
rect 17954 5284 17960 5296
rect 17727 5256 17960 5284
rect 17727 5253 17739 5256
rect 17681 5247 17739 5253
rect 17954 5244 17960 5256
rect 18012 5244 18018 5296
rect 18877 5287 18935 5293
rect 18877 5253 18889 5287
rect 18923 5284 18935 5287
rect 20806 5284 20812 5296
rect 18923 5256 20812 5284
rect 18923 5253 18935 5256
rect 18877 5247 18935 5253
rect 20806 5244 20812 5256
rect 20864 5244 20870 5296
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11296 5188 11713 5216
rect 11296 5176 11302 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 15565 5219 15623 5225
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 15654 5176 15660 5228
rect 15712 5216 15718 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15712 5188 15945 5216
rect 15712 5176 15718 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16540 5188 16957 5216
rect 16540 5176 16546 5188
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 19058 5176 19064 5228
rect 19116 5216 19122 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19116 5188 19441 5216
rect 19116 5176 19122 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 20346 5176 20352 5228
rect 20404 5216 20410 5228
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 20404 5188 20545 5216
rect 20404 5176 20410 5188
rect 20533 5185 20545 5188
rect 20579 5185 20591 5219
rect 20533 5179 20591 5185
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 8202 5148 8208 5160
rect 7147 5120 8208 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 8202 5108 8208 5120
rect 8260 5148 8266 5160
rect 10060 5148 10088 5176
rect 11054 5148 11060 5160
rect 8260 5120 10088 5148
rect 10152 5120 11060 5148
rect 8260 5108 8266 5120
rect 7368 5083 7426 5089
rect 7368 5049 7380 5083
rect 7414 5080 7426 5083
rect 7742 5080 7748 5092
rect 7414 5052 7748 5080
rect 7414 5049 7426 5052
rect 7368 5043 7426 5049
rect 7742 5040 7748 5052
rect 7800 5080 7806 5092
rect 10152 5080 10180 5120
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12529 5151 12587 5157
rect 12529 5148 12541 5151
rect 12492 5120 12541 5148
rect 12492 5108 12498 5120
rect 12529 5117 12541 5120
rect 12575 5117 12587 5151
rect 12529 5111 12587 5117
rect 12796 5151 12854 5157
rect 12796 5117 12808 5151
rect 12842 5148 12854 5151
rect 13722 5148 13728 5160
rect 12842 5120 13728 5148
rect 12842 5117 12854 5120
rect 12796 5111 12854 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 16853 5151 16911 5157
rect 16853 5148 16865 5151
rect 14424 5120 16865 5148
rect 14424 5108 14430 5120
rect 16853 5117 16865 5120
rect 16899 5148 16911 5151
rect 17126 5148 17132 5160
rect 16899 5120 17132 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 17126 5108 17132 5120
rect 17184 5108 17190 5160
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5148 18383 5151
rect 18598 5148 18604 5160
rect 18371 5120 18604 5148
rect 18371 5117 18383 5120
rect 18325 5111 18383 5117
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 18966 5108 18972 5160
rect 19024 5148 19030 5160
rect 19245 5151 19303 5157
rect 19245 5148 19257 5151
rect 19024 5120 19257 5148
rect 19024 5108 19030 5120
rect 19245 5117 19257 5120
rect 19291 5117 19303 5151
rect 20990 5148 20996 5160
rect 20951 5120 20996 5148
rect 19245 5111 19303 5117
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 7800 5052 10180 5080
rect 10312 5083 10370 5089
rect 7800 5040 7806 5052
rect 10312 5049 10324 5083
rect 10358 5080 10370 5083
rect 10358 5052 11284 5080
rect 10358 5049 10370 5052
rect 10312 5043 10370 5049
rect 11256 5024 11284 5052
rect 16022 5040 16028 5092
rect 16080 5080 16086 5092
rect 19337 5083 19395 5089
rect 19337 5080 19349 5083
rect 16080 5052 19349 5080
rect 16080 5040 16086 5052
rect 19337 5049 19349 5052
rect 19383 5049 19395 5083
rect 19337 5043 19395 5049
rect 20441 5083 20499 5089
rect 20441 5049 20453 5083
rect 20487 5080 20499 5083
rect 21450 5080 21456 5092
rect 20487 5052 21456 5080
rect 20487 5049 20499 5052
rect 20441 5043 20499 5049
rect 21450 5040 21456 5052
rect 21508 5040 21514 5092
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9217 5015 9275 5021
rect 9217 4981 9229 5015
rect 9263 5012 9275 5015
rect 9582 5012 9588 5024
rect 9263 4984 9588 5012
rect 9263 4981 9275 4984
rect 9217 4975 9275 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 11296 4984 13921 5012
rect 11296 4972 11302 4984
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 14182 5012 14188 5024
rect 14143 4984 14188 5012
rect 13909 4975 13967 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 14516 4984 15301 5012
rect 14516 4972 14522 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 15381 5015 15439 5021
rect 15381 4981 15393 5015
rect 15427 5012 15439 5015
rect 15470 5012 15476 5024
rect 15427 4984 15476 5012
rect 15427 4981 15439 4984
rect 15381 4975 15439 4981
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 16482 4972 16488 5024
rect 16540 5012 16546 5024
rect 16761 5015 16819 5021
rect 16761 5012 16773 5015
rect 16540 4984 16773 5012
rect 16540 4972 16546 4984
rect 16761 4981 16773 4984
rect 16807 4981 16819 5015
rect 16761 4975 16819 4981
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 18509 5015 18567 5021
rect 18509 5012 18521 5015
rect 18196 4984 18521 5012
rect 18196 4972 18202 4984
rect 18509 4981 18521 4984
rect 18555 4981 18567 5015
rect 18509 4975 18567 4981
rect 18874 4972 18880 5024
rect 18932 5012 18938 5024
rect 20346 5012 20352 5024
rect 18932 4984 20352 5012
rect 18932 4972 18938 4984
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 21174 5012 21180 5024
rect 21135 4984 21180 5012
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 7190 4808 7196 4820
rect 7151 4780 7196 4808
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 8205 4811 8263 4817
rect 8205 4777 8217 4811
rect 8251 4808 8263 4811
rect 8570 4808 8576 4820
rect 8251 4780 8576 4808
rect 8251 4777 8263 4780
rect 8205 4771 8263 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 10597 4811 10655 4817
rect 10597 4777 10609 4811
rect 10643 4808 10655 4811
rect 10686 4808 10692 4820
rect 10643 4780 10692 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 12710 4808 12716 4820
rect 12671 4780 12716 4808
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13081 4811 13139 4817
rect 13081 4777 13093 4811
rect 13127 4808 13139 4811
rect 14182 4808 14188 4820
rect 13127 4780 14188 4808
rect 13127 4777 13139 4780
rect 13081 4771 13139 4777
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 16850 4808 16856 4820
rect 15519 4780 16856 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 17313 4811 17371 4817
rect 17313 4777 17325 4811
rect 17359 4808 17371 4811
rect 20990 4808 20996 4820
rect 17359 4780 20996 4808
rect 17359 4777 17371 4780
rect 17313 4771 17371 4777
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 5350 4700 5356 4752
rect 5408 4740 5414 4752
rect 5408 4712 8708 4740
rect 5408 4700 5414 4712
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4641 7619 4675
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 7561 4635 7619 4641
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 6917 4471 6975 4477
rect 6917 4468 6929 4471
rect 5500 4440 6929 4468
rect 5500 4428 5506 4440
rect 6917 4437 6929 4440
rect 6963 4468 6975 4471
rect 7576 4468 7604 4635
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 8680 4672 8708 4712
rect 9582 4700 9588 4752
rect 9640 4740 9646 4752
rect 9769 4743 9827 4749
rect 9769 4740 9781 4743
rect 9640 4712 9781 4740
rect 9640 4700 9646 4712
rect 9769 4709 9781 4712
rect 9815 4740 9827 4743
rect 11698 4740 11704 4752
rect 9815 4712 11704 4740
rect 9815 4709 9827 4712
rect 9769 4703 9827 4709
rect 11698 4700 11704 4712
rect 11756 4740 11762 4752
rect 15841 4743 15899 4749
rect 15841 4740 15853 4743
rect 11756 4712 15853 4740
rect 11756 4700 11762 4712
rect 15841 4709 15853 4712
rect 15887 4740 15899 4743
rect 16574 4740 16580 4752
rect 15887 4712 16580 4740
rect 15887 4709 15899 4712
rect 15841 4703 15899 4709
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 17856 4743 17914 4749
rect 17856 4709 17868 4743
rect 17902 4740 17914 4743
rect 19794 4740 19800 4752
rect 17902 4712 19800 4740
rect 17902 4709 17914 4712
rect 17856 4703 17914 4709
rect 19794 4700 19800 4712
rect 19852 4740 19858 4752
rect 19852 4712 20024 4740
rect 19852 4700 19858 4712
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 8680 4644 10241 4672
rect 10229 4641 10241 4644
rect 10275 4672 10287 4675
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10275 4644 10977 4672
rect 10275 4641 10287 4644
rect 10229 4635 10287 4641
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4672 11851 4675
rect 11974 4672 11980 4684
rect 11839 4644 11980 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4672 12495 4675
rect 13173 4675 13231 4681
rect 13173 4672 13185 4675
rect 12483 4644 13185 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 6963 4440 7604 4468
rect 7668 4468 7696 4567
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 8662 4604 8668 4616
rect 7800 4576 7845 4604
rect 8623 4576 8668 4604
rect 7800 4564 7806 4576
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 8846 4604 8852 4616
rect 8807 4576 8852 4604
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 11238 4604 11244 4616
rect 11199 4576 11244 4604
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 8754 4496 8760 4548
rect 8812 4536 8818 4548
rect 11609 4539 11667 4545
rect 8812 4508 11376 4536
rect 8812 4496 8818 4508
rect 8478 4468 8484 4480
rect 7668 4440 8484 4468
rect 6963 4437 6975 4440
rect 6917 4431 6975 4437
rect 8478 4428 8484 4440
rect 8536 4468 8542 4480
rect 9309 4471 9367 4477
rect 9309 4468 9321 4471
rect 8536 4440 9321 4468
rect 8536 4428 8542 4440
rect 9309 4437 9321 4440
rect 9355 4468 9367 4471
rect 11238 4468 11244 4480
rect 9355 4440 11244 4468
rect 9355 4437 9367 4440
rect 9309 4431 9367 4437
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 11348 4468 11376 4508
rect 11609 4505 11621 4539
rect 11655 4536 11667 4539
rect 12434 4536 12440 4548
rect 11655 4508 12440 4536
rect 11655 4505 11667 4508
rect 11609 4499 11667 4505
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 12544 4468 12572 4644
rect 13173 4641 13185 4644
rect 13219 4641 13231 4675
rect 16206 4672 16212 4684
rect 16119 4644 16212 4672
rect 13173 4635 13231 4641
rect 16206 4632 16212 4644
rect 16264 4672 16270 4684
rect 16482 4672 16488 4684
rect 16264 4644 16488 4672
rect 16264 4632 16270 4644
rect 16482 4632 16488 4644
rect 16540 4672 16546 4684
rect 19058 4672 19064 4684
rect 16540 4644 19064 4672
rect 16540 4632 16546 4644
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 19886 4672 19892 4684
rect 19847 4644 19892 4672
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 19996 4672 20024 4712
rect 20901 4675 20959 4681
rect 19996 4644 20116 4672
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4604 13967 4607
rect 14550 4604 14556 4616
rect 13955 4576 14556 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 14550 4564 14556 4576
rect 14608 4604 14614 4616
rect 17034 4604 17040 4616
rect 14608 4576 17040 4604
rect 14608 4564 14614 4576
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 19978 4604 19984 4616
rect 19939 4576 19984 4604
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20088 4613 20116 4644
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 21266 4672 21272 4684
rect 20947 4644 21272 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4573 20131 4607
rect 20073 4567 20131 4573
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 12768 4508 14872 4536
rect 12768 4496 12774 4508
rect 11348 4440 12572 4468
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 14185 4471 14243 4477
rect 14185 4468 14197 4471
rect 13688 4440 14197 4468
rect 13688 4428 13694 4440
rect 14185 4437 14197 4440
rect 14231 4437 14243 4471
rect 14185 4431 14243 4437
rect 14458 4428 14464 4480
rect 14516 4468 14522 4480
rect 14737 4471 14795 4477
rect 14737 4468 14749 4471
rect 14516 4440 14749 4468
rect 14516 4428 14522 4440
rect 14737 4437 14749 4440
rect 14783 4437 14795 4471
rect 14844 4468 14872 4508
rect 16022 4496 16028 4548
rect 16080 4536 16086 4548
rect 16853 4539 16911 4545
rect 16853 4536 16865 4539
rect 16080 4508 16865 4536
rect 16080 4496 16086 4508
rect 16853 4505 16865 4508
rect 16899 4505 16911 4539
rect 16853 4499 16911 4505
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 21085 4539 21143 4545
rect 21085 4536 21097 4539
rect 19392 4508 21097 4536
rect 19392 4496 19398 4508
rect 21085 4505 21097 4508
rect 21131 4505 21143 4539
rect 21085 4499 21143 4505
rect 16577 4471 16635 4477
rect 16577 4468 16589 4471
rect 14844 4440 16589 4468
rect 14737 4431 14795 4437
rect 16577 4437 16589 4440
rect 16623 4468 16635 4471
rect 16666 4468 16672 4480
rect 16623 4440 16672 4468
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17034 4428 17040 4480
rect 17092 4468 17098 4480
rect 18782 4468 18788 4480
rect 17092 4440 18788 4468
rect 17092 4428 17098 4440
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 18966 4468 18972 4480
rect 18927 4440 18972 4468
rect 18966 4428 18972 4440
rect 19024 4428 19030 4480
rect 19518 4468 19524 4480
rect 19479 4440 19524 4468
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 20162 4428 20168 4480
rect 20220 4468 20226 4480
rect 21174 4468 21180 4480
rect 20220 4440 21180 4468
rect 20220 4428 20226 4440
rect 21174 4428 21180 4440
rect 21232 4428 21238 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 7193 4267 7251 4273
rect 7193 4233 7205 4267
rect 7239 4264 7251 4267
rect 7558 4264 7564 4276
rect 7239 4236 7564 4264
rect 7239 4233 7251 4236
rect 7193 4227 7251 4233
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 8938 4264 8944 4276
rect 7852 4236 8944 4264
rect 7852 4128 7880 4236
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 10410 4264 10416 4276
rect 10371 4236 10416 4264
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 11146 4264 11152 4276
rect 10704 4236 11152 4264
rect 10704 4128 10732 4236
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11238 4224 11244 4276
rect 11296 4264 11302 4276
rect 15657 4267 15715 4273
rect 15657 4264 15669 4267
rect 11296 4236 15669 4264
rect 11296 4224 11302 4236
rect 15657 4233 15669 4236
rect 15703 4264 15715 4267
rect 16206 4264 16212 4276
rect 15703 4236 16212 4264
rect 15703 4233 15715 4236
rect 15657 4227 15715 4233
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 18874 4224 18880 4276
rect 18932 4264 18938 4276
rect 18932 4236 19564 4264
rect 18932 4224 18938 4236
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 11517 4199 11575 4205
rect 11517 4196 11529 4199
rect 11112 4168 11529 4196
rect 11112 4156 11118 4168
rect 11517 4165 11529 4168
rect 11563 4196 11575 4199
rect 12710 4196 12716 4208
rect 11563 4168 12716 4196
rect 11563 4165 11575 4168
rect 11517 4159 11575 4165
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 14366 4196 14372 4208
rect 14016 4168 14372 4196
rect 10962 4128 10968 4140
rect 7760 4100 7880 4128
rect 9692 4100 10732 4128
rect 10923 4100 10968 4128
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 5350 4060 5356 4072
rect 3476 4032 5356 4060
rect 3476 4020 3482 4032
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 7760 4060 7788 4100
rect 6236 4032 7788 4060
rect 7837 4063 7895 4069
rect 6236 4020 6242 4032
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 7926 4060 7932 4072
rect 7883 4032 7932 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 9692 4060 9720 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 12066 4128 12072 4140
rect 12027 4100 12072 4128
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 14016 4137 14044 4168
rect 14366 4156 14372 4168
rect 14424 4156 14430 4208
rect 14737 4199 14795 4205
rect 14737 4165 14749 4199
rect 14783 4165 14795 4199
rect 14737 4159 14795 4165
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14752 4128 14780 4159
rect 17954 4156 17960 4208
rect 18012 4196 18018 4208
rect 18322 4196 18328 4208
rect 18012 4168 18328 4196
rect 18012 4156 18018 4168
rect 18322 4156 18328 4168
rect 18380 4156 18386 4208
rect 19536 4196 19564 4236
rect 19794 4224 19800 4276
rect 19852 4264 19858 4276
rect 19889 4267 19947 4273
rect 19889 4264 19901 4267
rect 19852 4236 19901 4264
rect 19852 4224 19858 4236
rect 19889 4233 19901 4236
rect 19935 4233 19947 4267
rect 19889 4227 19947 4233
rect 19978 4224 19984 4276
rect 20036 4264 20042 4276
rect 20165 4267 20223 4273
rect 20165 4264 20177 4267
rect 20036 4236 20177 4264
rect 20036 4224 20042 4236
rect 20165 4233 20177 4236
rect 20211 4233 20223 4267
rect 20165 4227 20223 4233
rect 21634 4196 21640 4208
rect 19536 4168 21640 4196
rect 21634 4156 21640 4168
rect 21692 4156 21698 4208
rect 14148 4100 14193 4128
rect 14384 4100 14780 4128
rect 14148 4088 14154 4100
rect 14384 4072 14412 4100
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 18230 4128 18236 4140
rect 17184 4100 18236 4128
rect 17184 4088 17190 4100
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 20717 4131 20775 4137
rect 20717 4128 20729 4131
rect 20496 4100 20729 4128
rect 20496 4088 20502 4100
rect 20717 4097 20729 4100
rect 20763 4097 20775 4131
rect 21358 4128 21364 4140
rect 21319 4100 21364 4128
rect 20717 4091 20775 4097
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 8444 4032 9720 4060
rect 9769 4063 9827 4069
rect 8444 4020 8450 4032
rect 9769 4029 9781 4063
rect 9815 4060 9827 4063
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9815 4032 10149 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 10137 4029 10149 4032
rect 10183 4060 10195 4063
rect 10686 4060 10692 4072
rect 10183 4032 10692 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10870 4060 10876 4072
rect 10831 4032 10876 4060
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 11238 4060 11244 4072
rect 11072 4032 11244 4060
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 5442 3992 5448 4004
rect 2924 3964 5448 3992
rect 2924 3952 2930 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 8104 3995 8162 4001
rect 8104 3961 8116 3995
rect 8150 3992 8162 3995
rect 8846 3992 8852 4004
rect 8150 3964 8852 3992
rect 8150 3961 8162 3964
rect 8104 3955 8162 3961
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 10781 3995 10839 4001
rect 10781 3961 10793 3995
rect 10827 3992 10839 3995
rect 11072 3992 11100 4032
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12986 4060 12992 4072
rect 12483 4032 12992 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 14366 4020 14372 4072
rect 14424 4020 14430 4072
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4060 14611 4063
rect 14642 4060 14648 4072
rect 14599 4032 14648 4060
rect 14599 4029 14611 4032
rect 14553 4023 14611 4029
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14792 4032 15117 4060
rect 14792 4020 14798 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 15378 4020 15384 4072
rect 15436 4060 15442 4072
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15436 4032 15945 4060
rect 15436 4020 15442 4032
rect 15933 4029 15945 4032
rect 15979 4060 15991 4063
rect 17586 4060 17592 4072
rect 15979 4032 17592 4060
rect 15979 4029 15991 4032
rect 15933 4023 15991 4029
rect 17586 4020 17592 4032
rect 17644 4060 17650 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 17644 4032 18521 4060
rect 17644 4020 17650 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 18776 4063 18834 4069
rect 18776 4029 18788 4063
rect 18822 4060 18834 4063
rect 20456 4060 20484 4088
rect 18822 4032 20484 4060
rect 20533 4063 20591 4069
rect 18822 4029 18834 4032
rect 18776 4023 18834 4029
rect 20533 4029 20545 4063
rect 20579 4060 20591 4063
rect 20806 4060 20812 4072
rect 20579 4032 20812 4060
rect 20579 4029 20591 4032
rect 20533 4023 20591 4029
rect 10827 3964 11100 3992
rect 10827 3961 10839 3964
rect 10781 3955 10839 3961
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 16200 3995 16258 4001
rect 13412 3964 13676 3992
rect 13412 3952 13418 3964
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 12342 3924 12348 3936
rect 5132 3896 12348 3924
rect 5132 3884 5138 3896
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 12483 3896 12541 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12529 3887 12587 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 12989 3927 13047 3933
rect 12989 3893 13001 3927
rect 13035 3924 13047 3927
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 13035 3896 13553 3924
rect 13035 3893 13047 3896
rect 12989 3887 13047 3893
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 13648 3924 13676 3964
rect 16200 3961 16212 3995
rect 16246 3992 16258 3995
rect 16246 3964 18460 3992
rect 16246 3961 16258 3964
rect 16200 3955 16258 3961
rect 13909 3927 13967 3933
rect 13909 3924 13921 3927
rect 13648 3896 13921 3924
rect 13541 3887 13599 3893
rect 13909 3893 13921 3896
rect 13955 3924 13967 3927
rect 15470 3924 15476 3936
rect 13955 3896 15476 3924
rect 13955 3893 13967 3896
rect 13909 3887 13967 3893
rect 15470 3884 15476 3896
rect 15528 3924 15534 3936
rect 17126 3924 17132 3936
rect 15528 3896 17132 3924
rect 15528 3884 15534 3896
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17310 3924 17316 3936
rect 17271 3896 17316 3924
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17586 3924 17592 3936
rect 17547 3896 17592 3924
rect 17586 3884 17592 3896
rect 17644 3924 17650 3936
rect 17770 3924 17776 3936
rect 17644 3896 17776 3924
rect 17644 3884 17650 3896
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18432 3924 18460 3964
rect 18874 3952 18880 4004
rect 18932 3992 18938 4004
rect 20162 3992 20168 4004
rect 18932 3964 20168 3992
rect 18932 3952 18938 3964
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 18966 3924 18972 3936
rect 18432 3896 18972 3924
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 20548 3924 20576 4023
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 19116 3896 20576 3924
rect 20625 3927 20683 3933
rect 19116 3884 19122 3896
rect 20625 3893 20637 3927
rect 20671 3924 20683 3927
rect 20898 3924 20904 3936
rect 20671 3896 20904 3924
rect 20671 3893 20683 3896
rect 20625 3887 20683 3893
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 8754 3720 8760 3732
rect 4028 3692 8760 3720
rect 4028 3680 4034 3692
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8904 3692 9045 3720
rect 8904 3680 8910 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 10652 3692 13124 3720
rect 10652 3680 10658 3692
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 9122 3652 9128 3664
rect 6788 3624 9128 3652
rect 6788 3612 6794 3624
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 10100 3624 11100 3652
rect 10100 3612 10106 3624
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7653 3587 7711 3593
rect 7653 3584 7665 3587
rect 7524 3556 7665 3584
rect 7524 3544 7530 3556
rect 7653 3553 7665 3556
rect 7699 3584 7711 3587
rect 7742 3584 7748 3596
rect 7699 3556 7748 3584
rect 7699 3553 7711 3556
rect 7653 3547 7711 3553
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 7920 3587 7978 3593
rect 7920 3553 7932 3587
rect 7966 3584 7978 3587
rect 8846 3584 8852 3596
rect 7966 3556 8852 3584
rect 7966 3553 7978 3556
rect 7920 3547 7978 3553
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10220 3587 10278 3593
rect 10220 3553 10232 3587
rect 10266 3584 10278 3587
rect 10962 3584 10968 3596
rect 10266 3556 10968 3584
rect 10266 3553 10278 3556
rect 10220 3547 10278 3553
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11072 3584 11100 3624
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11204 3624 11621 3652
rect 11204 3612 11210 3624
rect 11609 3621 11621 3624
rect 11655 3652 11667 3655
rect 12986 3652 12992 3664
rect 11655 3624 12992 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 12986 3612 12992 3624
rect 13044 3612 13050 3664
rect 13096 3652 13124 3692
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13817 3723 13875 3729
rect 13817 3720 13829 3723
rect 13228 3692 13829 3720
rect 13228 3680 13234 3692
rect 13817 3689 13829 3692
rect 13863 3720 13875 3723
rect 14090 3720 14096 3732
rect 13863 3692 14096 3720
rect 13863 3689 13875 3692
rect 13817 3683 13875 3689
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 14185 3723 14243 3729
rect 14185 3689 14197 3723
rect 14231 3720 14243 3723
rect 14274 3720 14280 3732
rect 14231 3692 14280 3720
rect 14231 3689 14243 3692
rect 14185 3683 14243 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 15841 3723 15899 3729
rect 15841 3689 15853 3723
rect 15887 3720 15899 3723
rect 19797 3723 19855 3729
rect 15887 3692 19472 3720
rect 15887 3689 15899 3692
rect 15841 3683 15899 3689
rect 14458 3652 14464 3664
rect 13096 3624 14464 3652
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 15381 3655 15439 3661
rect 15381 3621 15393 3655
rect 15427 3652 15439 3655
rect 17862 3652 17868 3664
rect 15427 3624 17868 3652
rect 15427 3621 15439 3624
rect 15381 3615 15439 3621
rect 12526 3584 12532 3596
rect 11072 3556 12532 3584
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12704 3587 12762 3593
rect 12704 3553 12716 3587
rect 12750 3584 12762 3587
rect 14550 3584 14556 3596
rect 12750 3556 14228 3584
rect 14511 3556 14556 3584
rect 12750 3553 12762 3556
rect 12704 3547 12762 3553
rect 11974 3516 11980 3528
rect 11935 3488 11980 3516
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12434 3516 12440 3528
rect 12395 3488 12440 3516
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 14200 3516 14228 3556
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 15286 3584 15292 3596
rect 14691 3556 15292 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15672 3593 15700 3624
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 18877 3655 18935 3661
rect 18877 3652 18889 3655
rect 18288 3624 18889 3652
rect 18288 3612 18294 3624
rect 18877 3621 18889 3624
rect 18923 3652 18935 3655
rect 19058 3652 19064 3664
rect 18923 3624 19064 3652
rect 18923 3621 18935 3624
rect 18877 3615 18935 3621
rect 19058 3612 19064 3624
rect 19116 3612 19122 3664
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3553 15715 3587
rect 15657 3547 15715 3553
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 16540 3556 16589 3584
rect 16540 3544 16546 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 17586 3584 17592 3596
rect 16724 3556 17592 3584
rect 16724 3544 16730 3556
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3584 17739 3587
rect 17770 3584 17776 3596
rect 17727 3556 17776 3584
rect 17727 3553 17739 3556
rect 17681 3547 17739 3553
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 18785 3587 18843 3593
rect 18785 3584 18797 3587
rect 17972 3556 18797 3584
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14200 3488 14749 3516
rect 14737 3485 14749 3488
rect 14783 3516 14795 3519
rect 15102 3516 15108 3528
rect 14783 3488 15108 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 16850 3516 16856 3528
rect 16763 3488 16856 3516
rect 16850 3476 16856 3488
rect 16908 3516 16914 3528
rect 17310 3516 17316 3528
rect 16908 3488 17316 3516
rect 16908 3476 16914 3488
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 13814 3408 13820 3460
rect 13872 3448 13878 3460
rect 14366 3448 14372 3460
rect 13872 3420 14372 3448
rect 13872 3408 13878 3420
rect 14366 3408 14372 3420
rect 14424 3408 14430 3460
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 17865 3451 17923 3457
rect 17865 3448 17877 3451
rect 17184 3420 17877 3448
rect 17184 3408 17190 3420
rect 17865 3417 17877 3420
rect 17911 3417 17923 3451
rect 17865 3411 17923 3417
rect 2314 3340 2320 3392
rect 2372 3380 2378 3392
rect 9490 3380 9496 3392
rect 2372 3352 9496 3380
rect 2372 3340 2378 3352
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 10870 3380 10876 3392
rect 9824 3352 10876 3380
rect 9824 3340 9830 3352
rect 10870 3340 10876 3352
rect 10928 3380 10934 3392
rect 11333 3383 11391 3389
rect 11333 3380 11345 3383
rect 10928 3352 11345 3380
rect 10928 3340 10934 3352
rect 11333 3349 11345 3352
rect 11379 3349 11391 3383
rect 11333 3343 11391 3349
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12802 3380 12808 3392
rect 11756 3352 12808 3380
rect 11756 3340 11762 3352
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 16022 3380 16028 3392
rect 13412 3352 16028 3380
rect 13412 3340 13418 3352
rect 16022 3340 16028 3352
rect 16080 3340 16086 3392
rect 16206 3380 16212 3392
rect 16167 3352 16212 3380
rect 16206 3340 16212 3352
rect 16264 3340 16270 3392
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 17310 3340 17316 3352
rect 17368 3380 17374 3392
rect 17972 3380 18000 3556
rect 18785 3553 18797 3556
rect 18831 3553 18843 3587
rect 19444 3584 19472 3692
rect 19797 3689 19809 3723
rect 19843 3720 19855 3723
rect 19886 3720 19892 3732
rect 19843 3692 19892 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 19521 3655 19579 3661
rect 19521 3621 19533 3655
rect 19567 3652 19579 3655
rect 19978 3652 19984 3664
rect 19567 3624 19984 3652
rect 19567 3621 19579 3624
rect 19521 3615 19579 3621
rect 19978 3612 19984 3624
rect 20036 3612 20042 3664
rect 19886 3584 19892 3596
rect 18785 3547 18843 3553
rect 18892 3556 19380 3584
rect 19444 3556 19892 3584
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18892 3516 18920 3556
rect 18380 3488 18920 3516
rect 19061 3519 19119 3525
rect 18380 3476 18386 3488
rect 19061 3485 19073 3519
rect 19107 3516 19119 3519
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 19107 3488 19257 3516
rect 19107 3485 19119 3488
rect 19061 3479 19119 3485
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19352 3516 19380 3556
rect 19886 3544 19892 3556
rect 19944 3544 19950 3596
rect 20162 3584 20168 3596
rect 20123 3556 20168 3584
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 20257 3587 20315 3593
rect 20257 3553 20269 3587
rect 20303 3584 20315 3587
rect 20901 3587 20959 3593
rect 20303 3556 20392 3584
rect 20303 3553 20315 3556
rect 20257 3547 20315 3553
rect 20180 3516 20208 3544
rect 19352 3488 20208 3516
rect 19245 3479 19303 3485
rect 20364 3448 20392 3556
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 21358 3584 21364 3596
rect 20947 3556 21364 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 20441 3519 20499 3525
rect 20441 3485 20453 3519
rect 20487 3516 20499 3519
rect 20625 3519 20683 3525
rect 20625 3516 20637 3519
rect 20487 3488 20637 3516
rect 20487 3485 20499 3488
rect 20441 3479 20499 3485
rect 20625 3485 20637 3488
rect 20671 3485 20683 3519
rect 20625 3479 20683 3485
rect 21174 3448 21180 3460
rect 20364 3420 21180 3448
rect 21174 3408 21180 3420
rect 21232 3408 21238 3460
rect 17368 3352 18000 3380
rect 18417 3383 18475 3389
rect 17368 3340 17374 3352
rect 18417 3349 18429 3383
rect 18463 3380 18475 3383
rect 18874 3380 18880 3392
rect 18463 3352 18880 3380
rect 18463 3349 18475 3352
rect 18417 3343 18475 3349
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 19245 3383 19303 3389
rect 19245 3349 19257 3383
rect 19291 3380 19303 3383
rect 20438 3380 20444 3392
rect 19291 3352 20444 3380
rect 19291 3349 19303 3352
rect 19245 3343 19303 3349
rect 20438 3340 20444 3352
rect 20496 3380 20502 3392
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 20496 3352 20637 3380
rect 20496 3340 20502 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 20625 3343 20683 3349
rect 20898 3340 20904 3392
rect 20956 3380 20962 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 20956 3352 21097 3380
rect 20956 3340 20962 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 8846 3176 8852 3188
rect 8807 3148 8852 3176
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9088 3148 10916 3176
rect 9088 3136 9094 3148
rect 8754 3068 8760 3120
rect 8812 3108 8818 3120
rect 9674 3108 9680 3120
rect 8812 3080 9680 3108
rect 8812 3068 8818 3080
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 10888 3108 10916 3148
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 11020 3148 11253 3176
rect 11020 3136 11026 3148
rect 11241 3145 11253 3148
rect 11287 3145 11299 3179
rect 11241 3139 11299 3145
rect 12529 3179 12587 3185
rect 12529 3145 12541 3179
rect 12575 3176 12587 3179
rect 12894 3176 12900 3188
rect 12575 3148 12900 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 15102 3176 15108 3188
rect 14516 3148 14688 3176
rect 15063 3148 15108 3176
rect 14516 3136 14522 3148
rect 13630 3108 13636 3120
rect 10888 3080 13636 3108
rect 13630 3068 13636 3080
rect 13688 3068 13694 3120
rect 14660 3108 14688 3148
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 18690 3176 18696 3188
rect 15212 3148 18696 3176
rect 15212 3108 15240 3148
rect 18690 3136 18696 3148
rect 18748 3136 18754 3188
rect 19150 3176 19156 3188
rect 18984 3148 19156 3176
rect 14660 3080 15240 3108
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 17589 3111 17647 3117
rect 17589 3108 17601 3111
rect 16632 3080 17601 3108
rect 16632 3068 16638 3080
rect 17589 3077 17601 3080
rect 17635 3077 17647 3111
rect 17589 3071 17647 3077
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 18049 3111 18107 3117
rect 18049 3108 18061 3111
rect 18012 3080 18061 3108
rect 18012 3068 18018 3080
rect 18049 3077 18061 3080
rect 18095 3077 18107 3111
rect 18049 3071 18107 3077
rect 18325 3111 18383 3117
rect 18325 3077 18337 3111
rect 18371 3108 18383 3111
rect 18417 3111 18475 3117
rect 18417 3108 18429 3111
rect 18371 3080 18429 3108
rect 18371 3077 18383 3080
rect 18325 3071 18383 3077
rect 18417 3077 18429 3080
rect 18463 3077 18475 3111
rect 18984 3108 19012 3148
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 19426 3176 19432 3188
rect 19387 3148 19432 3176
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 19610 3136 19616 3188
rect 19668 3176 19674 3188
rect 19668 3148 19932 3176
rect 19668 3136 19674 3148
rect 19794 3108 19800 3120
rect 18417 3071 18475 3077
rect 18708 3080 19012 3108
rect 19076 3080 19800 3108
rect 18708 3052 18736 3080
rect 7466 3040 7472 3052
rect 7427 3012 7472 3040
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 8628 3012 9137 3040
rect 8628 3000 8634 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 9490 3000 9496 3052
rect 9548 3040 9554 3052
rect 12618 3040 12624 3052
rect 9548 3012 9996 3040
rect 9548 3000 9554 3012
rect 7736 2975 7794 2981
rect 7736 2941 7748 2975
rect 7782 2972 7794 2975
rect 9674 2972 9680 2984
rect 7782 2944 9680 2972
rect 7782 2941 7794 2944
rect 7736 2935 7794 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9858 2972 9864 2984
rect 9819 2944 9864 2972
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 9968 2972 9996 3012
rect 11808 3012 12624 3040
rect 11514 2972 11520 2984
rect 9968 2944 11520 2972
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11808 2981 11836 3012
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 18690 3000 18696 3052
rect 18748 3000 18754 3052
rect 18874 3040 18880 3052
rect 18835 3012 18880 3040
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19076 3049 19104 3080
rect 19794 3068 19800 3080
rect 19852 3068 19858 3120
rect 19904 3108 19932 3148
rect 20717 3111 20775 3117
rect 20717 3108 20729 3111
rect 19904 3080 20729 3108
rect 20717 3077 20729 3080
rect 20763 3077 20775 3111
rect 20717 3071 20775 3077
rect 20993 3111 21051 3117
rect 20993 3077 21005 3111
rect 21039 3077 21051 3111
rect 20993 3071 21051 3077
rect 19061 3043 19119 3049
rect 19061 3009 19073 3043
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 19518 3000 19524 3052
rect 19576 3040 19582 3052
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19576 3012 19901 3040
rect 19576 3000 19582 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 21008 3040 21036 3071
rect 19981 3003 20039 3009
rect 20088 3012 21036 3040
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12032 2944 12909 2972
rect 12032 2932 12038 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 12897 2935 12955 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 15648 2975 15706 2981
rect 14424 2944 15240 2972
rect 14424 2932 14430 2944
rect 7834 2864 7840 2916
rect 7892 2904 7898 2916
rect 9950 2904 9956 2916
rect 7892 2876 9956 2904
rect 7892 2864 7898 2876
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 10128 2907 10186 2913
rect 10128 2873 10140 2907
rect 10174 2904 10186 2907
rect 13078 2904 13084 2916
rect 10174 2876 13084 2904
rect 10174 2873 10186 2876
rect 10128 2867 10186 2873
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 13992 2907 14050 2913
rect 13992 2873 14004 2907
rect 14038 2904 14050 2907
rect 14642 2904 14648 2916
rect 14038 2876 14648 2904
rect 14038 2873 14050 2876
rect 13992 2867 14050 2873
rect 14642 2864 14648 2876
rect 14700 2904 14706 2916
rect 15212 2904 15240 2944
rect 15648 2941 15660 2975
rect 15694 2972 15706 2975
rect 16850 2972 16856 2984
rect 15694 2944 16856 2972
rect 15694 2941 15706 2944
rect 15648 2935 15706 2941
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 17175 2944 17417 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 17405 2941 17417 2944
rect 17451 2972 17463 2975
rect 17678 2972 17684 2984
rect 17451 2944 17684 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 17678 2932 17684 2944
rect 17736 2932 17742 2984
rect 18046 2932 18052 2984
rect 18104 2972 18110 2984
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 18104 2944 18797 2972
rect 18104 2932 18110 2944
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 18966 2932 18972 2984
rect 19024 2972 19030 2984
rect 19996 2972 20024 3003
rect 19024 2944 20024 2972
rect 19024 2932 19030 2944
rect 18325 2907 18383 2913
rect 14700 2876 15148 2904
rect 15212 2876 18184 2904
rect 14700 2864 14706 2876
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 11606 2836 11612 2848
rect 5684 2808 11612 2836
rect 5684 2796 5690 2808
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11698 2796 11704 2848
rect 11756 2836 11762 2848
rect 11977 2839 12035 2845
rect 11977 2836 11989 2839
rect 11756 2808 11989 2836
rect 11756 2796 11762 2808
rect 11977 2805 11989 2808
rect 12023 2805 12035 2839
rect 15120 2836 15148 2876
rect 16761 2839 16819 2845
rect 16761 2836 16773 2839
rect 15120 2808 16773 2836
rect 11977 2799 12035 2805
rect 16761 2805 16773 2808
rect 16807 2805 16819 2839
rect 18156 2836 18184 2876
rect 18325 2873 18337 2907
rect 18371 2904 18383 2907
rect 19797 2907 19855 2913
rect 19797 2904 19809 2907
rect 18371 2876 19809 2904
rect 18371 2873 18383 2876
rect 18325 2867 18383 2873
rect 19797 2873 19809 2876
rect 19843 2873 19855 2907
rect 19797 2867 19855 2873
rect 20088 2836 20116 3012
rect 20717 2975 20775 2981
rect 20717 2941 20729 2975
rect 20763 2972 20775 2975
rect 20809 2975 20867 2981
rect 20809 2972 20821 2975
rect 20763 2944 20821 2972
rect 20763 2941 20775 2944
rect 20717 2935 20775 2941
rect 20809 2941 20821 2944
rect 20855 2941 20867 2975
rect 20809 2935 20867 2941
rect 20530 2864 20536 2916
rect 20588 2904 20594 2916
rect 21818 2904 21824 2916
rect 20588 2876 21824 2904
rect 20588 2864 20594 2876
rect 21818 2864 21824 2876
rect 21876 2864 21882 2916
rect 18156 2808 20116 2836
rect 20441 2839 20499 2845
rect 16761 2799 16819 2805
rect 20441 2805 20453 2839
rect 20487 2836 20499 2839
rect 20898 2836 20904 2848
rect 20487 2808 20904 2836
rect 20487 2805 20499 2808
rect 20441 2799 20499 2805
rect 20898 2796 20904 2808
rect 20956 2836 20962 2848
rect 21726 2836 21732 2848
rect 20956 2808 21732 2836
rect 20956 2796 20962 2808
rect 21726 2796 21732 2808
rect 21784 2796 21790 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8662 2632 8668 2644
rect 7975 2604 8668 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 10008 2604 10149 2632
rect 10008 2592 10014 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10137 2595 10195 2601
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 10686 2632 10692 2644
rect 10551 2604 10692 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 10152 2564 10180 2595
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 11296 2604 11529 2632
rect 11296 2592 11302 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 12161 2635 12219 2641
rect 12161 2601 12173 2635
rect 12207 2632 12219 2635
rect 12710 2632 12716 2644
rect 12207 2604 12716 2632
rect 12207 2601 12219 2604
rect 12161 2595 12219 2601
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 13078 2592 13084 2644
rect 13136 2632 13142 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 13136 2604 14013 2632
rect 13136 2592 13142 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 14001 2595 14059 2601
rect 14369 2635 14427 2641
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 14550 2632 14556 2644
rect 14415 2604 14556 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14734 2632 14740 2644
rect 14695 2604 14740 2632
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 15344 2604 15485 2632
rect 15344 2592 15350 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 15933 2635 15991 2641
rect 15933 2601 15945 2635
rect 15979 2632 15991 2635
rect 16206 2632 16212 2644
rect 15979 2604 16212 2632
rect 15979 2601 15991 2604
rect 15933 2595 15991 2601
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 16485 2635 16543 2641
rect 16485 2601 16497 2635
rect 16531 2601 16543 2635
rect 16485 2595 16543 2601
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17034 2632 17040 2644
rect 16991 2604 17040 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 10873 2567 10931 2573
rect 10873 2564 10885 2567
rect 10152 2536 10885 2564
rect 10873 2533 10885 2536
rect 10919 2533 10931 2567
rect 10873 2527 10931 2533
rect 10962 2524 10968 2576
rect 11020 2524 11026 2576
rect 12888 2567 12946 2573
rect 12888 2533 12900 2567
rect 12934 2564 12946 2567
rect 13170 2564 13176 2576
rect 12934 2536 13176 2564
rect 12934 2533 12946 2536
rect 12888 2527 12946 2533
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 14829 2567 14887 2573
rect 14829 2564 14841 2567
rect 13688 2536 14841 2564
rect 13688 2524 13694 2536
rect 14829 2533 14841 2536
rect 14875 2533 14887 2567
rect 14829 2527 14887 2533
rect 15841 2567 15899 2573
rect 15841 2533 15853 2567
rect 15887 2564 15899 2567
rect 16500 2564 16528 2595
rect 17034 2592 17040 2604
rect 17092 2632 17098 2644
rect 18046 2632 18052 2644
rect 17092 2604 18052 2632
rect 17092 2592 17098 2604
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18417 2635 18475 2641
rect 18417 2601 18429 2635
rect 18463 2632 18475 2635
rect 19242 2632 19248 2644
rect 18463 2604 19248 2632
rect 18463 2601 18475 2604
rect 18417 2595 18475 2601
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 15887 2536 16528 2564
rect 16592 2536 16865 2564
rect 15887 2533 15899 2536
rect 15841 2527 15899 2533
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 7576 2468 8309 2496
rect 7282 2252 7288 2304
rect 7340 2292 7346 2304
rect 7576 2301 7604 2468
rect 8297 2465 8309 2468
rect 8343 2465 8355 2499
rect 8297 2459 8355 2465
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 8478 2496 8484 2508
rect 8435 2468 8484 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 8478 2456 8484 2468
rect 8536 2496 8542 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8536 2468 8953 2496
rect 8536 2456 8542 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 10980 2496 11008 2524
rect 11977 2499 12035 2505
rect 10980 2468 11100 2496
rect 8941 2459 8999 2465
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8846 2428 8852 2440
rect 8619 2400 8852 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 10962 2428 10968 2440
rect 9907 2400 10968 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11072 2437 11100 2468
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 12066 2496 12072 2508
rect 12023 2468 12072 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12492 2468 12633 2496
rect 12492 2456 12498 2468
rect 12621 2465 12633 2468
rect 12667 2496 12679 2499
rect 13722 2496 13728 2508
rect 12667 2468 13728 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 16592 2496 16620 2536
rect 16853 2533 16865 2536
rect 16899 2564 16911 2567
rect 17954 2564 17960 2576
rect 16899 2536 17960 2564
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 17954 2524 17960 2536
rect 18012 2524 18018 2576
rect 14568 2468 16620 2496
rect 17681 2499 17739 2505
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 9401 2363 9459 2369
rect 9401 2329 9413 2363
rect 9447 2360 9459 2363
rect 11790 2360 11796 2372
rect 9447 2332 11796 2360
rect 9447 2329 9459 2332
rect 9401 2323 9459 2329
rect 11790 2320 11796 2332
rect 11848 2320 11854 2372
rect 7561 2295 7619 2301
rect 7561 2292 7573 2295
rect 7340 2264 7573 2292
rect 7340 2252 7346 2264
rect 7561 2261 7573 2264
rect 7607 2261 7619 2295
rect 11808 2292 11836 2320
rect 14568 2292 14596 2468
rect 17681 2465 17693 2499
rect 17727 2496 17739 2499
rect 18432 2496 18460 2595
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 19610 2632 19616 2644
rect 19571 2604 19616 2632
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 21269 2635 21327 2641
rect 21269 2632 21281 2635
rect 20180 2604 21281 2632
rect 18598 2524 18604 2576
rect 18656 2564 18662 2576
rect 19061 2567 19119 2573
rect 19061 2564 19073 2567
rect 18656 2536 19073 2564
rect 18656 2524 18662 2536
rect 19061 2533 19073 2536
rect 19107 2533 19119 2567
rect 20070 2564 20076 2576
rect 19061 2527 19119 2533
rect 19904 2536 20076 2564
rect 17727 2468 18460 2496
rect 18785 2499 18843 2505
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 18785 2465 18797 2499
rect 18831 2496 18843 2499
rect 19904 2496 19932 2536
rect 20070 2524 20076 2536
rect 20128 2524 20134 2576
rect 18831 2468 19932 2496
rect 19981 2499 20039 2505
rect 18831 2465 18843 2468
rect 18785 2459 18843 2465
rect 19981 2465 19993 2499
rect 20027 2496 20039 2499
rect 20180 2496 20208 2604
rect 21269 2601 21281 2604
rect 21315 2632 21327 2635
rect 21818 2632 21824 2644
rect 21315 2604 21824 2632
rect 21315 2601 21327 2604
rect 21269 2595 21327 2601
rect 21818 2592 21824 2604
rect 21876 2592 21882 2644
rect 20027 2468 20208 2496
rect 20533 2499 20591 2505
rect 20027 2465 20039 2468
rect 19981 2459 20039 2465
rect 20533 2465 20545 2499
rect 20579 2496 20591 2499
rect 20898 2496 20904 2508
rect 20579 2468 20904 2496
rect 20579 2465 20591 2468
rect 20533 2459 20591 2465
rect 20898 2456 20904 2468
rect 20956 2456 20962 2508
rect 14642 2388 14648 2440
rect 14700 2428 14706 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14700 2400 15025 2428
rect 14700 2388 14706 2400
rect 15013 2397 15025 2400
rect 15059 2428 15071 2431
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15059 2400 16037 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 16850 2320 16856 2372
rect 16908 2360 16914 2372
rect 17052 2360 17080 2391
rect 17218 2388 17224 2440
rect 17276 2428 17282 2440
rect 17276 2400 20760 2428
rect 17276 2388 17282 2400
rect 20732 2369 20760 2400
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 16908 2332 17080 2360
rect 17144 2332 20177 2360
rect 16908 2320 16914 2332
rect 11808 2264 14596 2292
rect 7561 2255 7619 2261
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 17144 2292 17172 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 20165 2323 20223 2329
rect 20717 2363 20775 2369
rect 20717 2329 20729 2363
rect 20763 2329 20775 2363
rect 20717 2323 20775 2329
rect 16080 2264 17172 2292
rect 16080 2252 16086 2264
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 17736 2264 17877 2292
rect 17736 2252 17742 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 16390 2088 16396 2100
rect 11204 2060 16396 2088
rect 11204 2048 11210 2060
rect 16390 2048 16396 2060
rect 16448 2048 16454 2100
rect 1762 1368 1768 1420
rect 1820 1408 1826 1420
rect 8754 1408 8760 1420
rect 1820 1380 8760 1408
rect 1820 1368 1826 1380
rect 8754 1368 8760 1380
rect 8812 1368 8818 1420
rect 15470 1368 15476 1420
rect 15528 1408 15534 1420
rect 17218 1408 17224 1420
rect 15528 1380 17224 1408
rect 15528 1368 15534 1380
rect 17218 1368 17224 1380
rect 17276 1368 17282 1420
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 20444 20043 20496 20052
rect 20444 20009 20453 20043
rect 20453 20009 20487 20043
rect 20487 20009 20496 20043
rect 20444 20000 20496 20009
rect 21088 20043 21140 20052
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 20260 19907 20312 19916
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 20812 19864 20864 19916
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 20996 19499 21048 19508
rect 20996 19465 21005 19499
rect 21005 19465 21039 19499
rect 21039 19465 21048 19499
rect 20996 19456 21048 19465
rect 5724 19252 5776 19304
rect 18512 19252 18564 19304
rect 20168 19252 20220 19304
rect 20352 19252 20404 19304
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 19248 19116 19300 19168
rect 20536 19116 20588 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 20260 18912 20312 18964
rect 21088 18955 21140 18964
rect 21088 18921 21097 18955
rect 21097 18921 21131 18955
rect 21131 18921 21140 18955
rect 21088 18912 21140 18921
rect 11704 18776 11756 18828
rect 15844 18819 15896 18828
rect 15844 18785 15853 18819
rect 15853 18785 15887 18819
rect 15887 18785 15896 18819
rect 15844 18776 15896 18785
rect 18512 18887 18564 18896
rect 16856 18776 16908 18828
rect 18512 18853 18521 18887
rect 18521 18853 18555 18887
rect 18555 18853 18564 18887
rect 18512 18844 18564 18853
rect 20168 18887 20220 18896
rect 19892 18819 19944 18828
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 20168 18853 20177 18887
rect 20177 18853 20211 18887
rect 20211 18853 20220 18887
rect 20168 18844 20220 18853
rect 20812 18844 20864 18896
rect 20720 18776 20772 18828
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 20352 18300 20404 18352
rect 8852 18164 8904 18216
rect 20812 18207 20864 18216
rect 20812 18173 20821 18207
rect 20821 18173 20855 18207
rect 20855 18173 20864 18207
rect 20812 18164 20864 18173
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 21088 17867 21140 17876
rect 21088 17833 21097 17867
rect 21097 17833 21131 17867
rect 21131 17833 21140 17867
rect 21088 17824 21140 17833
rect 8392 17688 8444 17740
rect 20168 17688 20220 17740
rect 20720 17620 20772 17672
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 18788 17323 18840 17332
rect 18788 17289 18797 17323
rect 18797 17289 18831 17323
rect 18831 17289 18840 17323
rect 18788 17280 18840 17289
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 20168 17187 20220 17196
rect 11244 17119 11296 17128
rect 11244 17085 11253 17119
rect 11253 17085 11287 17119
rect 11287 17085 11296 17119
rect 11244 17076 11296 17085
rect 17960 17076 18012 17128
rect 13084 17008 13136 17060
rect 20168 17153 20177 17187
rect 20177 17153 20211 17187
rect 20211 17153 20220 17187
rect 20168 17144 20220 17153
rect 20260 17076 20312 17128
rect 20720 17008 20772 17060
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 21088 16779 21140 16788
rect 21088 16745 21097 16779
rect 21097 16745 21131 16779
rect 21131 16745 21140 16779
rect 21088 16736 21140 16745
rect 17960 16711 18012 16720
rect 17960 16677 17969 16711
rect 17969 16677 18003 16711
rect 18003 16677 18012 16711
rect 17960 16668 18012 16677
rect 18052 16668 18104 16720
rect 18788 16600 18840 16652
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 20996 16235 21048 16244
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 20260 16056 20312 16108
rect 19800 15988 19852 16040
rect 20812 16031 20864 16040
rect 20812 15997 20821 16031
rect 20821 15997 20855 16031
rect 20855 15997 20864 16031
rect 20812 15988 20864 15997
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 18052 15580 18104 15632
rect 14004 15512 14056 15564
rect 15200 15512 15252 15564
rect 20720 15512 20772 15564
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 20996 15147 21048 15156
rect 20996 15113 21005 15147
rect 21005 15113 21039 15147
rect 21039 15113 21048 15147
rect 20996 15104 21048 15113
rect 15200 14968 15252 15020
rect 11060 14900 11112 14952
rect 18696 14900 18748 14952
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 20628 14560 20680 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 20812 14492 20864 14544
rect 8576 14424 8628 14476
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 18788 14424 18840 14476
rect 20720 14356 20772 14408
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 20720 13923 20772 13932
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 20720 13880 20772 13889
rect 10968 13812 11020 13864
rect 18696 13812 18748 13864
rect 20628 13812 20680 13864
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 17868 13472 17920 13524
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 21088 13515 21140 13524
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 16580 13404 16632 13456
rect 12992 13336 13044 13388
rect 18788 13336 18840 13388
rect 20536 13336 20588 13388
rect 19984 13268 20036 13320
rect 16488 13132 16540 13184
rect 20260 13132 20312 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 14280 12792 14332 12844
rect 20536 12835 20588 12844
rect 19524 12724 19576 12776
rect 19984 12724 20036 12776
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 20444 12724 20496 12776
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 20628 12588 20680 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 15844 12384 15896 12436
rect 16856 12427 16908 12436
rect 16856 12393 16865 12427
rect 16865 12393 16899 12427
rect 16899 12393 16908 12427
rect 16856 12384 16908 12393
rect 18052 12384 18104 12436
rect 21088 12427 21140 12436
rect 21088 12393 21097 12427
rect 21097 12393 21131 12427
rect 21131 12393 21140 12427
rect 21088 12384 21140 12393
rect 13176 12316 13228 12368
rect 20168 12316 20220 12368
rect 20444 12316 20496 12368
rect 15016 12248 15068 12300
rect 18144 12291 18196 12300
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 18144 12257 18178 12291
rect 18178 12257 18196 12291
rect 18144 12248 18196 12257
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 19156 12180 19208 12232
rect 13360 12044 13412 12096
rect 19892 12112 19944 12164
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 12256 11840 12308 11892
rect 17408 11840 17460 11892
rect 10968 11704 11020 11756
rect 11796 11704 11848 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 20904 11840 20956 11892
rect 15292 11636 15344 11688
rect 16764 11636 16816 11688
rect 17868 11636 17920 11688
rect 15936 11568 15988 11620
rect 16672 11568 16724 11620
rect 19248 11568 19300 11620
rect 20352 11568 20404 11620
rect 20628 11636 20680 11688
rect 20904 11568 20956 11620
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 19340 11500 19392 11552
rect 19432 11500 19484 11552
rect 22100 11500 22152 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 4068 11296 4120 11348
rect 13176 11296 13228 11348
rect 13360 11339 13412 11348
rect 13360 11305 13369 11339
rect 13369 11305 13403 11339
rect 13403 11305 13412 11339
rect 13360 11296 13412 11305
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 18144 11296 18196 11348
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 19156 11339 19208 11348
rect 19156 11305 19165 11339
rect 19165 11305 19199 11339
rect 19199 11305 19208 11339
rect 19156 11296 19208 11305
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 16856 11228 16908 11280
rect 17408 11228 17460 11280
rect 12164 11203 12216 11212
rect 12164 11169 12196 11203
rect 12196 11169 12216 11203
rect 12164 11160 12216 11169
rect 15568 11203 15620 11212
rect 15568 11169 15602 11203
rect 15602 11169 15620 11203
rect 15568 11160 15620 11169
rect 19340 11160 19392 11212
rect 19892 11160 19944 11212
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 12624 11092 12676 11144
rect 13820 11135 13872 11144
rect 13820 11101 13829 11135
rect 13829 11101 13863 11135
rect 13863 11101 13872 11135
rect 13820 11092 13872 11101
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 15292 11135 15344 11144
rect 13912 11092 13964 11101
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20352 11135 20404 11144
rect 20352 11101 20361 11135
rect 20361 11101 20395 11135
rect 20395 11101 20404 11135
rect 20352 11092 20404 11101
rect 14188 10956 14240 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 13912 10795 13964 10804
rect 13912 10761 13921 10795
rect 13921 10761 13955 10795
rect 13955 10761 13964 10795
rect 13912 10752 13964 10761
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 15752 10752 15804 10804
rect 17316 10752 17368 10804
rect 12440 10548 12492 10600
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 16856 10616 16908 10668
rect 19432 10616 19484 10668
rect 16948 10548 17000 10600
rect 17868 10548 17920 10600
rect 13912 10480 13964 10532
rect 15752 10480 15804 10532
rect 18328 10523 18380 10532
rect 18328 10489 18362 10523
rect 18362 10489 18380 10523
rect 18328 10480 18380 10489
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 17224 10455 17276 10464
rect 17224 10421 17233 10455
rect 17233 10421 17267 10455
rect 17267 10421 17276 10455
rect 17224 10412 17276 10421
rect 18052 10412 18104 10464
rect 19432 10455 19484 10464
rect 19432 10421 19441 10455
rect 19441 10421 19475 10455
rect 19475 10421 19484 10455
rect 19432 10412 19484 10421
rect 21088 10455 21140 10464
rect 21088 10421 21097 10455
rect 21097 10421 21131 10455
rect 21131 10421 21140 10455
rect 21088 10412 21140 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 20260 10251 20312 10260
rect 20260 10217 20269 10251
rect 20269 10217 20303 10251
rect 20303 10217 20312 10251
rect 20260 10208 20312 10217
rect 9588 10140 9640 10192
rect 16212 10140 16264 10192
rect 16580 10115 16632 10124
rect 16580 10081 16589 10115
rect 16589 10081 16623 10115
rect 16623 10081 16632 10115
rect 16580 10072 16632 10081
rect 12164 10004 12216 10056
rect 16948 10072 17000 10124
rect 18052 10072 18104 10124
rect 18144 10072 18196 10124
rect 19892 10072 19944 10124
rect 21088 10140 21140 10192
rect 20904 10115 20956 10124
rect 13360 9936 13412 9988
rect 14188 9936 14240 9988
rect 18328 10004 18380 10056
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 664 9868 716 9920
rect 9588 9868 9640 9920
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 15752 9868 15804 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 13636 9460 13688 9512
rect 14188 9664 14240 9716
rect 17868 9596 17920 9648
rect 16672 9528 16724 9580
rect 18144 9528 18196 9580
rect 15752 9460 15804 9512
rect 18420 9460 18472 9512
rect 19432 9460 19484 9512
rect 10508 9392 10560 9444
rect 14740 9392 14792 9444
rect 10968 9324 11020 9376
rect 11244 9324 11296 9376
rect 13268 9324 13320 9376
rect 15384 9324 15436 9376
rect 19800 9392 19852 9444
rect 20628 9392 20680 9444
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 16396 9324 16448 9376
rect 17224 9324 17276 9376
rect 19708 9367 19760 9376
rect 19708 9333 19717 9367
rect 19717 9333 19751 9367
rect 19751 9333 19760 9367
rect 19708 9324 19760 9333
rect 19984 9324 20036 9376
rect 20168 9324 20220 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 9680 9120 9732 9172
rect 11612 9163 11664 9172
rect 11612 9129 11621 9163
rect 11621 9129 11655 9163
rect 11655 9129 11664 9163
rect 11612 9120 11664 9129
rect 10048 8984 10100 9036
rect 10968 8984 11020 9036
rect 14740 9120 14792 9172
rect 16120 9120 16172 9172
rect 20536 9120 20588 9172
rect 13544 9052 13596 9104
rect 19432 9052 19484 9104
rect 12440 8984 12492 9036
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 9496 8916 9548 8968
rect 13636 8984 13688 9036
rect 15384 8984 15436 9036
rect 15844 8984 15896 9036
rect 16120 8984 16172 9036
rect 16856 8984 16908 9036
rect 18972 8984 19024 9036
rect 19892 8984 19944 9036
rect 18788 8916 18840 8968
rect 19708 8916 19760 8968
rect 10416 8780 10468 8832
rect 11796 8780 11848 8832
rect 14188 8780 14240 8832
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 16856 8780 16908 8832
rect 17960 8780 18012 8832
rect 20720 8848 20772 8900
rect 19892 8780 19944 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 10968 8576 11020 8628
rect 11796 8576 11848 8628
rect 16120 8576 16172 8628
rect 16580 8576 16632 8628
rect 17500 8576 17552 8628
rect 20628 8576 20680 8628
rect 20904 8576 20956 8628
rect 13636 8508 13688 8560
rect 11244 8440 11296 8492
rect 9220 8304 9272 8356
rect 14372 8372 14424 8424
rect 14188 8304 14240 8356
rect 18604 8508 18656 8560
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 16672 8372 16724 8424
rect 10048 8236 10100 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 16028 8304 16080 8356
rect 19708 8415 19760 8424
rect 19708 8381 19742 8415
rect 19742 8381 19760 8415
rect 19708 8372 19760 8381
rect 18512 8304 18564 8356
rect 17224 8279 17276 8288
rect 17224 8245 17233 8279
rect 17233 8245 17267 8279
rect 17267 8245 17276 8279
rect 17224 8236 17276 8245
rect 18604 8279 18656 8288
rect 18604 8245 18613 8279
rect 18613 8245 18647 8279
rect 18647 8245 18656 8279
rect 18604 8236 18656 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 10508 8075 10560 8084
rect 10508 8041 10517 8075
rect 10517 8041 10551 8075
rect 10551 8041 10560 8075
rect 10508 8032 10560 8041
rect 11704 8032 11756 8084
rect 14004 8075 14056 8084
rect 14004 8041 14013 8075
rect 14013 8041 14047 8075
rect 14047 8041 14056 8075
rect 14004 8032 14056 8041
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 16212 8032 16264 8084
rect 18512 8032 18564 8084
rect 20260 8032 20312 8084
rect 10968 7964 11020 8016
rect 11704 7896 11756 7948
rect 12808 7896 12860 7948
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12532 7828 12584 7880
rect 13268 7828 13320 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 11244 7760 11296 7812
rect 11796 7760 11848 7812
rect 14740 7828 14792 7880
rect 8944 7692 8996 7744
rect 12072 7692 12124 7744
rect 12348 7692 12400 7744
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 17224 7896 17276 7948
rect 19892 7896 19944 7948
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 16028 7828 16080 7880
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 18880 7760 18932 7812
rect 17868 7692 17920 7744
rect 19708 7828 19760 7880
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 20628 7828 20680 7880
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 8852 7531 8904 7540
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 11980 7488 12032 7540
rect 13820 7488 13872 7540
rect 16764 7488 16816 7540
rect 18696 7488 18748 7540
rect 20076 7488 20128 7540
rect 20260 7420 20312 7472
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13912 7352 13964 7404
rect 16672 7352 16724 7404
rect 17224 7352 17276 7404
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 20168 7352 20220 7404
rect 11244 7284 11296 7336
rect 11336 7284 11388 7336
rect 12532 7284 12584 7336
rect 17960 7284 18012 7336
rect 19708 7327 19760 7336
rect 19708 7293 19717 7327
rect 19717 7293 19751 7327
rect 19751 7293 19760 7327
rect 19708 7284 19760 7293
rect 14464 7259 14516 7268
rect 14464 7225 14473 7259
rect 14473 7225 14507 7259
rect 14507 7225 14516 7259
rect 14464 7216 14516 7225
rect 14648 7216 14700 7268
rect 19524 7216 19576 7268
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 10876 7148 10928 7200
rect 13912 7148 13964 7200
rect 14556 7191 14608 7200
rect 14556 7157 14565 7191
rect 14565 7157 14599 7191
rect 14599 7157 14608 7191
rect 14556 7148 14608 7157
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 17224 7191 17276 7200
rect 16304 7148 16356 7157
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 18144 7148 18196 7200
rect 18880 7148 18932 7200
rect 19156 7148 19208 7200
rect 20076 7148 20128 7200
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 9404 6944 9456 6996
rect 11152 6944 11204 6996
rect 12532 6944 12584 6996
rect 16672 6987 16724 6996
rect 16672 6953 16681 6987
rect 16681 6953 16715 6987
rect 16715 6953 16724 6987
rect 16672 6944 16724 6953
rect 19984 6944 20036 6996
rect 8760 6808 8812 6860
rect 12440 6808 12492 6860
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 13268 6604 13320 6656
rect 14556 6604 14608 6656
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 16028 6808 16080 6860
rect 16580 6808 16632 6860
rect 19156 6876 19208 6928
rect 17592 6808 17644 6860
rect 19064 6851 19116 6860
rect 19064 6817 19098 6851
rect 19098 6817 19116 6851
rect 19064 6808 19116 6817
rect 16948 6783 17000 6792
rect 16948 6749 16957 6783
rect 16957 6749 16991 6783
rect 16991 6749 17000 6783
rect 16948 6740 17000 6749
rect 20168 6715 20220 6724
rect 20168 6681 20177 6715
rect 20177 6681 20211 6715
rect 20211 6681 20220 6715
rect 20168 6672 20220 6681
rect 17868 6604 17920 6656
rect 18144 6604 18196 6656
rect 20628 6604 20680 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 8760 6400 8812 6452
rect 9312 6400 9364 6452
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 13084 6443 13136 6452
rect 13084 6409 13093 6443
rect 13093 6409 13127 6443
rect 13127 6409 13136 6443
rect 13084 6400 13136 6409
rect 16028 6443 16080 6452
rect 16028 6409 16037 6443
rect 16037 6409 16071 6443
rect 16071 6409 16080 6443
rect 16028 6400 16080 6409
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 16028 6264 16080 6316
rect 8208 6196 8260 6248
rect 13636 6196 13688 6248
rect 8300 6128 8352 6180
rect 9496 6171 9548 6180
rect 9496 6137 9505 6171
rect 9505 6137 9539 6171
rect 9539 6137 9548 6171
rect 9496 6128 9548 6137
rect 10692 6128 10744 6180
rect 13912 6128 13964 6180
rect 14464 6128 14516 6180
rect 16488 6196 16540 6248
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 17500 6239 17552 6248
rect 17500 6205 17509 6239
rect 17509 6205 17543 6239
rect 17543 6205 17552 6239
rect 17500 6196 17552 6205
rect 19064 6400 19116 6452
rect 18144 6196 18196 6248
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 9680 6060 9732 6112
rect 10876 6060 10928 6112
rect 11244 6060 11296 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 11796 6060 11848 6112
rect 12072 6060 12124 6112
rect 12716 6060 12768 6112
rect 14004 6060 14056 6112
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 16948 6060 17000 6112
rect 17592 6060 17644 6112
rect 20168 6128 20220 6180
rect 20352 6060 20404 6112
rect 20444 6060 20496 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 8392 5856 8444 5908
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 14372 5856 14424 5908
rect 16212 5856 16264 5908
rect 16672 5856 16724 5908
rect 7564 5720 7616 5772
rect 9956 5788 10008 5840
rect 10048 5720 10100 5772
rect 11152 5720 11204 5772
rect 13360 5788 13412 5840
rect 12440 5720 12492 5772
rect 14096 5720 14148 5772
rect 7196 5652 7248 5704
rect 8300 5652 8352 5704
rect 15752 5788 15804 5840
rect 17868 5856 17920 5908
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 14740 5652 14792 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 9128 5559 9180 5568
rect 9128 5525 9137 5559
rect 9137 5525 9171 5559
rect 9171 5525 9180 5559
rect 9128 5516 9180 5525
rect 9496 5516 9548 5568
rect 11060 5516 11112 5568
rect 12072 5559 12124 5568
rect 12072 5525 12081 5559
rect 12081 5525 12115 5559
rect 12115 5525 12124 5559
rect 13728 5559 13780 5568
rect 12072 5516 12124 5525
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 15476 5584 15528 5636
rect 17776 5788 17828 5840
rect 18696 5720 18748 5772
rect 19984 5720 20036 5772
rect 20904 5763 20956 5772
rect 16028 5652 16080 5704
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 16488 5584 16540 5636
rect 18972 5652 19024 5704
rect 19064 5652 19116 5704
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 20352 5652 20404 5661
rect 21640 5652 21692 5704
rect 19524 5584 19576 5636
rect 21548 5584 21600 5636
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 22008 5559 22060 5568
rect 22008 5525 22017 5559
rect 22017 5525 22051 5559
rect 22051 5525 22060 5559
rect 22008 5516 22060 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 8300 5312 8352 5364
rect 9036 5312 9088 5364
rect 11152 5312 11204 5364
rect 15752 5312 15804 5364
rect 16764 5312 16816 5364
rect 16856 5312 16908 5364
rect 19156 5312 19208 5364
rect 19984 5355 20036 5364
rect 19984 5321 19993 5355
rect 19993 5321 20027 5355
rect 20027 5321 20036 5355
rect 19984 5312 20036 5321
rect 9220 5176 9272 5228
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 11244 5176 11296 5228
rect 17960 5244 18012 5296
rect 20812 5244 20864 5296
rect 15660 5176 15712 5228
rect 16488 5176 16540 5228
rect 19064 5176 19116 5228
rect 20352 5176 20404 5228
rect 8208 5108 8260 5160
rect 7748 5040 7800 5092
rect 11060 5108 11112 5160
rect 12440 5108 12492 5160
rect 13728 5108 13780 5160
rect 14372 5108 14424 5160
rect 17132 5108 17184 5160
rect 18604 5108 18656 5160
rect 18972 5108 19024 5160
rect 20996 5151 21048 5160
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 16028 5040 16080 5092
rect 21456 5040 21508 5092
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 9588 4972 9640 5024
rect 11244 4972 11296 5024
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 14464 4972 14516 5024
rect 15476 4972 15528 5024
rect 16488 4972 16540 5024
rect 18144 4972 18196 5024
rect 18880 4972 18932 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 8576 4768 8628 4820
rect 10692 4768 10744 4820
rect 12716 4811 12768 4820
rect 12716 4777 12725 4811
rect 12725 4777 12759 4811
rect 12759 4777 12768 4811
rect 12716 4768 12768 4777
rect 14188 4768 14240 4820
rect 16856 4768 16908 4820
rect 20996 4768 21048 4820
rect 5356 4700 5408 4752
rect 8576 4675 8628 4684
rect 5448 4428 5500 4480
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 9588 4700 9640 4752
rect 11704 4700 11756 4752
rect 16580 4700 16632 4752
rect 19800 4700 19852 4752
rect 11980 4632 12032 4684
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 8668 4607 8720 4616
rect 7748 4564 7800 4573
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 8852 4607 8904 4616
rect 8852 4573 8861 4607
rect 8861 4573 8895 4607
rect 8895 4573 8904 4607
rect 8852 4564 8904 4573
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 8760 4496 8812 4548
rect 8484 4428 8536 4480
rect 11244 4428 11296 4480
rect 12440 4496 12492 4548
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 16488 4632 16540 4684
rect 19064 4632 19116 4684
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 14556 4564 14608 4616
rect 17040 4564 17092 4616
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 21272 4632 21324 4684
rect 12716 4496 12768 4548
rect 13636 4428 13688 4480
rect 14464 4428 14516 4480
rect 16028 4496 16080 4548
rect 19340 4496 19392 4548
rect 16672 4428 16724 4480
rect 17040 4428 17092 4480
rect 18788 4428 18840 4480
rect 18972 4471 19024 4480
rect 18972 4437 18981 4471
rect 18981 4437 19015 4471
rect 19015 4437 19024 4471
rect 18972 4428 19024 4437
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19524 4428 19576 4437
rect 20168 4428 20220 4480
rect 21180 4428 21232 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 8944 4224 8996 4276
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 10416 4267 10468 4276
rect 10416 4233 10425 4267
rect 10425 4233 10459 4267
rect 10459 4233 10468 4267
rect 10416 4224 10468 4233
rect 11152 4224 11204 4276
rect 11244 4224 11296 4276
rect 16212 4224 16264 4276
rect 18880 4224 18932 4276
rect 11060 4156 11112 4208
rect 12716 4156 12768 4208
rect 10968 4131 11020 4140
rect 3424 4020 3476 4072
rect 5356 4020 5408 4072
rect 6184 4020 6236 4072
rect 7932 4020 7984 4072
rect 8392 4020 8444 4072
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 14372 4156 14424 4208
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 17960 4156 18012 4208
rect 18328 4156 18380 4208
rect 19800 4224 19852 4276
rect 19984 4224 20036 4276
rect 21640 4156 21692 4208
rect 14096 4088 14148 4097
rect 17132 4088 17184 4140
rect 18236 4088 18288 4140
rect 20444 4088 20496 4140
rect 21364 4131 21416 4140
rect 21364 4097 21373 4131
rect 21373 4097 21407 4131
rect 21407 4097 21416 4131
rect 21364 4088 21416 4097
rect 10692 4020 10744 4072
rect 10876 4063 10928 4072
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 2872 3952 2924 4004
rect 5448 3952 5500 4004
rect 8852 3952 8904 4004
rect 11244 4020 11296 4072
rect 12992 4020 13044 4072
rect 14372 4020 14424 4072
rect 14648 4020 14700 4072
rect 14740 4020 14792 4072
rect 15384 4020 15436 4072
rect 17592 4020 17644 4072
rect 13360 3952 13412 4004
rect 5080 3884 5132 3936
rect 12348 3884 12400 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 15476 3884 15528 3936
rect 17132 3884 17184 3936
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 17592 3927 17644 3936
rect 17592 3893 17601 3927
rect 17601 3893 17635 3927
rect 17635 3893 17644 3927
rect 17592 3884 17644 3893
rect 17776 3884 17828 3936
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 18880 3952 18932 4004
rect 20168 3952 20220 4004
rect 18972 3884 19024 3936
rect 19064 3884 19116 3936
rect 20812 4020 20864 4072
rect 20904 3884 20956 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 3976 3680 4028 3732
rect 8760 3680 8812 3732
rect 8852 3680 8904 3732
rect 10600 3680 10652 3732
rect 6736 3612 6788 3664
rect 9128 3612 9180 3664
rect 10048 3612 10100 3664
rect 7472 3544 7524 3596
rect 7748 3544 7800 3596
rect 8852 3544 8904 3596
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 10968 3544 11020 3596
rect 11152 3612 11204 3664
rect 12992 3612 13044 3664
rect 13176 3680 13228 3732
rect 14096 3680 14148 3732
rect 14280 3680 14332 3732
rect 14464 3612 14516 3664
rect 12532 3544 12584 3596
rect 14556 3587 14608 3596
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15292 3544 15344 3596
rect 17868 3612 17920 3664
rect 18236 3612 18288 3664
rect 19064 3612 19116 3664
rect 16488 3544 16540 3596
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 17592 3544 17644 3596
rect 17776 3544 17828 3596
rect 15108 3476 15160 3528
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 17316 3476 17368 3528
rect 13820 3408 13872 3460
rect 14372 3408 14424 3460
rect 17132 3408 17184 3460
rect 2320 3340 2372 3392
rect 9496 3340 9548 3392
rect 9772 3340 9824 3392
rect 10876 3340 10928 3392
rect 11704 3340 11756 3392
rect 12808 3340 12860 3392
rect 13360 3340 13412 3392
rect 16028 3340 16080 3392
rect 16212 3383 16264 3392
rect 16212 3349 16221 3383
rect 16221 3349 16255 3383
rect 16255 3349 16264 3383
rect 16212 3340 16264 3349
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 19892 3680 19944 3732
rect 19984 3612 20036 3664
rect 18328 3476 18380 3528
rect 19892 3544 19944 3596
rect 20168 3587 20220 3596
rect 20168 3553 20177 3587
rect 20177 3553 20211 3587
rect 20211 3553 20220 3587
rect 20168 3544 20220 3553
rect 21364 3544 21416 3596
rect 21180 3408 21232 3460
rect 17316 3340 17368 3349
rect 18880 3340 18932 3392
rect 20444 3340 20496 3392
rect 20904 3340 20956 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 9036 3136 9088 3188
rect 8760 3068 8812 3120
rect 9680 3068 9732 3120
rect 10968 3136 11020 3188
rect 12900 3136 12952 3188
rect 14464 3136 14516 3188
rect 15108 3179 15160 3188
rect 13636 3068 13688 3120
rect 15108 3145 15117 3179
rect 15117 3145 15151 3179
rect 15151 3145 15160 3179
rect 15108 3136 15160 3145
rect 18696 3136 18748 3188
rect 16580 3068 16632 3120
rect 17960 3068 18012 3120
rect 19156 3136 19208 3188
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 19616 3136 19668 3188
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 8576 3000 8628 3052
rect 9496 3000 9548 3052
rect 9680 2932 9732 2984
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 11520 2932 11572 2984
rect 12624 3000 12676 3052
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 18696 3000 18748 3052
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 19800 3068 19852 3120
rect 19524 3000 19576 3052
rect 11980 2932 12032 2984
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 14372 2932 14424 2984
rect 7840 2864 7892 2916
rect 9956 2864 10008 2916
rect 13084 2864 13136 2916
rect 14648 2864 14700 2916
rect 16856 2932 16908 2984
rect 17684 2932 17736 2984
rect 18052 2932 18104 2984
rect 18972 2932 19024 2984
rect 5632 2796 5684 2848
rect 11612 2796 11664 2848
rect 11704 2796 11756 2848
rect 20536 2864 20588 2916
rect 21824 2864 21876 2916
rect 20904 2796 20956 2848
rect 21732 2796 21784 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 8668 2592 8720 2644
rect 9956 2592 10008 2644
rect 10692 2592 10744 2644
rect 11244 2592 11296 2644
rect 12716 2592 12768 2644
rect 13084 2592 13136 2644
rect 14556 2592 14608 2644
rect 14740 2635 14792 2644
rect 14740 2601 14749 2635
rect 14749 2601 14783 2635
rect 14783 2601 14792 2635
rect 14740 2592 14792 2601
rect 15292 2592 15344 2644
rect 16212 2592 16264 2644
rect 10968 2524 11020 2576
rect 13176 2524 13228 2576
rect 13636 2524 13688 2576
rect 17040 2592 17092 2644
rect 18052 2592 18104 2644
rect 7288 2252 7340 2304
rect 8484 2456 8536 2508
rect 8852 2388 8904 2440
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 12072 2456 12124 2508
rect 12440 2456 12492 2508
rect 13728 2456 13780 2508
rect 17960 2524 18012 2576
rect 11796 2320 11848 2372
rect 19248 2592 19300 2644
rect 19616 2635 19668 2644
rect 19616 2601 19625 2635
rect 19625 2601 19659 2635
rect 19659 2601 19668 2635
rect 19616 2592 19668 2601
rect 18604 2524 18656 2576
rect 20076 2524 20128 2576
rect 21824 2592 21876 2644
rect 20904 2456 20956 2508
rect 14648 2388 14700 2440
rect 16856 2320 16908 2372
rect 17224 2388 17276 2440
rect 16028 2252 16080 2304
rect 17684 2252 17736 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 11152 2048 11204 2100
rect 16396 2048 16448 2100
rect 1768 1368 1820 1420
rect 8760 1368 8812 1420
rect 15476 1368 15528 1420
rect 17224 1368 17276 1420
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 18694 22672 18750 22681
rect 18694 22607 18750 22616
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 5736 19310 5764 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 17236 19394 17264 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 16592 19366 17264 19394
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4066 11520 4122 11529
rect 4066 11455 4122 11464
rect 4080 11354 4108 11455
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 664 9920 716 9926
rect 664 9862 716 9868
rect 202 3496 258 3505
rect 202 3431 258 3440
rect 216 800 244 3431
rect 676 800 704 9862
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 5368 4078 5396 4694
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 1214 3632 1270 3641
rect 1214 3567 1270 3576
rect 1228 800 1256 3567
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 1768 1420 1820 1426
rect 1768 1362 1820 1368
rect 1780 800 1808 1362
rect 2332 800 2360 3334
rect 2884 800 2912 3946
rect 3436 800 3464 4014
rect 5460 4010 5488 4422
rect 7024 4185 7052 19110
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 4826 7236 5646
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7576 4282 7604 5714
rect 8220 5166 8248 6190
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5710 8340 6122
rect 8404 5914 8432 17682
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8312 5370 8340 5646
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4622 7788 5034
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7010 4176 7066 4185
rect 8220 4162 8248 5102
rect 8588 4826 8616 14418
rect 8864 7546 8892 18158
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9600 9926 9628 10134
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9692 9178 9720 14418
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10980 11762 11008 13806
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11072 9568 11100 14894
rect 11256 12594 11284 17070
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11256 12566 11376 12594
rect 11348 12356 11376 12566
rect 11164 12328 11376 12356
rect 11164 9636 11192 12328
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11164 9608 11284 9636
rect 10980 9540 11100 9568
rect 10598 9480 10654 9489
rect 10508 9444 10560 9450
rect 10598 9415 10654 9424
rect 10508 9386 10560 9392
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8772 6458 8800 6802
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 7010 4111 7066 4120
rect 7944 4134 8248 4162
rect 7944 4078 7972 4134
rect 6184 4072 6236 4078
rect 7932 4072 7984 4078
rect 6184 4014 6236 4020
rect 7760 4020 7932 4026
rect 7760 4014 7984 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3988 800 4016 3674
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4802 2952 4858 2961
rect 4802 2887 4858 2896
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1442 4844 2887
rect 4540 1414 4844 1442
rect 4540 800 4568 1414
rect 5092 800 5120 3878
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 800 5672 2790
rect 6196 800 6224 4014
rect 7760 3998 7972 4014
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6748 800 6776 3606
rect 7760 3602 7788 3998
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7484 3058 7512 3538
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7760 2922 7880 2938
rect 7760 2916 7892 2922
rect 7760 2910 7840 2916
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7300 800 7328 2246
rect 7760 1442 7788 2910
rect 7840 2858 7892 2864
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 7760 1414 7880 1442
rect 7852 800 7880 1414
rect 8404 800 8432 4014
rect 8496 2514 8524 4422
rect 8588 3058 8616 4626
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8680 2650 8708 4558
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8772 3738 8800 4490
rect 8864 4010 8892 4558
rect 8956 4282 8984 7686
rect 9048 5370 9076 8910
rect 9508 8634 9536 8910
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9140 5030 9168 5510
rect 9232 5234 9260 8298
rect 10060 8294 10088 8978
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 8090 10088 8230
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 6458 9352 7142
rect 9416 7002 9444 7346
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9508 5574 9536 6122
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8864 3738 8892 3946
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9140 3670 9168 4966
rect 9232 4282 9260 5170
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8864 3194 8892 3538
rect 9508 3398 9536 5510
rect 9600 5030 9628 6054
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4758 9628 4966
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8772 1426 8800 3062
rect 8864 2446 8892 3130
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8760 1420 8812 1426
rect 8760 1362 8812 1368
rect 9048 898 9076 3130
rect 9692 3126 9720 6054
rect 9956 5840 10008 5846
rect 9954 5808 9956 5817
rect 10008 5808 10010 5817
rect 9954 5743 10010 5752
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10060 5234 10088 5714
rect 10048 5228 10100 5234
rect 9968 5188 10048 5216
rect 9968 3602 9996 5188
rect 10048 5170 10100 5176
rect 10428 4282 10456 8774
rect 10520 8090 10548 9386
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10612 6458 10640 9415
rect 10980 9382 11008 9540
rect 11256 9489 11284 9608
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11242 9480 11298 9489
rect 11242 9415 11298 9424
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 8634 11008 8978
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10980 8022 11008 8570
rect 11256 8498 11284 9318
rect 11624 9178 11652 9522
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11716 8090 11744 18770
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11808 8838 11836 11698
rect 12162 11248 12218 11257
rect 12162 11183 12164 11192
rect 12216 11183 12218 11192
rect 12164 11154 12216 11160
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 4826 10732 6122
rect 10888 6118 10916 7142
rect 11164 7002 11192 7346
rect 11256 7342 11284 7754
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11716 7410 11744 7890
rect 11808 7818 11836 8570
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11992 7546 12020 7822
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11348 6798 11376 7278
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 11164 5778 11192 6258
rect 12084 6118 12112 7686
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11796 6112 11848 6118
rect 12072 6112 12124 6118
rect 11796 6054 11848 6060
rect 11992 6072 12072 6100
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5166 11100 5510
rect 11164 5370 11192 5714
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11256 5234 11284 6054
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11256 4622 11284 4966
rect 11716 4758 11744 6054
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 11072 4214 11100 4558
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 4282 11284 4422
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11060 4208 11112 4214
rect 10506 4176 10562 4185
rect 10506 4111 10562 4120
rect 10690 4176 10746 4185
rect 11060 4150 11112 4156
rect 10690 4111 10746 4120
rect 10968 4140 11020 4146
rect 10520 3777 10548 4111
rect 10704 4078 10732 4111
rect 10968 4082 11020 4088
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 3890 10916 4014
rect 10704 3862 10916 3890
rect 10506 3768 10562 3777
rect 10506 3703 10562 3712
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9956 3596 10008 3602
rect 9876 3556 9956 3584
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 8956 870 9076 898
rect 8956 800 8984 870
rect 9508 800 9536 2994
rect 9680 2984 9732 2990
rect 9784 2972 9812 3334
rect 9876 2990 9904 3556
rect 9956 3538 10008 3544
rect 9732 2944 9812 2972
rect 9864 2984 9916 2990
rect 9680 2926 9732 2932
rect 9864 2926 9916 2932
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9968 2650 9996 2858
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10060 800 10088 3606
rect 10612 800 10640 3674
rect 10704 2650 10732 3862
rect 10980 3720 11008 4082
rect 10888 3692 11008 3720
rect 10888 3398 10916 3692
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10980 3194 11008 3538
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10980 2582 11008 3130
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10968 2440 11020 2446
rect 11072 2428 11100 4150
rect 11164 3670 11192 4218
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11256 2650 11284 4014
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11518 3088 11574 3097
rect 11518 3023 11574 3032
rect 11532 2990 11560 3023
rect 11520 2984 11572 2990
rect 11716 2938 11744 3334
rect 11520 2926 11572 2932
rect 11624 2910 11744 2938
rect 11624 2854 11652 2910
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11020 2400 11100 2428
rect 10968 2382 11020 2388
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11164 800 11192 2042
rect 11716 800 11744 2790
rect 11808 2378 11836 6054
rect 11992 4690 12020 6072
rect 12072 6054 12124 6060
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 12084 4146 12112 5510
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12176 4026 12204 9998
rect 12084 3998 12204 4026
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 2990 12020 3470
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 12084 2514 12112 3998
rect 12268 3924 12296 11834
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 9042 12480 10542
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 3942 12388 7686
rect 12452 7410 12480 8978
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 6866 12480 7346
rect 12544 7342 12572 7822
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12544 7002 12572 7278
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12452 5166 12480 5714
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12452 4554 12480 5102
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12176 3896 12296 3924
rect 12348 3936 12400 3942
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 12176 800 12204 3896
rect 12348 3878 12400 3884
rect 12452 3534 12480 4490
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12452 2514 12480 3470
rect 12544 3369 12572 3538
rect 12530 3360 12586 3369
rect 12530 3295 12586 3304
rect 12636 3058 12664 11086
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 7954 12848 8230
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 4826 12756 6054
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12728 4214 12756 4490
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12820 3398 12848 7890
rect 13004 4078 13032 13330
rect 13096 6458 13124 17002
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13188 11354 13216 12310
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11354 13400 12038
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13266 9616 13322 9625
rect 13266 9551 13268 9560
rect 13320 9551 13322 9560
rect 13268 9522 13320 9528
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 7886 13308 9318
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13280 6662 13308 7822
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13372 6338 13400 9930
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13556 7886 13584 9046
rect 13648 9042 13676 9454
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13280 6310 13400 6338
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12912 3194 12940 3878
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13004 3058 13032 3606
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13096 2922 13124 4082
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13188 3058 13216 3674
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 13096 2650 13124 2858
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12728 800 12756 2586
rect 13188 2582 13216 2994
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13280 800 13308 6310
rect 13648 6254 13676 8502
rect 13832 7546 13860 11086
rect 13924 10810 13952 11086
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13924 7410 13952 10474
rect 14016 8090 14044 15506
rect 15212 15026 15240 15506
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10606 14228 10950
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 9994 14228 10542
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13924 7206 13952 7346
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13372 4622 13400 5782
rect 13740 5574 13768 6258
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 5166 13768 5510
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13358 4176 13414 4185
rect 13358 4111 13414 4120
rect 13372 4010 13400 4111
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13360 3392 13412 3398
rect 13358 3360 13360 3369
rect 13412 3360 13414 3369
rect 13358 3295 13414 3304
rect 13648 3126 13676 4422
rect 13924 3641 13952 6122
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5914 14044 6054
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14108 5778 14136 9862
rect 14200 9722 14228 9930
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8362 14228 8774
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4826 14228 4966
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 3738 14136 4082
rect 14292 3738 14320 12786
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15856 12442 15884 18770
rect 16592 13462 16620 19366
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18524 18902 18552 19246
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15028 11762 15056 12242
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15304 11150 15332 11630
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15580 10810 15608 11154
rect 15764 10810 15792 12174
rect 15948 11626 15976 12174
rect 15936 11620 15988 11626
rect 15936 11562 15988 11568
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15764 9926 15792 10474
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 10198 16252 10406
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 14462 9616 14518 9625
rect 14462 9551 14518 9560
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 8090 14412 8366
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14476 7392 14504 9551
rect 15764 9518 15792 9862
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14752 9178 14780 9386
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14752 7886 14780 9114
rect 15396 9042 15424 9318
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15764 7954 15792 9454
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16132 9178 16160 9318
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14384 7364 14504 7392
rect 14384 5914 14412 7364
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14476 6186 14504 7210
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6662 14596 7142
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14384 5817 14412 5850
rect 14370 5808 14426 5817
rect 14370 5743 14426 5752
rect 14384 5166 14412 5743
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14384 4214 14412 5102
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4486 14504 4966
rect 14568 4622 14596 6598
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 13910 3632 13966 3641
rect 13910 3567 13966 3576
rect 14384 3466 14412 4014
rect 14476 3670 14504 4422
rect 14660 4078 14688 7210
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 5710 14780 6598
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 15764 5846 15792 7890
rect 15856 7886 15884 8978
rect 16132 8634 16160 8978
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 16040 7886 16068 8298
rect 16224 8090 16252 9318
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16040 6458 16068 6802
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16040 6322 16068 6394
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15488 5030 15516 5578
rect 15672 5234 15700 5714
rect 16040 5710 16068 6258
rect 16224 5914 16252 7142
rect 16316 6458 16344 7142
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15764 5370 15792 5646
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 13648 2582 13676 3062
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13740 2514 13768 2926
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13832 800 13860 3402
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14384 800 14412 2926
rect 14476 1442 14504 3130
rect 14568 2650 14596 3538
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14660 2446 14688 2858
rect 14752 2650 14780 4014
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15120 3194 15148 3470
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15304 2650 15332 3538
rect 15396 3058 15424 4014
rect 15488 3942 15516 4966
rect 16040 4554 16068 5034
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 16040 3398 16068 4490
rect 16224 4282 16252 4626
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 16224 2650 16252 3334
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 14476 1414 14964 1442
rect 14936 800 14964 1414
rect 15476 1420 15528 1426
rect 15476 1362 15528 1368
rect 15488 800 15516 1362
rect 16040 800 16068 2246
rect 16408 2106 16436 9318
rect 16500 6254 16528 13126
rect 16868 12442 16896 18770
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17972 16726 18000 17070
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18064 15638 18092 16662
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18708 15042 18736 22607
rect 20626 22264 20682 22273
rect 20626 22199 20682 22208
rect 19246 21720 19302 21729
rect 19246 21655 19302 21664
rect 19260 19174 19288 21655
rect 20442 21312 20498 21321
rect 20442 21247 20498 21256
rect 20456 20058 20484 21247
rect 20534 20904 20590 20913
rect 20534 20839 20590 20848
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 20180 18902 20208 19246
rect 20272 18970 20300 19858
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 18786 18048 18842 18057
rect 18786 17983 18842 17992
rect 18800 17338 18828 17983
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18616 15014 18736 15042
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17880 12238 17908 13466
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 12442 18092 12582
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16684 11354 16712 11562
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 8634 16620 10066
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16684 8838 16712 9522
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8430 16712 8774
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16592 6866 16620 7822
rect 16776 7546 16804 11630
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11286 16896 11494
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16868 10674 16896 11222
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16960 10606 16988 11086
rect 17328 10810 17356 12174
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17420 11286 17448 11834
rect 17880 11694 17908 12174
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17880 10606 17908 11630
rect 18156 11354 18184 12242
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 16960 10130 16988 10542
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 17236 9382 17264 10406
rect 17880 9654 17908 10542
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10130 18092 10406
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 18064 9466 18092 10066
rect 18156 9586 18184 10066
rect 18340 10062 18368 10474
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18616 9625 18644 15014
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18708 13870 18736 14894
rect 18800 14634 18828 16594
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 18800 14606 18920 14634
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18800 13394 18828 14418
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18800 11257 18828 11290
rect 18786 11248 18842 11257
rect 18786 11183 18842 11192
rect 18602 9616 18658 9625
rect 18144 9580 18196 9586
rect 18602 9551 18658 9560
rect 18144 9522 18196 9528
rect 18420 9512 18472 9518
rect 18064 9438 18184 9466
rect 18472 9472 18644 9500
rect 18420 9454 18472 9460
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8838 16896 8978
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16684 7002 16712 7346
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16500 5642 16528 6190
rect 16684 5914 16712 6190
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16500 5234 16528 5578
rect 16776 5370 16804 6054
rect 16868 5710 16896 8774
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17236 7954 17264 8230
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17236 7410 17264 7890
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16960 6118 16988 6734
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16868 5370 16896 5646
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16500 4690 16528 4966
rect 16868 4826 16896 5306
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 16856 4820 16908 4826
rect 16592 4758 16620 4789
rect 16856 4762 16908 4768
rect 16580 4752 16632 4758
rect 16578 4720 16580 4729
rect 16632 4720 16634 4729
rect 16488 4684 16540 4690
rect 16578 4655 16634 4664
rect 16488 4626 16540 4632
rect 16592 4570 16620 4655
rect 16500 4542 16620 4570
rect 17040 4616 17092 4622
rect 17144 4593 17172 5102
rect 17040 4558 17092 4564
rect 17130 4584 17186 4593
rect 16500 3602 16528 4542
rect 17052 4486 17080 4558
rect 17130 4519 17186 4528
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16684 3602 16712 4422
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16396 2100 16448 2106
rect 16396 2042 16448 2048
rect 16592 800 16620 3062
rect 16868 2990 16896 3470
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16868 2378 16896 2926
rect 17052 2650 17080 4422
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17144 3942 17172 4082
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 17144 800 17172 3402
rect 17236 2961 17264 7142
rect 17512 6254 17540 8570
rect 17682 7984 17738 7993
rect 17682 7919 17738 7928
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17604 6118 17632 6802
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17604 4622 17632 6054
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17604 4078 17632 4558
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17328 3534 17356 3878
rect 17604 3602 17632 3878
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 3097 17356 3334
rect 17314 3088 17370 3097
rect 17314 3023 17370 3032
rect 17222 2952 17278 2961
rect 17222 2887 17278 2896
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17236 1426 17264 2382
rect 17224 1420 17276 1426
rect 17224 1362 17276 1368
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12714 0 12770 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17604 241 17632 3538
rect 17696 2990 17724 7919
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17880 6662 17908 7686
rect 17972 7342 18000 8774
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17788 3942 17816 5782
rect 17880 5148 17908 5850
rect 17960 5296 18012 5302
rect 17958 5264 17960 5273
rect 18012 5264 18014 5273
rect 17958 5199 18014 5208
rect 17880 5120 18000 5148
rect 17972 4214 18000 5120
rect 17960 4208 18012 4214
rect 17866 4176 17922 4185
rect 17960 4150 18012 4156
rect 17866 4111 17922 4120
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17880 3670 17908 4111
rect 18064 4026 18092 7375
rect 18156 7206 18184 9438
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18616 8566 18644 9472
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 8090 18552 8298
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6254 18184 6598
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18616 5250 18644 8230
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18708 7546 18736 7822
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18524 5222 18644 5250
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 17972 3998 18092 4026
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17788 3482 17816 3538
rect 17972 3482 18000 3998
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17788 3454 18000 3482
rect 17972 3126 18000 3454
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18064 2990 18092 3878
rect 17684 2984 17736 2990
rect 18052 2984 18104 2990
rect 17684 2926 17736 2932
rect 17958 2952 18014 2961
rect 18052 2926 18104 2932
rect 17958 2887 18014 2896
rect 17972 2582 18000 2887
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 800 17724 2246
rect 18064 2009 18092 2586
rect 18050 2000 18106 2009
rect 18050 1935 18106 1944
rect 18156 1442 18184 4966
rect 18524 4729 18552 5222
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18510 4720 18566 4729
rect 18510 4655 18566 4664
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18328 4208 18380 4214
rect 18328 4150 18380 4156
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18248 3670 18276 4082
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18340 3534 18368 4150
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 2582 18644 5102
rect 18708 3913 18736 5714
rect 18800 4486 18828 8910
rect 18892 7818 18920 14606
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19168 11354 19196 12174
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11626 19288 12038
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19352 11218 19380 11494
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19444 11150 19472 11494
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10674 19472 11086
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19444 9518 19472 10406
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19444 9110 19472 9454
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18984 8498 19012 8978
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 19536 7698 19564 12718
rect 19614 9752 19670 9761
rect 19614 9687 19670 9696
rect 19444 7670 19564 7698
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 18892 5030 18920 7142
rect 19168 6934 19196 7142
rect 19246 7032 19302 7041
rect 19246 6967 19302 6976
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 19076 6458 19104 6802
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19076 5710 19104 6394
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 18984 5166 19012 5646
rect 19076 5234 19104 5646
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18878 4720 18934 4729
rect 18878 4655 18934 4664
rect 19064 4684 19116 4690
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18892 4282 18920 4655
rect 19064 4626 19116 4632
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18694 3904 18750 3913
rect 18892 3890 18920 3946
rect 18984 3942 19012 4422
rect 19076 3942 19104 4626
rect 18694 3839 18750 3848
rect 18800 3862 18920 3890
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18694 3224 18750 3233
rect 18694 3159 18696 3168
rect 18748 3159 18750 3168
rect 18696 3130 18748 3136
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18708 2689 18736 2994
rect 18694 2680 18750 2689
rect 18694 2615 18750 2624
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1414 18276 1442
rect 18248 800 18276 1414
rect 18800 800 18828 3862
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3058 18920 3334
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18984 2990 19012 3878
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19076 3369 19104 3606
rect 19062 3360 19118 3369
rect 19062 3295 19118 3304
rect 19168 3194 19196 5306
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 19260 2650 19288 6967
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19352 800 19380 4490
rect 19444 3194 19472 7670
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 19536 5642 19564 7210
rect 19524 5636 19576 5642
rect 19524 5578 19576 5584
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19536 3058 19564 4422
rect 19628 3194 19656 9687
rect 19812 9450 19840 15982
rect 19904 12170 19932 18770
rect 20364 18358 20392 19246
rect 20548 19174 20576 20839
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 20180 17202 20208 17682
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20272 16114 20300 17070
rect 20442 16688 20498 16697
rect 20442 16623 20498 16632
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20456 15706 20484 16623
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20640 14618 20668 22199
rect 21086 20360 21142 20369
rect 21086 20295 21142 20304
rect 21100 20058 21128 20295
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20994 19952 21050 19961
rect 20812 19916 20864 19922
rect 20994 19887 21050 19896
rect 20812 19858 20864 19864
rect 20824 18902 20852 19858
rect 21008 19514 21036 19887
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21086 19408 21142 19417
rect 21086 19343 21142 19352
rect 20994 19000 21050 19009
rect 21100 18970 21128 19343
rect 20994 18935 21050 18944
rect 21088 18964 21140 18970
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20732 17678 20760 18770
rect 21008 18426 21036 18935
rect 21088 18906 21140 18912
rect 21086 18592 21142 18601
rect 21086 18527 21142 18536
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20824 17082 20852 18158
rect 21100 17882 21128 18527
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 20994 17640 21050 17649
rect 20994 17575 21050 17584
rect 21008 17338 21036 17575
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21086 17232 21142 17241
rect 21086 17167 21142 17176
rect 20732 17066 20852 17082
rect 20720 17060 20852 17066
rect 20772 17054 20852 17060
rect 20720 17002 20772 17008
rect 21100 16794 21128 17167
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 20994 16280 21050 16289
rect 20994 16215 20996 16224
rect 21048 16215 21050 16224
rect 20996 16186 21048 16192
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20442 14376 20498 14385
rect 20442 14311 20498 14320
rect 20456 13530 20484 14311
rect 20640 13870 20668 14554
rect 20732 14414 20760 15506
rect 20824 14550 20852 15982
rect 21086 15736 21142 15745
rect 21086 15671 21088 15680
rect 21140 15671 21142 15680
rect 21088 15642 21140 15648
rect 20994 15328 21050 15337
rect 20994 15263 21050 15272
rect 21008 15162 21036 15263
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21086 14920 21142 14929
rect 21086 14855 21142 14864
rect 21100 14618 21128 14855
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 21086 13968 21142 13977
rect 20720 13932 20772 13938
rect 21086 13903 21142 13912
rect 20720 13874 20772 13880
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19996 12782 20024 13262
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19904 10130 19932 11154
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 8974 19748 9318
rect 19904 9042 19932 10066
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19720 8430 19748 8910
rect 19904 8838 19932 8978
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19904 7954 19932 8774
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7342 19748 7822
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7410 19840 7686
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19904 7154 19932 7890
rect 19996 7410 20024 9318
rect 20088 7546 20116 12242
rect 20180 9382 20208 12310
rect 20272 12073 20300 13126
rect 20548 12850 20576 13330
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12374 20484 12718
rect 20640 12646 20668 12677
rect 20628 12640 20680 12646
rect 20626 12608 20628 12617
rect 20680 12608 20682 12617
rect 20626 12543 20682 12552
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20258 12064 20314 12073
rect 20258 11999 20314 12008
rect 20272 11354 20300 11999
rect 20640 11694 20668 12543
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20258 11248 20314 11257
rect 20258 11183 20314 11192
rect 20272 10266 20300 11183
rect 20364 11150 20392 11562
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20534 10296 20590 10305
rect 20260 10260 20312 10266
rect 20534 10231 20590 10240
rect 20260 10202 20312 10208
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20272 8090 20300 10202
rect 20548 9178 20576 10231
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20640 8634 20668 9386
rect 20732 8906 20760 13874
rect 21100 13530 21128 13903
rect 21270 13560 21326 13569
rect 21088 13524 21140 13530
rect 21270 13495 21326 13504
rect 21088 13466 21140 13472
rect 21086 13016 21142 13025
rect 21284 12986 21312 13495
rect 21086 12951 21142 12960
rect 21272 12980 21324 12986
rect 21100 12442 21128 12951
rect 21272 12922 21324 12928
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20916 11898 20944 12242
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20902 11656 20958 11665
rect 20902 11591 20904 11600
rect 20956 11591 20958 11600
rect 20904 11562 20956 11568
rect 20916 11218 20944 11562
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20902 10704 20958 10713
rect 20902 10639 20958 10648
rect 20916 10130 20944 10639
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21100 10198 21128 10406
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20916 8634 20944 10066
rect 21362 9344 21418 9353
rect 21362 9279 21418 9288
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20534 8392 20590 8401
rect 20534 8327 20590 8336
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20272 7478 20300 7822
rect 20260 7472 20312 7478
rect 20260 7414 20312 7420
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 19720 7126 19932 7154
rect 19720 3505 19748 7126
rect 19996 7002 20024 7346
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19996 5370 20024 5714
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 19812 4282 19840 4694
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19706 3496 19762 3505
rect 19706 3431 19762 3440
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19628 2650 19656 3130
rect 19812 3126 19840 4218
rect 19904 3738 19932 4626
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 4282 20024 4558
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19982 3768 20038 3777
rect 19892 3732 19944 3738
rect 19982 3703 20038 3712
rect 19892 3674 19944 3680
rect 19996 3670 20024 3703
rect 19984 3664 20036 3670
rect 19984 3606 20036 3612
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19904 3505 19932 3538
rect 19890 3496 19946 3505
rect 19890 3431 19946 3440
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 20088 2582 20116 7142
rect 20180 6730 20208 7346
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20180 6186 20208 6666
rect 20272 6633 20300 7414
rect 20258 6624 20314 6633
rect 20258 6559 20314 6568
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20364 5710 20392 6054
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20364 5234 20392 5646
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20180 4010 20208 4422
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20076 2576 20128 2582
rect 20076 2518 20128 2524
rect 20180 2417 20208 3538
rect 20364 2961 20392 4966
rect 20456 4146 20484 6054
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20456 3398 20484 4082
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20350 2952 20406 2961
rect 20548 2922 20576 8327
rect 20640 7886 20668 8570
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20732 6746 20760 7142
rect 20732 6718 20852 6746
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20350 2887 20406 2896
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 20166 2408 20222 2417
rect 20166 2343 20222 2352
rect 20640 921 20668 6598
rect 20824 5302 20852 6718
rect 20994 6080 21050 6089
rect 20994 6015 21050 6024
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20812 5296 20864 5302
rect 20916 5273 20944 5714
rect 20812 5238 20864 5244
rect 20902 5264 20958 5273
rect 20902 5199 20958 5208
rect 21008 5166 21036 6015
rect 21270 5672 21326 5681
rect 21270 5607 21326 5616
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 21008 4826 21036 5102
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20902 4584 20958 4593
rect 20902 4519 20958 4528
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 19890 912 19946 921
rect 19890 847 19946 856
rect 20442 912 20498 921
rect 20442 847 20498 856
rect 20626 912 20682 921
rect 20626 847 20682 856
rect 19904 800 19932 847
rect 20456 800 20484 847
rect 17590 232 17646 241
rect 17590 167 17646 176
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19890 0 19946 800
rect 20442 0 20498 800
rect 20824 649 20852 4014
rect 20916 3942 20944 4519
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20994 3496 21050 3505
rect 20994 3431 21050 3440
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20916 3233 20944 3334
rect 20902 3224 20958 3233
rect 20902 3159 20958 3168
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20916 2514 20944 2790
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 21008 800 21036 3431
rect 21100 1057 21128 5510
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21192 4486 21220 4966
rect 21284 4690 21312 5607
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21180 4480 21232 4486
rect 21180 4422 21232 4428
rect 21284 3777 21312 4626
rect 21376 4146 21404 9279
rect 21730 8936 21786 8945
rect 21730 8871 21786 8880
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21270 3768 21326 3777
rect 21270 3703 21326 3712
rect 21376 3602 21404 4082
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 21192 2689 21220 3402
rect 21178 2680 21234 2689
rect 21178 2615 21234 2624
rect 21192 1601 21220 2615
rect 21468 2009 21496 5034
rect 21454 2000 21510 2009
rect 21454 1935 21510 1944
rect 21178 1592 21234 1601
rect 21178 1527 21234 1536
rect 21086 1048 21142 1057
rect 21086 983 21142 992
rect 21560 800 21588 5578
rect 21652 4214 21680 5646
rect 21640 4208 21692 4214
rect 21640 4150 21692 4156
rect 21652 1057 21680 4150
rect 21744 2854 21772 8871
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22020 4729 22048 5510
rect 22006 4720 22062 4729
rect 22006 4655 22062 4664
rect 21824 2916 21876 2922
rect 21824 2858 21876 2864
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21836 2650 21864 2858
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21638 1048 21694 1057
rect 21638 983 21694 992
rect 22112 800 22140 11494
rect 22650 3632 22706 3641
rect 22650 3567 22706 3576
rect 22664 800 22692 3567
rect 20810 640 20866 649
rect 20810 575 20866 584
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
<< via2 >>
rect 18694 22616 18750 22672
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4066 11464 4122 11520
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 202 3440 258 3496
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 1214 3576 1270 3632
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7010 4120 7066 4176
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10598 9424 10654 9480
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4802 2896 4858 2952
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 9954 5788 9956 5808
rect 9956 5788 10008 5808
rect 10008 5788 10010 5808
rect 9954 5752 10010 5788
rect 11242 9424 11298 9480
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 12162 11212 12218 11248
rect 12162 11192 12164 11212
rect 12164 11192 12216 11212
rect 12216 11192 12218 11212
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 10506 4120 10562 4176
rect 10690 4120 10746 4176
rect 10506 3712 10562 3768
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11518 3032 11574 3088
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12530 3304 12586 3360
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 13266 9580 13322 9616
rect 13266 9560 13268 9580
rect 13268 9560 13320 9580
rect 13320 9560 13322 9580
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 13358 4120 13414 4176
rect 13358 3340 13360 3360
rect 13360 3340 13412 3360
rect 13412 3340 13414 3360
rect 13358 3304 13414 3340
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14462 9560 14518 9616
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14370 5752 14426 5808
rect 13910 3576 13966 3632
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 20626 22208 20682 22264
rect 19246 21664 19302 21720
rect 20442 21256 20498 21312
rect 20534 20848 20590 20904
rect 18786 17992 18842 18048
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18786 11192 18842 11248
rect 18602 9560 18658 9616
rect 16578 4700 16580 4720
rect 16580 4700 16632 4720
rect 16632 4700 16634 4720
rect 16578 4664 16634 4700
rect 17130 4528 17186 4584
rect 17682 7928 17738 7984
rect 17314 3032 17370 3088
rect 17222 2896 17278 2952
rect 18050 7384 18106 7440
rect 17958 5244 17960 5264
rect 17960 5244 18012 5264
rect 18012 5244 18014 5264
rect 17958 5208 18014 5244
rect 17866 4120 17922 4176
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 17958 2896 18014 2952
rect 18050 1944 18106 2000
rect 18510 4664 18566 4720
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 19614 9696 19670 9752
rect 19246 6976 19302 7032
rect 18878 4664 18934 4720
rect 18694 3848 18750 3904
rect 18694 3188 18750 3224
rect 18694 3168 18696 3188
rect 18696 3168 18748 3188
rect 18748 3168 18750 3188
rect 18694 2624 18750 2680
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19062 3304 19118 3360
rect 20442 16632 20498 16688
rect 21086 20304 21142 20360
rect 20994 19896 21050 19952
rect 21086 19352 21142 19408
rect 20994 18944 21050 19000
rect 21086 18536 21142 18592
rect 20994 17584 21050 17640
rect 21086 17176 21142 17232
rect 20994 16244 21050 16280
rect 20994 16224 20996 16244
rect 20996 16224 21048 16244
rect 21048 16224 21050 16244
rect 20442 14320 20498 14376
rect 21086 15700 21142 15736
rect 21086 15680 21088 15700
rect 21088 15680 21140 15700
rect 21140 15680 21142 15700
rect 20994 15272 21050 15328
rect 21086 14864 21142 14920
rect 21086 13912 21142 13968
rect 20626 12588 20628 12608
rect 20628 12588 20680 12608
rect 20680 12588 20682 12608
rect 20626 12552 20682 12588
rect 20258 12008 20314 12064
rect 20258 11192 20314 11248
rect 20534 10240 20590 10296
rect 21270 13504 21326 13560
rect 21086 12960 21142 13016
rect 20902 11620 20958 11656
rect 20902 11600 20904 11620
rect 20904 11600 20956 11620
rect 20956 11600 20958 11620
rect 20902 10648 20958 10704
rect 21362 9288 21418 9344
rect 20534 8336 20590 8392
rect 19706 3440 19762 3496
rect 19982 3712 20038 3768
rect 19890 3440 19946 3496
rect 20258 6568 20314 6624
rect 20350 2896 20406 2952
rect 20166 2352 20222 2408
rect 20994 6024 21050 6080
rect 20902 5208 20958 5264
rect 21270 5616 21326 5672
rect 20902 4528 20958 4584
rect 19890 856 19946 912
rect 20442 856 20498 912
rect 20626 856 20682 912
rect 17590 176 17646 232
rect 20994 3440 21050 3496
rect 20902 3168 20958 3224
rect 21730 8880 21786 8936
rect 21270 3712 21326 3768
rect 21178 2624 21234 2680
rect 21454 1944 21510 2000
rect 21178 1536 21234 1592
rect 21086 992 21142 1048
rect 22006 4664 22062 4720
rect 21638 992 21694 1048
rect 22650 3576 22706 3632
rect 20810 584 20866 640
<< metal3 >>
rect 18689 22674 18755 22677
rect 22200 22674 23000 22704
rect 18689 22672 23000 22674
rect 18689 22616 18694 22672
rect 18750 22616 23000 22672
rect 18689 22614 23000 22616
rect 18689 22611 18755 22614
rect 22200 22584 23000 22614
rect 20621 22266 20687 22269
rect 22200 22266 23000 22296
rect 20621 22264 23000 22266
rect 20621 22208 20626 22264
rect 20682 22208 23000 22264
rect 20621 22206 23000 22208
rect 20621 22203 20687 22206
rect 22200 22176 23000 22206
rect 19241 21722 19307 21725
rect 22200 21722 23000 21752
rect 19241 21720 23000 21722
rect 19241 21664 19246 21720
rect 19302 21664 23000 21720
rect 19241 21662 23000 21664
rect 19241 21659 19307 21662
rect 22200 21632 23000 21662
rect 20437 21314 20503 21317
rect 22200 21314 23000 21344
rect 20437 21312 23000 21314
rect 20437 21256 20442 21312
rect 20498 21256 23000 21312
rect 20437 21254 23000 21256
rect 20437 21251 20503 21254
rect 22200 21224 23000 21254
rect 20529 20906 20595 20909
rect 22200 20906 23000 20936
rect 20529 20904 23000 20906
rect 20529 20848 20534 20904
rect 20590 20848 23000 20904
rect 20529 20846 23000 20848
rect 20529 20843 20595 20846
rect 22200 20816 23000 20846
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 21081 20362 21147 20365
rect 22200 20362 23000 20392
rect 21081 20360 23000 20362
rect 21081 20304 21086 20360
rect 21142 20304 23000 20360
rect 21081 20302 23000 20304
rect 21081 20299 21147 20302
rect 22200 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 20989 19954 21055 19957
rect 22200 19954 23000 19984
rect 20989 19952 23000 19954
rect 20989 19896 20994 19952
rect 21050 19896 23000 19952
rect 20989 19894 23000 19896
rect 20989 19891 21055 19894
rect 22200 19864 23000 19894
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 21081 19410 21147 19413
rect 22200 19410 23000 19440
rect 21081 19408 23000 19410
rect 21081 19352 21086 19408
rect 21142 19352 23000 19408
rect 21081 19350 23000 19352
rect 21081 19347 21147 19350
rect 22200 19320 23000 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 20989 19002 21055 19005
rect 22200 19002 23000 19032
rect 20989 19000 23000 19002
rect 20989 18944 20994 19000
rect 21050 18944 23000 19000
rect 20989 18942 23000 18944
rect 20989 18939 21055 18942
rect 22200 18912 23000 18942
rect 21081 18594 21147 18597
rect 22200 18594 23000 18624
rect 21081 18592 23000 18594
rect 21081 18536 21086 18592
rect 21142 18536 23000 18592
rect 21081 18534 23000 18536
rect 21081 18531 21147 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 22200 18504 23000 18534
rect 18270 18463 18590 18464
rect 18781 18050 18847 18053
rect 22200 18050 23000 18080
rect 18781 18048 23000 18050
rect 18781 17992 18786 18048
rect 18842 17992 23000 18048
rect 18781 17990 23000 17992
rect 18781 17987 18847 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 20989 17642 21055 17645
rect 22200 17642 23000 17672
rect 20989 17640 23000 17642
rect 20989 17584 20994 17640
rect 21050 17584 23000 17640
rect 20989 17582 23000 17584
rect 20989 17579 21055 17582
rect 22200 17552 23000 17582
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 21081 17234 21147 17237
rect 22200 17234 23000 17264
rect 21081 17232 23000 17234
rect 21081 17176 21086 17232
rect 21142 17176 23000 17232
rect 21081 17174 23000 17176
rect 21081 17171 21147 17174
rect 22200 17144 23000 17174
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 20437 16690 20503 16693
rect 22200 16690 23000 16720
rect 20437 16688 23000 16690
rect 20437 16632 20442 16688
rect 20498 16632 23000 16688
rect 20437 16630 23000 16632
rect 20437 16627 20503 16630
rect 22200 16600 23000 16630
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 20989 16282 21055 16285
rect 22200 16282 23000 16312
rect 20989 16280 23000 16282
rect 20989 16224 20994 16280
rect 21050 16224 23000 16280
rect 20989 16222 23000 16224
rect 20989 16219 21055 16222
rect 22200 16192 23000 16222
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 21081 15738 21147 15741
rect 22200 15738 23000 15768
rect 21081 15736 23000 15738
rect 21081 15680 21086 15736
rect 21142 15680 23000 15736
rect 21081 15678 23000 15680
rect 21081 15675 21147 15678
rect 22200 15648 23000 15678
rect 20989 15330 21055 15333
rect 22200 15330 23000 15360
rect 20989 15328 23000 15330
rect 20989 15272 20994 15328
rect 21050 15272 23000 15328
rect 20989 15270 23000 15272
rect 20989 15267 21055 15270
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 22200 15240 23000 15270
rect 18270 15199 18590 15200
rect 21081 14922 21147 14925
rect 22200 14922 23000 14952
rect 21081 14920 23000 14922
rect 21081 14864 21086 14920
rect 21142 14864 23000 14920
rect 21081 14862 23000 14864
rect 21081 14859 21147 14862
rect 22200 14832 23000 14862
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 20437 14378 20503 14381
rect 22200 14378 23000 14408
rect 20437 14376 23000 14378
rect 20437 14320 20442 14376
rect 20498 14320 23000 14376
rect 20437 14318 23000 14320
rect 20437 14315 20503 14318
rect 22200 14288 23000 14318
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 21081 13970 21147 13973
rect 22200 13970 23000 14000
rect 21081 13968 23000 13970
rect 21081 13912 21086 13968
rect 21142 13912 23000 13968
rect 21081 13910 23000 13912
rect 21081 13907 21147 13910
rect 22200 13880 23000 13910
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 21265 13562 21331 13565
rect 22200 13562 23000 13592
rect 21265 13560 23000 13562
rect 21265 13504 21270 13560
rect 21326 13504 23000 13560
rect 21265 13502 23000 13504
rect 21265 13499 21331 13502
rect 22200 13472 23000 13502
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 21081 13018 21147 13021
rect 22200 13018 23000 13048
rect 21081 13016 23000 13018
rect 21081 12960 21086 13016
rect 21142 12960 23000 13016
rect 21081 12958 23000 12960
rect 21081 12955 21147 12958
rect 22200 12928 23000 12958
rect 20621 12610 20687 12613
rect 22200 12610 23000 12640
rect 20621 12608 23000 12610
rect 20621 12552 20626 12608
rect 20682 12552 23000 12608
rect 20621 12550 23000 12552
rect 20621 12547 20687 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 22200 12520 23000 12550
rect 14805 12479 15125 12480
rect 20253 12066 20319 12069
rect 22200 12066 23000 12096
rect 20253 12064 23000 12066
rect 20253 12008 20258 12064
rect 20314 12008 23000 12064
rect 20253 12006 23000 12008
rect 20253 12003 20319 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 22200 11976 23000 12006
rect 18270 11935 18590 11936
rect 20897 11658 20963 11661
rect 22200 11658 23000 11688
rect 20897 11656 23000 11658
rect 20897 11600 20902 11656
rect 20958 11600 23000 11656
rect 20897 11598 23000 11600
rect 20897 11595 20963 11598
rect 22200 11568 23000 11598
rect 0 11522 800 11552
rect 4061 11522 4127 11525
rect 0 11520 4127 11522
rect 0 11464 4066 11520
rect 4122 11464 4127 11520
rect 0 11462 4127 11464
rect 0 11432 800 11462
rect 4061 11459 4127 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 12157 11250 12223 11253
rect 18781 11250 18847 11253
rect 12157 11248 18847 11250
rect 12157 11192 12162 11248
rect 12218 11192 18786 11248
rect 18842 11192 18847 11248
rect 12157 11190 18847 11192
rect 12157 11187 12223 11190
rect 18781 11187 18847 11190
rect 20253 11250 20319 11253
rect 22200 11250 23000 11280
rect 20253 11248 23000 11250
rect 20253 11192 20258 11248
rect 20314 11192 23000 11248
rect 20253 11190 23000 11192
rect 20253 11187 20319 11190
rect 22200 11160 23000 11190
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 20897 10706 20963 10709
rect 22200 10706 23000 10736
rect 20897 10704 23000 10706
rect 20897 10648 20902 10704
rect 20958 10648 23000 10704
rect 20897 10646 23000 10648
rect 20897 10643 20963 10646
rect 22200 10616 23000 10646
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 20529 10298 20595 10301
rect 22200 10298 23000 10328
rect 20529 10296 23000 10298
rect 20529 10240 20534 10296
rect 20590 10240 23000 10296
rect 20529 10238 23000 10240
rect 20529 10235 20595 10238
rect 22200 10208 23000 10238
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 19609 9754 19675 9757
rect 22200 9754 23000 9784
rect 19609 9752 23000 9754
rect 19609 9696 19614 9752
rect 19670 9696 23000 9752
rect 19609 9694 23000 9696
rect 19609 9691 19675 9694
rect 22200 9664 23000 9694
rect 13261 9618 13327 9621
rect 14457 9618 14523 9621
rect 18597 9618 18663 9621
rect 13261 9616 18663 9618
rect 13261 9560 13266 9616
rect 13322 9560 14462 9616
rect 14518 9560 18602 9616
rect 18658 9560 18663 9616
rect 13261 9558 18663 9560
rect 13261 9555 13327 9558
rect 14457 9555 14523 9558
rect 18597 9555 18663 9558
rect 10593 9482 10659 9485
rect 11237 9482 11303 9485
rect 10593 9480 11303 9482
rect 10593 9424 10598 9480
rect 10654 9424 11242 9480
rect 11298 9424 11303 9480
rect 10593 9422 11303 9424
rect 10593 9419 10659 9422
rect 11237 9419 11303 9422
rect 21357 9346 21423 9349
rect 22200 9346 23000 9376
rect 21357 9344 23000 9346
rect 21357 9288 21362 9344
rect 21418 9288 23000 9344
rect 21357 9286 23000 9288
rect 21357 9283 21423 9286
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 22200 9256 23000 9286
rect 14805 9215 15125 9216
rect 21725 8938 21791 8941
rect 22200 8938 23000 8968
rect 21725 8936 23000 8938
rect 21725 8880 21730 8936
rect 21786 8880 23000 8936
rect 21725 8878 23000 8880
rect 21725 8875 21791 8878
rect 22200 8848 23000 8878
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 20529 8394 20595 8397
rect 22200 8394 23000 8424
rect 20529 8392 23000 8394
rect 20529 8336 20534 8392
rect 20590 8336 23000 8392
rect 20529 8334 23000 8336
rect 20529 8331 20595 8334
rect 22200 8304 23000 8334
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 17677 7986 17743 7989
rect 22200 7986 23000 8016
rect 17677 7984 23000 7986
rect 17677 7928 17682 7984
rect 17738 7928 23000 7984
rect 17677 7926 23000 7928
rect 17677 7923 17743 7926
rect 22200 7896 23000 7926
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 22200 7578 23000 7608
rect 18692 7518 23000 7578
rect 18045 7442 18111 7445
rect 18692 7442 18752 7518
rect 22200 7488 23000 7518
rect 18045 7440 18752 7442
rect 18045 7384 18050 7440
rect 18106 7384 18752 7440
rect 18045 7382 18752 7384
rect 18045 7379 18111 7382
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 19241 7034 19307 7037
rect 22200 7034 23000 7064
rect 19241 7032 23000 7034
rect 19241 6976 19246 7032
rect 19302 6976 23000 7032
rect 19241 6974 23000 6976
rect 19241 6971 19307 6974
rect 22200 6944 23000 6974
rect 20253 6626 20319 6629
rect 22200 6626 23000 6656
rect 20253 6624 23000 6626
rect 20253 6568 20258 6624
rect 20314 6568 23000 6624
rect 20253 6566 23000 6568
rect 20253 6563 20319 6566
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 22200 6536 23000 6566
rect 18270 6495 18590 6496
rect 20989 6082 21055 6085
rect 22200 6082 23000 6112
rect 20989 6080 23000 6082
rect 20989 6024 20994 6080
rect 21050 6024 23000 6080
rect 20989 6022 23000 6024
rect 20989 6019 21055 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 22200 5992 23000 6022
rect 14805 5951 15125 5952
rect 9949 5810 10015 5813
rect 14365 5810 14431 5813
rect 9949 5808 14431 5810
rect 9949 5752 9954 5808
rect 10010 5752 14370 5808
rect 14426 5752 14431 5808
rect 9949 5750 14431 5752
rect 9949 5747 10015 5750
rect 14365 5747 14431 5750
rect 21265 5674 21331 5677
rect 22200 5674 23000 5704
rect 21265 5672 23000 5674
rect 21265 5616 21270 5672
rect 21326 5616 23000 5672
rect 21265 5614 23000 5616
rect 21265 5611 21331 5614
rect 22200 5584 23000 5614
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 17953 5266 18019 5269
rect 20897 5266 20963 5269
rect 22200 5266 23000 5296
rect 17953 5264 23000 5266
rect 17953 5208 17958 5264
rect 18014 5208 20902 5264
rect 20958 5208 23000 5264
rect 17953 5206 23000 5208
rect 17953 5203 18019 5206
rect 20897 5203 20963 5206
rect 22200 5176 23000 5206
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 16573 4722 16639 4725
rect 18505 4722 18571 4725
rect 18873 4722 18939 4725
rect 16573 4720 18939 4722
rect 16573 4664 16578 4720
rect 16634 4664 18510 4720
rect 18566 4664 18878 4720
rect 18934 4664 18939 4720
rect 16573 4662 18939 4664
rect 16573 4659 16639 4662
rect 18505 4659 18571 4662
rect 18873 4659 18939 4662
rect 22001 4722 22067 4725
rect 22200 4722 23000 4752
rect 22001 4720 23000 4722
rect 22001 4664 22006 4720
rect 22062 4664 23000 4720
rect 22001 4662 23000 4664
rect 22001 4659 22067 4662
rect 22200 4632 23000 4662
rect 17125 4586 17191 4589
rect 20897 4586 20963 4589
rect 17125 4584 20963 4586
rect 17125 4528 17130 4584
rect 17186 4528 20902 4584
rect 20958 4528 20963 4584
rect 17125 4526 20963 4528
rect 17125 4523 17191 4526
rect 20897 4523 20963 4526
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 22200 4314 23000 4344
rect 18692 4254 23000 4314
rect 7005 4178 7071 4181
rect 10501 4178 10567 4181
rect 7005 4176 10567 4178
rect 7005 4120 7010 4176
rect 7066 4120 10506 4176
rect 10562 4120 10567 4176
rect 7005 4118 10567 4120
rect 7005 4115 7071 4118
rect 10501 4115 10567 4118
rect 10685 4178 10751 4181
rect 13353 4178 13419 4181
rect 10685 4176 13419 4178
rect 10685 4120 10690 4176
rect 10746 4120 13358 4176
rect 13414 4120 13419 4176
rect 10685 4118 13419 4120
rect 10685 4115 10751 4118
rect 13353 4115 13419 4118
rect 17861 4178 17927 4181
rect 18692 4178 18752 4254
rect 22200 4224 23000 4254
rect 17861 4176 18752 4178
rect 17861 4120 17866 4176
rect 17922 4120 18752 4176
rect 17861 4118 18752 4120
rect 17861 4115 17927 4118
rect 18689 3906 18755 3909
rect 22200 3906 23000 3936
rect 18689 3904 23000 3906
rect 18689 3848 18694 3904
rect 18750 3848 23000 3904
rect 18689 3846 23000 3848
rect 18689 3843 18755 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 10501 3770 10567 3773
rect 19977 3770 20043 3773
rect 21265 3770 21331 3773
rect 10501 3768 14106 3770
rect 10501 3712 10506 3768
rect 10562 3712 14106 3768
rect 10501 3710 14106 3712
rect 10501 3707 10567 3710
rect 1209 3634 1275 3637
rect 13905 3634 13971 3637
rect 1209 3632 13971 3634
rect 1209 3576 1214 3632
rect 1270 3576 13910 3632
rect 13966 3576 13971 3632
rect 1209 3574 13971 3576
rect 14046 3634 14106 3710
rect 19977 3768 21331 3770
rect 19977 3712 19982 3768
rect 20038 3712 21270 3768
rect 21326 3712 21331 3768
rect 19977 3710 21331 3712
rect 19977 3707 20043 3710
rect 21265 3707 21331 3710
rect 22645 3634 22711 3637
rect 14046 3632 22711 3634
rect 14046 3576 22650 3632
rect 22706 3576 22711 3632
rect 14046 3574 22711 3576
rect 1209 3571 1275 3574
rect 13905 3571 13971 3574
rect 22645 3571 22711 3574
rect 197 3498 263 3501
rect 19701 3498 19767 3501
rect 197 3496 19767 3498
rect 197 3440 202 3496
rect 258 3440 19706 3496
rect 19762 3440 19767 3496
rect 197 3438 19767 3440
rect 197 3435 263 3438
rect 19701 3435 19767 3438
rect 19885 3498 19951 3501
rect 20989 3498 21055 3501
rect 19885 3496 21055 3498
rect 19885 3440 19890 3496
rect 19946 3440 20994 3496
rect 21050 3440 21055 3496
rect 19885 3438 21055 3440
rect 19885 3435 19951 3438
rect 20989 3435 21055 3438
rect 12525 3362 12591 3365
rect 13353 3362 13419 3365
rect 12525 3360 13419 3362
rect 12525 3304 12530 3360
rect 12586 3304 13358 3360
rect 13414 3304 13419 3360
rect 12525 3302 13419 3304
rect 12525 3299 12591 3302
rect 13353 3299 13419 3302
rect 19057 3362 19123 3365
rect 22200 3362 23000 3392
rect 19057 3360 23000 3362
rect 19057 3304 19062 3360
rect 19118 3304 23000 3360
rect 19057 3302 23000 3304
rect 19057 3299 19123 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 22200 3272 23000 3302
rect 18270 3231 18590 3232
rect 18689 3226 18755 3229
rect 20897 3226 20963 3229
rect 18689 3224 20963 3226
rect 18689 3168 18694 3224
rect 18750 3168 20902 3224
rect 20958 3168 20963 3224
rect 18689 3166 20963 3168
rect 18689 3163 18755 3166
rect 20897 3163 20963 3166
rect 11513 3090 11579 3093
rect 17309 3090 17375 3093
rect 11513 3088 17375 3090
rect 11513 3032 11518 3088
rect 11574 3032 17314 3088
rect 17370 3032 17375 3088
rect 11513 3030 17375 3032
rect 11513 3027 11579 3030
rect 17309 3027 17375 3030
rect 4797 2954 4863 2957
rect 17217 2954 17283 2957
rect 4797 2952 17283 2954
rect 4797 2896 4802 2952
rect 4858 2896 17222 2952
rect 17278 2896 17283 2952
rect 4797 2894 17283 2896
rect 4797 2891 4863 2894
rect 17217 2891 17283 2894
rect 17953 2954 18019 2957
rect 20345 2954 20411 2957
rect 22200 2954 23000 2984
rect 17953 2952 23000 2954
rect 17953 2896 17958 2952
rect 18014 2896 20350 2952
rect 20406 2896 23000 2952
rect 17953 2894 23000 2896
rect 17953 2891 18019 2894
rect 20345 2891 20411 2894
rect 22200 2864 23000 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 18689 2682 18755 2685
rect 21173 2682 21239 2685
rect 18689 2680 21239 2682
rect 18689 2624 18694 2680
rect 18750 2624 21178 2680
rect 21234 2624 21239 2680
rect 18689 2622 21239 2624
rect 18689 2619 18755 2622
rect 21173 2619 21239 2622
rect 20161 2410 20227 2413
rect 22200 2410 23000 2440
rect 20161 2408 23000 2410
rect 20161 2352 20166 2408
rect 20222 2352 23000 2408
rect 20161 2350 23000 2352
rect 20161 2347 20227 2350
rect 22200 2320 23000 2350
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 18045 2002 18111 2005
rect 21449 2002 21515 2005
rect 22200 2002 23000 2032
rect 18045 2000 23000 2002
rect 18045 1944 18050 2000
rect 18106 1944 21454 2000
rect 21510 1944 23000 2000
rect 18045 1942 23000 1944
rect 18045 1939 18111 1942
rect 21449 1939 21515 1942
rect 22200 1912 23000 1942
rect 21173 1594 21239 1597
rect 22200 1594 23000 1624
rect 21173 1592 23000 1594
rect 21173 1536 21178 1592
rect 21234 1536 23000 1592
rect 21173 1534 23000 1536
rect 21173 1531 21239 1534
rect 22200 1504 23000 1534
rect 21081 1050 21147 1053
rect 19934 1048 21147 1050
rect 19934 992 21086 1048
rect 21142 992 21147 1048
rect 19934 990 21147 992
rect 19934 917 19994 990
rect 21081 987 21147 990
rect 21633 1050 21699 1053
rect 22200 1050 23000 1080
rect 21633 1048 23000 1050
rect 21633 992 21638 1048
rect 21694 992 23000 1048
rect 21633 990 23000 992
rect 21633 987 21699 990
rect 22200 960 23000 990
rect 19885 912 19994 917
rect 19885 856 19890 912
rect 19946 856 19994 912
rect 19885 854 19994 856
rect 20437 914 20503 917
rect 20621 914 20687 917
rect 20437 912 20687 914
rect 20437 856 20442 912
rect 20498 856 20626 912
rect 20682 856 20687 912
rect 20437 854 20687 856
rect 19885 851 19951 854
rect 20437 851 20503 854
rect 20621 851 20687 854
rect 20805 642 20871 645
rect 22200 642 23000 672
rect 20805 640 23000 642
rect 20805 584 20810 640
rect 20866 584 23000 640
rect 20805 582 23000 584
rect 20805 579 20871 582
rect 22200 552 23000 582
rect 17585 234 17651 237
rect 22200 234 23000 264
rect 17585 232 23000 234
rect 17585 176 17590 232
rect 17646 176 23000 232
rect 17585 174 23000 176
rect 17585 171 17651 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608910539
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608910539
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608910539
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7360 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_83
timestamp 1608910539
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1608910539
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1608910539
transform 1 0 7452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7452 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1608910539
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1608910539
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608910539
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _42_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9108 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1608910539
transform 1 0 9752 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1608910539
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96
timestamp 1608910539
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9844 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_111
timestamp 1608910539
transform 1 0 11316 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_111
timestamp 1608910539
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1608910539
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_115
timestamp 1608910539
transform 1 0 11684 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1608910539
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1608910539
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1608910539
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12512 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1608910539
transform 1 0 13340 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1608910539
transform 1 0 14076 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14352 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13708 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_153
timestamp 1608910539
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1608910539
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608910539
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15364 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1608910539
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1608910539
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1608910539
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1608910539
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16468 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_186
timestamp 1608910539
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1608910539
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608910539
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608910539
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608910539
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1608910539
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_189
timestamp 1608910539
transform 1 0 18492 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18400 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 18768 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1608910539
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_198
timestamp 1608910539
transform 1 0 19320 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1608910539
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 19412 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608910539
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1608910539
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_212
timestamp 1608910539
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1608910539
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1608910539
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608910539
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_218
timestamp 1608910539
transform 1 0 21160 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1608910539
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608910539
transform 1 0 20792 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1608910539
transform 1 0 21528 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_220
timestamp 1608910539
transform 1 0 21344 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608910539
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608910539
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608910539
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp 1608910539
transform 1 0 7360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7636 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1608910539
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1608910539
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9936 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1608910539
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1608910539
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1608910539
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1608910539
transform 1 0 11960 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_139
timestamp 1608910539
transform 1 0 13892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp 1608910539
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_156
timestamp 1608910539
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608910539
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16192 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1608910539
transform 1 0 15640 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1608910539
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_178
timestamp 1608910539
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_173
timestamp 1608910539
transform 1 0 17020 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608910539
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1608910539
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1608910539
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1608910539
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 18400 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 19780 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1608910539
transform 1 0 21252 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1608910539
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608910539
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608910539
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1608910539
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_67
timestamp 1608910539
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1608910539
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1608910539
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1608910539
transform 1 0 9292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10396 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608910539
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_114
timestamp 1608910539
transform 1 0 11592 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1608910539
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1608910539
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1608910539
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1608910539
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1608910539
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1608910539
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15916 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608910539
transform 1 0 14536 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1608910539
transform 1 0 15088 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_187
timestamp 1608910539
transform 1 0 18308 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1608910539
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_177
timestamp 1608910539
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_205
timestamp 1608910539
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20148 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18492 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1608910539
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_216
timestamp 1608910539
transform 1 0 20976 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1608910539
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608910539
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_56
timestamp 1608910539
transform 1 0 6256 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608910539
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1608910539
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1608910539
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8188 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1608910539
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_95
timestamp 1608910539
transform 1 0 9844 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1608910539
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_86
timestamp 1608910539
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_124
timestamp 1608910539
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1608910539
transform 1 0 12236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1608910539
transform 1 0 11868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1608910539
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1608910539
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_140
timestamp 1608910539
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_135
timestamp 1608910539
transform 1 0 13524 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12696 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1608910539
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_157
timestamp 1608910539
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 15364 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_161
timestamp 1608910539
transform 1 0 15916 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15732 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_165
timestamp 1608910539
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 1608910539
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_173
timestamp 1608910539
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_169
timestamp 1608910539
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1608910539
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 17572 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1608910539
transform 1 0 19412 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_195
timestamp 1608910539
transform 1 0 19044 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19504 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1608910539
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1608910539
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1608910539
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608910539
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1608910539
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8740 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7084 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp 1608910539
transform 1 0 9936 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_92
timestamp 1608910539
transform 1 0 9568 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10028 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1608910539
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1608910539
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12512 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608910539
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1608910539
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1608910539
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608910539
transform 1 0 14168 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1608910539
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_159
timestamp 1608910539
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_149
timestamp 1608910539
transform 1 0 14812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 14904 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1608910539
transform 1 0 15916 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1608910539
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_175
timestamp 1608910539
transform 1 0 17204 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1608910539
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608910539
transform 1 0 18308 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_202
timestamp 1608910539
transform 1 0 19688 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_191
timestamp 1608910539
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18860 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 19964 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1608910539
transform 1 0 21344 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_214
timestamp 1608910539
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608910539
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608910539
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608910539
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_56
timestamp 1608910539
transform 1 0 6256 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608910539
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1608910539
transform 1 0 7360 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_80
timestamp 1608910539
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1608910539
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_64
timestamp 1608910539
transform 1 0 6992 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7452 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608910539
transform 1 0 8648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1608910539
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1608910539
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1608910539
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9108 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1608910539
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_96
timestamp 1608910539
transform 1 0 9936 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_95
timestamp 1608910539
transform 1 0 9844 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10120 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1608910539
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1608910539
transform 1 0 11592 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1608910539
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_116
timestamp 1608910539
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1608910539
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12328 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_143
timestamp 1608910539
transform 1 0 14260 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1608910539
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_126
timestamp 1608910539
transform 1 0 12696 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1608910539
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13064 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13984 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_163
timestamp 1608910539
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_163
timestamp 1608910539
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1608910539
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16284 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16376 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14628 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_174
timestamp 1608910539
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_175
timestamp 1608910539
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1608910539
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 17296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1608910539
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_184
timestamp 1608910539
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1608910539
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1608910539
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1608910539
transform 1 0 17756 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_7_200
timestamp 1608910539
transform 1 0 19504 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1608910539
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1608910539
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18768 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19780 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1608910539
transform 1 0 21252 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1608910539
transform 1 0 21252 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1608910539
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608910539
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608910539
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1608910539
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7912 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1608910539
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11316 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_131
timestamp 1608910539
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1608910539
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13340 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1608910539
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1608910539
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16928 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1608910539
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_188
timestamp 1608910539
transform 1 0 18400 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 18768 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1608910539
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1608910539
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1608910539
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608910539
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1608910539
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1608910539
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_82
timestamp 1608910539
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_74
timestamp 1608910539
transform 1 0 7912 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1608910539
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1608910539
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1608910539
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8832 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608910539
transform 1 0 9844 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1608910539
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_112
timestamp 1608910539
transform 1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608910539
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1608910539
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14076 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1608910539
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1608910539
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15824 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15088 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_186
timestamp 1608910539
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1608910539
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1608910539
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16836 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_207
timestamp 1608910539
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1608910539
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_192
timestamp 1608910539
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1608910539
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19320 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1608910539
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_218
timestamp 1608910539
transform 1 0 21160 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 20332 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608910539
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608910539
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608910539
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608910539
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_80
timestamp 1608910539
transform 1 0 8464 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 1608910539
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_95
timestamp 1608910539
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608910539
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_122
timestamp 1608910539
transform 1 0 12328 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_111
timestamp 1608910539
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1608910539
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1608910539
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13984 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12972 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1608910539
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1608910539
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1608910539
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1608910539
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18216 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16560 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_201
timestamp 1608910539
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_195
timestamp 1608910539
transform 1 0 19044 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1608910539
transform 1 0 19320 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1608910539
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1608910539
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1608910539
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608910539
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608910539
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608910539
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608910539
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1608910539
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8096 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1608910539
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9752 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1608910539
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1608910539
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1608910539
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1608910539
transform 1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1608910539
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_128
timestamp 1608910539
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13524 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1608910539
transform 1 0 13064 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_159
timestamp 1608910539
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_155
timestamp 1608910539
transform 1 0 15364 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15824 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_187
timestamp 1608910539
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1608910539
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1608910539
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608910539
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp 1608910539
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1608910539
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19412 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1608910539
transform 1 0 18952 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1608910539
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1608910539
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1608910539
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608910539
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608910539
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1608910539
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608910539
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1608910539
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_96
timestamp 1608910539
transform 1 0 9936 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608910539
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10212 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1608910539
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11868 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1608910539
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1608910539
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_184
timestamp 1608910539
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_179
timestamp 1608910539
transform 1 0 17572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1608910539
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp 1608910539
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18216 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1608910539
transform 1 0 16928 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1608910539
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_195
timestamp 1608910539
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1608910539
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1608910539
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1608910539
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608910539
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608910539
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608910539
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1608910539
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1608910539
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1608910539
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1608910539
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608910539
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1608910539
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1608910539
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1608910539
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_98
timestamp 1608910539
transform 1 0 10120 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1608910539
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1608910539
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1608910539
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1608910539
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1608910539
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_106
timestamp 1608910539
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11040 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1608910539
transform 1 0 12972 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 1608910539
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13340 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1608910539
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_139
timestamp 1608910539
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_137
timestamp 1608910539
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13892 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608910539
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1608910539
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1608910539
transform 1 0 15364 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_164
timestamp 1608910539
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_160
timestamp 1608910539
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_156
timestamp 1608910539
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15732 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 16376 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1608910539
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1608910539
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1608910539
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_168
timestamp 1608910539
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1608910539
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_184
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608910539
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1608910539
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18308 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16836 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_202
timestamp 1608910539
transform 1 0 19688 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_198
timestamp 1608910539
transform 1 0 19320 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1608910539
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18492 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19964 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1608910539
transform 1 0 21252 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1608910539
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1608910539
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608910539
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1608910539
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1608910539
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1608910539
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1608910539
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1608910539
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1608910539
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_123
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1608910539
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12512 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1608910539
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14168 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1608910539
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15824 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1608910539
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1608910539
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16836 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1608910539
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19688 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_222
timestamp 1608910539
transform 1 0 21528 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_218
timestamp 1608910539
transform 1 0 21160 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608910539
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608910539
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1608910539
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1608910539
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1608910539
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_117
timestamp 1608910539
transform 1 0 11868 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1608910539
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12144 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1608910539
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_132
timestamp 1608910539
transform 1 0 13248 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_126
timestamp 1608910539
transform 1 0 12696 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608910539
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_147
timestamp 1608910539
transform 1 0 14628 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1608910539
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16928 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1608910539
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_188
timestamp 1608910539
transform 1 0 18400 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18768 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1608910539
transform 1 0 21252 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1608910539
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608910539
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1608910539
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1608910539
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1608910539
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1608910539
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1608910539
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1608910539
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1608910539
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1608910539
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_154
timestamp 1608910539
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1608910539
transform 1 0 14628 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15456 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608910539
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_187
timestamp 1608910539
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1608910539
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1608910539
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1608910539
transform 1 0 18124 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17112 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_191
timestamp 1608910539
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18860 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1608910539
transform 1 0 21528 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_218
timestamp 1608910539
transform 1 0 21160 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_213
timestamp 1608910539
transform 1 0 20700 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1608910539
transform 1 0 20332 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1608910539
transform 1 0 20792 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608910539
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608910539
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1608910539
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1608910539
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1608910539
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1608910539
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1608910539
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1608910539
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1608910539
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1608910539
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1608910539
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1608910539
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17848 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_204
timestamp 1608910539
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_198
timestamp 1608910539
transform 1 0 19320 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1608910539
transform 1 0 19596 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1608910539
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608910539
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608910539
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608910539
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608910539
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608910539
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608910539
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608910539
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1608910539
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1608910539
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608910539
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608910539
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1608910539
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608910539
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608910539
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13524 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1608910539
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1608910539
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16192 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1608910539
transform 1 0 18032 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1608910539
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_187
timestamp 1608910539
transform 1 0 18308 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1608910539
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1608910539
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_196
timestamp 1608910539
transform 1 0 19136 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1608910539
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1608910539
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_195
timestamp 1608910539
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1608910539
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19596 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608910539
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608910539
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_215
timestamp 1608910539
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20332 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1608910539
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1608910539
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608910539
transform 1 0 21068 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608910539
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1608910539
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1608910539
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608910539
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1608910539
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1608910539
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_98
timestamp 1608910539
transform 1 0 10120 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1608910539
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1608910539
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1608910539
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_106
timestamp 1608910539
transform 1 0 10856 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11132 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1608910539
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1608910539
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1608910539
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_204
timestamp 1608910539
transform 1 0 19872 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_196
timestamp 1608910539
transform 1 0 19136 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20148 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1608910539
transform 1 0 21252 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608910539
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608910539
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1608910539
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608910539
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_80
timestamp 1608910539
transform 1 0 8464 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1608910539
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8740 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1608910539
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1608910539
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1608910539
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1608910539
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_135
timestamp 1608910539
transform 1 0 13524 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1608910539
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1608910539
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1608910539
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1608910539
transform 1 0 19688 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1608910539
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1608910539
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608910539
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1608910539
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1608910539
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1608910539
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1608910539
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1608910539
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1608910539
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1608910539
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1608910539
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_110
timestamp 1608910539
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11592 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1608910539
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1608910539
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1608910539
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1608910539
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_208
timestamp 1608910539
transform 1 0 20240 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1608910539
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1608910539
transform 1 0 21528 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1608910539
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608910539
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1608910539
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1608910539
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1608910539
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1608910539
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1608910539
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1608910539
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1608910539
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1608910539
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1608910539
transform 1 0 14076 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1608910539
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14352 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1608910539
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1608910539
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1608910539
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_202
timestamp 1608910539
transform 1 0 19688 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1608910539
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608910539
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1608910539
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1608910539
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1608910539
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1608910539
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1608910539
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608910539
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1608910539
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1608910539
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1608910539
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1608910539
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1608910539
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1608910539
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1608910539
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1608910539
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1608910539
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1608910539
transform 1 0 19136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1608910539
transform 1 0 21528 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1608910539
transform 1 0 21160 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_210
timestamp 1608910539
transform 1 0 20424 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608910539
transform 1 0 20792 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1608910539
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1608910539
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1608910539
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1608910539
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608910539
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1608910539
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1608910539
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1608910539
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1608910539
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1608910539
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1608910539
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1608910539
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1608910539
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1608910539
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_116
timestamp 1608910539
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1608910539
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1608910539
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11224 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1608910539
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1608910539
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1608910539
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1608910539
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1608910539
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1608910539
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1608910539
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_186
timestamp 1608910539
transform 1 0 18216 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_178
timestamp 1608910539
transform 1 0 17480 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17664 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_202
timestamp 1608910539
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_194
timestamp 1608910539
transform 1 0 18952 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_198
timestamp 1608910539
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608910539
transform 1 0 18584 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1608910539
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1608910539
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_218
timestamp 1608910539
transform 1 0 21160 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608910539
transform 1 0 20792 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1608910539
transform 1 0 21528 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1608910539
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1608910539
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1608910539
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1608910539
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1608910539
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1608910539
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_68
timestamp 1608910539
transform 1 0 7360 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8280 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1608910539
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1608910539
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1608910539
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1608910539
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1608910539
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1608910539
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1608910539
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1608910539
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1608910539
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1608910539
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1608910539
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1608910539
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1608910539
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608910539
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1608910539
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1608910539
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_96
timestamp 1608910539
transform 1 0 9936 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_86
timestamp 1608910539
transform 1 0 9016 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9384 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1608910539
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_108
timestamp 1608910539
transform 1 0 11040 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1608910539
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1608910539
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1608910539
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1608910539
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_208
timestamp 1608910539
transform 1 0 20240 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1608910539
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1608910539
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_218
timestamp 1608910539
transform 1 0 21160 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608910539
transform 1 0 20792 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1608910539
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608910539
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1608910539
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1608910539
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1608910539
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1608910539
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_125
timestamp 1608910539
transform 1 0 12604 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_117
timestamp 1608910539
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1608910539
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12052 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_137
timestamp 1608910539
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1608910539
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_154
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1608910539
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15824 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_178
timestamp 1608910539
transform 1 0 17480 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18216 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_192
timestamp 1608910539
transform 1 0 18768 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1608910539
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1608910539
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1608910539
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1608910539
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1608910539
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608910539
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1608910539
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1608910539
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1608910539
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1608910539
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1608910539
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1608910539
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1608910539
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_106
timestamp 1608910539
transform 1 0 10856 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1608910539
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1608910539
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1608910539
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1608910539
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1608910539
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_196
timestamp 1608910539
transform 1 0 19136 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 19688 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608910539
transform 1 0 20240 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1608910539
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1608910539
transform 1 0 21160 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1608910539
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608910539
transform 1 0 20792 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608910539
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608910539
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1608910539
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608910539
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1608910539
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1608910539
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1608910539
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1608910539
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1608910539
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1608910539
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1608910539
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1608910539
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_202
timestamp 1608910539
transform 1 0 19688 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1608910539
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 20240 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1608910539
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1608910539
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1608910539
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1608910539
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1608910539
transform 1 0 6256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1608910539
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_75
timestamp 1608910539
transform 1 0 8004 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_87
timestamp 1608910539
transform 1 0 9108 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1608910539
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_199
timestamp 1608910539
transform 1 0 19412 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1608910539
transform 1 0 21528 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_211
timestamp 1608910539
transform 1 0 20516 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5722 22200 5778 23000 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_1_
port 2 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 ccff_tail
port 4 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 5 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[10]
port 6 nsew signal input
rlabel metal3 s 22200 8848 23000 8968 6 chanx_right_in[11]
port 7 nsew signal input
rlabel metal3 s 22200 9256 23000 9376 6 chanx_right_in[12]
port 8 nsew signal input
rlabel metal3 s 22200 9664 23000 9784 6 chanx_right_in[13]
port 9 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[14]
port 10 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[15]
port 11 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[16]
port 12 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[17]
port 13 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[18]
port 14 nsew signal input
rlabel metal3 s 22200 12520 23000 12640 6 chanx_right_in[19]
port 15 nsew signal input
rlabel metal3 s 22200 4224 23000 4344 6 chanx_right_in[1]
port 16 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[2]
port 17 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 18 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[4]
port 19 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[5]
port 20 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[6]
port 21 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[7]
port 22 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[8]
port 23 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[9]
port 24 nsew signal input
rlabel metal3 s 22200 12928 23000 13048 6 chanx_right_out[0]
port 25 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[10]
port 26 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[11]
port 27 nsew signal tristate
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[12]
port 28 nsew signal tristate
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[13]
port 29 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[14]
port 30 nsew signal tristate
rlabel metal3 s 22200 19864 23000 19984 6 chanx_right_out[15]
port 31 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[16]
port 32 nsew signal tristate
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[17]
port 33 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[18]
port 34 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[19]
port 35 nsew signal tristate
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[1]
port 36 nsew signal tristate
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[2]
port 37 nsew signal tristate
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[3]
port 38 nsew signal tristate
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[4]
port 39 nsew signal tristate
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[5]
port 40 nsew signal tristate
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[6]
port 41 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[7]
port 42 nsew signal tristate
rlabel metal3 s 22200 16600 23000 16720 6 chanx_right_out[8]
port 43 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[9]
port 44 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 chany_bottom_in[0]
port 45 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_in[10]
port 46 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_in[11]
port 47 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[12]
port 48 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[13]
port 49 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 chany_bottom_in[14]
port 50 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[15]
port 51 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[16]
port 52 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[17]
port 53 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[18]
port 54 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 chany_bottom_in[19]
port 55 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 chany_bottom_in[1]
port 56 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_in[2]
port 57 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_in[3]
port 58 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 chany_bottom_in[4]
port 59 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_in[5]
port 60 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_in[6]
port 61 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_in[7]
port 62 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[8]
port 63 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_in[9]
port 64 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_out[0]
port 65 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 chany_bottom_out[10]
port 66 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[11]
port 67 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[12]
port 68 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[13]
port 69 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[14]
port 70 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[15]
port 71 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[16]
port 72 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[17]
port 73 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[18]
port 74 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[19]
port 75 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_out[1]
port 76 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[2]
port 77 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[3]
port 78 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_out[4]
port 79 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[5]
port 80 nsew signal tristate
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_out[6]
port 81 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[7]
port 82 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[8]
port 83 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[9]
port 84 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 prog_clk_0_E_in
port 85 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 86 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 87 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 88 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 89 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 90 nsew signal input
rlabel metal3 s 22200 2320 23000 2440 6 right_bottom_grid_pin_39_
port 91 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 92 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_41_
port 93 nsew signal input
rlabel metal3 s 22200 22584 23000 22704 6 right_top_grid_pin_1_
port 94 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 95 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 96 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 97 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 98 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 99 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
