magic
tech sky130A
magscale 1 2
timestamp 1608762545
<< checkpaint >>
rect -1260 -1260 24060 24060
<< locali >>
rect 9413 18751 9447 18921
rect 12265 16983 12299 17289
rect 9505 13175 9539 13481
rect 12265 13175 12299 13481
rect 15117 13243 15151 13481
rect 13461 9979 13495 10149
rect 13921 6103 13955 6205
rect 19073 5559 19107 5797
rect 10241 4607 10275 4709
<< viali >>
rect 13461 20009 13495 20043
rect 15669 20009 15703 20043
rect 16037 20009 16071 20043
rect 7205 19941 7239 19975
rect 19625 19941 19659 19975
rect 20729 19941 20763 19975
rect 3617 19873 3651 19907
rect 4528 19873 4562 19907
rect 6929 19873 6963 19907
rect 7941 19873 7975 19907
rect 8033 19873 8067 19907
rect 13277 19873 13311 19907
rect 15485 19873 15519 19907
rect 15853 19873 15887 19907
rect 18337 19873 18371 19907
rect 19349 19873 19383 19907
rect 19901 19873 19935 19907
rect 20453 19873 20487 19907
rect 4261 19805 4295 19839
rect 8125 19805 8159 19839
rect 18521 19805 18555 19839
rect 20177 19805 20211 19839
rect 3801 19669 3835 19703
rect 5641 19669 5675 19703
rect 7573 19669 7607 19703
rect 6285 19465 6319 19499
rect 3801 19329 3835 19363
rect 4721 19329 4755 19363
rect 9229 19329 9263 19363
rect 9873 19329 9907 19363
rect 12817 19329 12851 19363
rect 16129 19329 16163 19363
rect 4445 19261 4479 19295
rect 4537 19261 4571 19295
rect 4905 19261 4939 19295
rect 6929 19261 6963 19295
rect 9597 19261 9631 19295
rect 10149 19261 10183 19295
rect 10517 19261 10551 19295
rect 11437 19261 11471 19295
rect 11805 19261 11839 19295
rect 12541 19261 12575 19295
rect 13093 19261 13127 19295
rect 13461 19261 13495 19295
rect 13829 19261 13863 19295
rect 14197 19261 14231 19295
rect 14565 19261 14599 19295
rect 14933 19261 14967 19295
rect 15301 19261 15335 19295
rect 15945 19261 15979 19295
rect 16497 19261 16531 19295
rect 16865 19261 16899 19295
rect 17417 19261 17451 19295
rect 17693 19261 17727 19295
rect 18337 19261 18371 19295
rect 19073 19261 19107 19295
rect 20453 19261 20487 19295
rect 20729 19261 20763 19295
rect 3525 19193 3559 19227
rect 3617 19193 3651 19227
rect 5172 19193 5206 19227
rect 7196 19193 7230 19227
rect 9045 19193 9079 19227
rect 17141 19193 17175 19227
rect 18613 19193 18647 19227
rect 19717 19193 19751 19227
rect 3157 19125 3191 19159
rect 4077 19125 4111 19159
rect 8309 19125 8343 19159
rect 8585 19125 8619 19159
rect 8953 19125 8987 19159
rect 10333 19125 10367 19159
rect 10701 19125 10735 19159
rect 11621 19125 11655 19159
rect 11989 19125 12023 19159
rect 13277 19125 13311 19159
rect 13645 19125 13679 19159
rect 14013 19125 14047 19159
rect 14381 19125 14415 19159
rect 14749 19125 14783 19159
rect 15117 19125 15151 19159
rect 15485 19125 15519 19159
rect 16681 19125 16715 19159
rect 3249 18921 3283 18955
rect 4537 18921 4571 18955
rect 5457 18921 5491 18955
rect 5825 18921 5859 18955
rect 9413 18921 9447 18955
rect 16773 18921 16807 18955
rect 5181 18853 5215 18887
rect 3157 18785 3191 18819
rect 4445 18785 4479 18819
rect 4905 18785 4939 18819
rect 6285 18785 6319 18819
rect 6552 18785 6586 18819
rect 8208 18785 8242 18819
rect 10885 18853 10919 18887
rect 14565 18853 14599 18887
rect 15577 18853 15611 18887
rect 20545 18853 20579 18887
rect 10057 18785 10091 18819
rect 10609 18785 10643 18819
rect 11612 18785 11646 18819
rect 13084 18785 13118 18819
rect 14289 18785 14323 18819
rect 15301 18785 15335 18819
rect 16589 18785 16623 18819
rect 17969 18785 18003 18819
rect 18521 18785 18555 18819
rect 19165 18785 19199 18819
rect 19717 18785 19751 18819
rect 20269 18785 20303 18819
rect 3387 18717 3421 18751
rect 4721 18717 4755 18751
rect 5917 18717 5951 18751
rect 6101 18717 6135 18751
rect 7941 18717 7975 18751
rect 9413 18717 9447 18751
rect 10149 18717 10183 18751
rect 10241 18717 10275 18751
rect 11345 18717 11379 18751
rect 12817 18717 12851 18751
rect 18153 18717 18187 18751
rect 18705 18717 18739 18751
rect 19349 18717 19383 18751
rect 19901 18717 19935 18751
rect 12725 18649 12759 18683
rect 2789 18581 2823 18615
rect 4077 18581 4111 18615
rect 7665 18581 7699 18615
rect 9321 18581 9355 18615
rect 9689 18581 9723 18615
rect 14197 18581 14231 18615
rect 2145 18377 2179 18411
rect 4445 18377 4479 18411
rect 7297 18377 7331 18411
rect 9229 18377 9263 18411
rect 12449 18377 12483 18411
rect 13277 18377 13311 18411
rect 17233 18377 17267 18411
rect 1961 18309 1995 18343
rect 4353 18309 4387 18343
rect 2697 18241 2731 18275
rect 4905 18241 4939 18275
rect 4997 18241 5031 18275
rect 6285 18241 6319 18275
rect 7849 18241 7883 18275
rect 8585 18241 8619 18275
rect 8677 18241 8711 18275
rect 9873 18241 9907 18275
rect 13093 18241 13127 18275
rect 13829 18241 13863 18275
rect 19625 18241 19659 18275
rect 20729 18241 20763 18275
rect 1777 18173 1811 18207
rect 2513 18173 2547 18207
rect 2973 18173 3007 18207
rect 6101 18173 6135 18207
rect 8493 18173 8527 18207
rect 9597 18173 9631 18207
rect 10241 18173 10275 18207
rect 12909 18173 12943 18207
rect 13737 18173 13771 18207
rect 17049 18173 17083 18207
rect 19349 18173 19383 18207
rect 19901 18173 19935 18207
rect 20453 18173 20487 18207
rect 2605 18105 2639 18139
rect 3240 18105 3274 18139
rect 6009 18105 6043 18139
rect 7665 18105 7699 18139
rect 10508 18105 10542 18139
rect 13645 18105 13679 18139
rect 20177 18105 20211 18139
rect 4813 18037 4847 18071
rect 5641 18037 5675 18071
rect 7757 18037 7791 18071
rect 8125 18037 8159 18071
rect 9689 18037 9723 18071
rect 11621 18037 11655 18071
rect 12817 18037 12851 18071
rect 1685 17833 1719 17867
rect 6469 17833 6503 17867
rect 7205 17833 7239 17867
rect 8033 17833 8067 17867
rect 10977 17833 11011 17867
rect 11437 17833 11471 17867
rect 13001 17833 13035 17867
rect 21097 17833 21131 17867
rect 2136 17765 2170 17799
rect 4782 17765 4816 17799
rect 6377 17765 6411 17799
rect 13093 17765 13127 17799
rect 1501 17697 1535 17731
rect 1869 17697 1903 17731
rect 7573 17697 7607 17731
rect 8401 17697 8435 17731
rect 10517 17697 10551 17731
rect 11345 17697 11379 17731
rect 12173 17697 12207 17731
rect 13728 17697 13762 17731
rect 20269 17697 20303 17731
rect 20913 17697 20947 17731
rect 4537 17629 4571 17663
rect 6561 17629 6595 17663
rect 7665 17629 7699 17663
rect 7849 17629 7883 17663
rect 8493 17629 8527 17663
rect 8677 17629 8711 17663
rect 10609 17629 10643 17663
rect 10793 17629 10827 17663
rect 11529 17629 11563 17663
rect 12265 17629 12299 17663
rect 12357 17629 12391 17663
rect 13277 17629 13311 17663
rect 13461 17629 13495 17663
rect 20545 17629 20579 17663
rect 10149 17561 10183 17595
rect 3249 17493 3283 17527
rect 5917 17493 5951 17527
rect 6009 17493 6043 17527
rect 11805 17493 11839 17527
rect 12633 17493 12667 17527
rect 14841 17493 14875 17527
rect 1961 17289 1995 17323
rect 4629 17289 4663 17323
rect 6837 17289 6871 17323
rect 8401 17289 8435 17323
rect 10977 17289 11011 17323
rect 11437 17289 11471 17323
rect 12265 17289 12299 17323
rect 19901 17289 19935 17323
rect 20269 17289 20303 17323
rect 21189 17289 21223 17323
rect 2145 17221 2179 17255
rect 2697 17153 2731 17187
rect 3525 17153 3559 17187
rect 4353 17153 4387 17187
rect 5181 17153 5215 17187
rect 6009 17153 6043 17187
rect 6101 17153 6135 17187
rect 7481 17153 7515 17187
rect 8125 17153 8159 17187
rect 9045 17153 9079 17187
rect 9597 17153 9631 17187
rect 11897 17153 11931 17187
rect 11989 17153 12023 17187
rect 1777 17085 1811 17119
rect 2605 17085 2639 17119
rect 4997 17085 5031 17119
rect 5917 17085 5951 17119
rect 9864 17085 9898 17119
rect 11161 17085 11195 17119
rect 2513 17017 2547 17051
rect 3433 17017 3467 17051
rect 4169 17017 4203 17051
rect 5089 17017 5123 17051
rect 7297 17017 7331 17051
rect 11805 17017 11839 17051
rect 12449 17221 12483 17255
rect 12909 17153 12943 17187
rect 13093 17153 13127 17187
rect 12817 17085 12851 17119
rect 13277 17085 13311 17119
rect 14749 17085 14783 17119
rect 19717 17085 19751 17119
rect 20085 17085 20119 17119
rect 20453 17085 20487 17119
rect 21005 17085 21039 17119
rect 13544 17017 13578 17051
rect 14994 17017 15028 17051
rect 20729 17017 20763 17051
rect 2973 16949 3007 16983
rect 3341 16949 3375 16983
rect 3801 16949 3835 16983
rect 4261 16949 4295 16983
rect 5549 16949 5583 16983
rect 7205 16949 7239 16983
rect 8769 16949 8803 16983
rect 8861 16949 8895 16983
rect 12265 16949 12299 16983
rect 14657 16949 14691 16983
rect 16129 16949 16163 16983
rect 1593 16745 1627 16779
rect 1777 16745 1811 16779
rect 2145 16745 2179 16779
rect 2605 16745 2639 16779
rect 3617 16745 3651 16779
rect 4537 16745 4571 16779
rect 5733 16745 5767 16779
rect 6193 16745 6227 16779
rect 6653 16745 6687 16779
rect 8677 16745 8711 16779
rect 10057 16745 10091 16779
rect 10885 16745 10919 16779
rect 11713 16745 11747 16779
rect 12081 16745 12115 16779
rect 12633 16745 12667 16779
rect 13093 16745 13127 16779
rect 13461 16745 13495 16779
rect 14749 16745 14783 16779
rect 16957 16745 16991 16779
rect 21097 16745 21131 16779
rect 2237 16677 2271 16711
rect 4905 16677 4939 16711
rect 9045 16677 9079 16711
rect 13001 16677 13035 16711
rect 15546 16677 15580 16711
rect 1409 16609 1443 16643
rect 2973 16609 3007 16643
rect 3433 16609 3467 16643
rect 5825 16609 5859 16643
rect 6561 16609 6595 16643
rect 7205 16609 7239 16643
rect 7472 16609 7506 16643
rect 11253 16609 11287 16643
rect 11345 16609 11379 16643
rect 12173 16609 12207 16643
rect 13829 16609 13863 16643
rect 14657 16609 14691 16643
rect 15301 16609 15335 16643
rect 16773 16609 16807 16643
rect 20269 16609 20303 16643
rect 20545 16609 20579 16643
rect 20913 16609 20947 16643
rect 2421 16541 2455 16575
rect 3065 16541 3099 16575
rect 3249 16541 3283 16575
rect 4997 16541 5031 16575
rect 5089 16541 5123 16575
rect 5917 16541 5951 16575
rect 6745 16541 6779 16575
rect 9137 16541 9171 16575
rect 9229 16541 9263 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 11529 16541 11563 16575
rect 12265 16541 12299 16575
rect 13185 16541 13219 16575
rect 13921 16541 13955 16575
rect 14105 16541 14139 16575
rect 14841 16541 14875 16575
rect 8585 16473 8619 16507
rect 9689 16473 9723 16507
rect 16681 16473 16715 16507
rect 5365 16405 5399 16439
rect 14289 16405 14323 16439
rect 1593 16201 1627 16235
rect 3709 16201 3743 16235
rect 4445 16201 4479 16235
rect 8217 16201 8251 16235
rect 8861 16201 8895 16235
rect 12265 16201 12299 16235
rect 13093 16201 13127 16235
rect 13921 16201 13955 16235
rect 14749 16201 14783 16235
rect 18245 16201 18279 16235
rect 20361 16201 20395 16235
rect 20729 16201 20763 16235
rect 1961 16133 1995 16167
rect 4997 16065 5031 16099
rect 9413 16065 9447 16099
rect 10517 16065 10551 16099
rect 10885 16065 10919 16099
rect 13553 16065 13587 16099
rect 13737 16065 13771 16099
rect 14473 16065 14507 16099
rect 15301 16065 15335 16099
rect 16957 16065 16991 16099
rect 19809 16065 19843 16099
rect 1409 15997 1443 16031
rect 1777 15997 1811 16031
rect 2329 15997 2363 16031
rect 2596 15997 2630 16031
rect 5273 15997 5307 16031
rect 6837 15997 6871 16031
rect 9229 15997 9263 16031
rect 15209 15997 15243 16031
rect 18061 15997 18095 16031
rect 19533 15997 19567 16031
rect 20177 15997 20211 16031
rect 20545 15997 20579 16031
rect 20913 15997 20947 16031
rect 4353 15929 4387 15963
rect 5540 15929 5574 15963
rect 7082 15929 7116 15963
rect 9321 15929 9355 15963
rect 10333 15929 10367 15963
rect 11152 15929 11186 15963
rect 14289 15929 14323 15963
rect 16773 15929 16807 15963
rect 4813 15861 4847 15895
rect 4905 15861 4939 15895
rect 6653 15861 6687 15895
rect 8677 15861 8711 15895
rect 9965 15861 9999 15895
rect 10425 15861 10459 15895
rect 13461 15861 13495 15895
rect 14381 15861 14415 15895
rect 15117 15861 15151 15895
rect 16405 15861 16439 15895
rect 16865 15861 16899 15895
rect 17233 15861 17267 15895
rect 21097 15861 21131 15895
rect 2053 15657 2087 15691
rect 2881 15657 2915 15691
rect 3341 15657 3375 15691
rect 6837 15657 6871 15691
rect 8769 15657 8803 15691
rect 9137 15657 9171 15691
rect 12081 15657 12115 15691
rect 12449 15657 12483 15691
rect 13369 15657 13403 15691
rect 13737 15657 13771 15691
rect 14197 15657 14231 15691
rect 15301 15657 15335 15691
rect 18061 15657 18095 15691
rect 18153 15657 18187 15691
rect 20269 15657 20303 15691
rect 1777 15589 1811 15623
rect 2421 15589 2455 15623
rect 3709 15589 3743 15623
rect 6377 15589 6411 15623
rect 1501 15521 1535 15555
rect 3249 15521 3283 15555
rect 4712 15521 4746 15555
rect 7205 15521 7239 15555
rect 7297 15521 7331 15555
rect 9229 15521 9263 15555
rect 10140 15521 10174 15555
rect 14565 15521 14599 15555
rect 16488 15521 16522 15555
rect 18521 15521 18555 15555
rect 20085 15521 20119 15555
rect 20453 15521 20487 15555
rect 20913 15521 20947 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 3433 15453 3467 15487
rect 4445 15453 4479 15487
rect 6469 15453 6503 15487
rect 6653 15453 6687 15487
rect 7481 15453 7515 15487
rect 7665 15453 7699 15487
rect 9413 15453 9447 15487
rect 9873 15453 9907 15487
rect 12541 15453 12575 15487
rect 12633 15453 12667 15487
rect 13829 15453 13863 15487
rect 14013 15453 14047 15487
rect 14657 15453 14691 15487
rect 14749 15453 14783 15487
rect 16221 15453 16255 15487
rect 18245 15453 18279 15487
rect 18797 15453 18831 15487
rect 6009 15385 6043 15419
rect 17601 15385 17635 15419
rect 5825 15317 5859 15351
rect 11253 15317 11287 15351
rect 17693 15317 17727 15351
rect 20637 15317 20671 15351
rect 21097 15317 21131 15351
rect 1593 15113 1627 15147
rect 2697 15113 2731 15147
rect 3065 15113 3099 15147
rect 7205 15113 7239 15147
rect 8033 15113 8067 15147
rect 11529 15113 11563 15147
rect 17049 15113 17083 15147
rect 18061 15113 18095 15147
rect 19625 15113 19659 15147
rect 10241 15045 10275 15079
rect 12725 15045 12759 15079
rect 21097 15045 21131 15079
rect 4077 14977 4111 15011
rect 4813 14977 4847 15011
rect 5917 14977 5951 15011
rect 7757 14977 7791 15011
rect 8493 14977 8527 15011
rect 8585 14977 8619 15011
rect 8861 14977 8895 15011
rect 11345 14977 11379 15011
rect 12081 14977 12115 15011
rect 13369 14977 13403 15011
rect 14197 14977 14231 15011
rect 15577 14977 15611 15011
rect 17693 14977 17727 15011
rect 18613 14977 18647 15011
rect 1409 14909 1443 14943
rect 1777 14909 1811 14943
rect 2145 14909 2179 14943
rect 2513 14909 2547 14943
rect 2881 14909 2915 14943
rect 7573 14909 7607 14943
rect 7665 14909 7699 14943
rect 8401 14909 8435 14943
rect 15844 14909 15878 14943
rect 17509 14909 17543 14943
rect 18429 14909 18463 14943
rect 19441 14909 19475 14943
rect 19809 14909 19843 14943
rect 20177 14909 20211 14943
rect 20545 14909 20579 14943
rect 20913 14909 20947 14943
rect 4629 14841 4663 14875
rect 9128 14841 9162 14875
rect 13093 14841 13127 14875
rect 17417 14841 17451 14875
rect 1961 14773 1995 14807
rect 2329 14773 2363 14807
rect 3433 14773 3467 14807
rect 3801 14773 3835 14807
rect 3893 14773 3927 14807
rect 4261 14773 4295 14807
rect 4721 14773 4755 14807
rect 5365 14773 5399 14807
rect 5733 14773 5767 14807
rect 5825 14773 5859 14807
rect 10701 14773 10735 14807
rect 11069 14773 11103 14807
rect 11161 14773 11195 14807
rect 11897 14773 11931 14807
rect 11989 14773 12023 14807
rect 13185 14773 13219 14807
rect 13553 14773 13587 14807
rect 13921 14773 13955 14807
rect 14013 14773 14047 14807
rect 16957 14773 16991 14807
rect 18521 14773 18555 14807
rect 19993 14773 20027 14807
rect 20361 14773 20395 14807
rect 20729 14773 20763 14807
rect 3157 14569 3191 14603
rect 5457 14569 5491 14603
rect 6009 14569 6043 14603
rect 6837 14569 6871 14603
rect 7665 14569 7699 14603
rect 9965 14569 9999 14603
rect 10333 14569 10367 14603
rect 10793 14569 10827 14603
rect 11621 14569 11655 14603
rect 13921 14569 13955 14603
rect 14841 14569 14875 14603
rect 15761 14569 15795 14603
rect 2237 14501 2271 14535
rect 4344 14501 4378 14535
rect 6377 14501 6411 14535
rect 17500 14501 17534 14535
rect 19901 14501 19935 14535
rect 20453 14501 20487 14535
rect 1593 14433 1627 14467
rect 1961 14433 1995 14467
rect 2513 14433 2547 14467
rect 3525 14433 3559 14467
rect 7205 14433 7239 14467
rect 7849 14433 7883 14467
rect 7948 14433 7982 14467
rect 8208 14433 8242 14467
rect 11161 14433 11195 14467
rect 11989 14433 12023 14467
rect 12541 14433 12575 14467
rect 12808 14433 12842 14467
rect 14197 14433 14231 14467
rect 14749 14433 14783 14467
rect 16129 14433 16163 14467
rect 19625 14433 19659 14467
rect 20177 14433 20211 14467
rect 20913 14433 20947 14467
rect 3617 14365 3651 14399
rect 3801 14365 3835 14399
rect 4077 14365 4111 14399
rect 6469 14365 6503 14399
rect 6561 14365 6595 14399
rect 7297 14365 7331 14399
rect 7481 14365 7515 14399
rect 10425 14365 10459 14399
rect 10609 14365 10643 14399
rect 11253 14365 11287 14399
rect 11345 14365 11379 14399
rect 12081 14365 12115 14399
rect 12173 14365 12207 14399
rect 15025 14365 15059 14399
rect 16221 14365 16255 14399
rect 16405 14365 16439 14399
rect 17233 14365 17267 14399
rect 9321 14297 9355 14331
rect 14381 14297 14415 14331
rect 1777 14229 1811 14263
rect 2697 14229 2731 14263
rect 14013 14229 14047 14263
rect 18613 14229 18647 14263
rect 21097 14229 21131 14263
rect 4169 14025 4203 14059
rect 5917 14025 5951 14059
rect 9505 14025 9539 14059
rect 11529 14025 11563 14059
rect 16773 14025 16807 14059
rect 18061 14025 18095 14059
rect 19717 14025 19751 14059
rect 6009 13957 6043 13991
rect 17049 13957 17083 13991
rect 10057 13889 10091 13923
rect 10977 13889 11011 13923
rect 11161 13889 11195 13923
rect 12173 13889 12207 13923
rect 15393 13889 15427 13923
rect 17693 13889 17727 13923
rect 18613 13889 18647 13923
rect 19441 13889 19475 13923
rect 20177 13889 20211 13923
rect 20361 13889 20395 13923
rect 20729 13889 20763 13923
rect 1593 13821 1627 13855
rect 1961 13821 1995 13855
rect 2237 13821 2271 13855
rect 2789 13821 2823 13855
rect 4537 13821 4571 13855
rect 6193 13821 6227 13855
rect 6837 13821 6871 13855
rect 7104 13821 7138 13855
rect 9965 13821 9999 13855
rect 12449 13821 12483 13855
rect 13921 13821 13955 13855
rect 14177 13821 14211 13855
rect 15660 13821 15694 13855
rect 20545 13821 20579 13855
rect 3056 13753 3090 13787
rect 4804 13753 4838 13787
rect 9873 13753 9907 13787
rect 11989 13753 12023 13787
rect 12716 13753 12750 13787
rect 17417 13753 17451 13787
rect 18429 13753 18463 13787
rect 19257 13753 19291 13787
rect 20085 13753 20119 13787
rect 1777 13685 1811 13719
rect 8217 13685 8251 13719
rect 10333 13685 10367 13719
rect 10701 13685 10735 13719
rect 10793 13685 10827 13719
rect 11897 13685 11931 13719
rect 13829 13685 13863 13719
rect 15301 13685 15335 13719
rect 17509 13685 17543 13719
rect 18521 13685 18555 13719
rect 18889 13685 18923 13719
rect 19349 13685 19383 13719
rect 2973 13481 3007 13515
rect 4077 13481 4111 13515
rect 4905 13481 4939 13515
rect 5733 13481 5767 13515
rect 6561 13481 6595 13515
rect 8309 13481 8343 13515
rect 8677 13481 8711 13515
rect 9045 13481 9079 13515
rect 9505 13481 9539 13515
rect 1869 13413 1903 13447
rect 4537 13413 4571 13447
rect 9137 13413 9171 13447
rect 1593 13345 1627 13379
rect 2513 13345 2547 13379
rect 3341 13345 3375 13379
rect 4445 13345 4479 13379
rect 5273 13345 5307 13379
rect 6101 13345 6135 13379
rect 6193 13345 6227 13379
rect 6929 13345 6963 13379
rect 8217 13345 8251 13379
rect 2605 13277 2639 13311
rect 2789 13277 2823 13311
rect 3433 13277 3467 13311
rect 3617 13277 3651 13311
rect 4629 13277 4663 13311
rect 5365 13277 5399 13311
rect 5457 13277 5491 13311
rect 6377 13277 6411 13311
rect 7021 13277 7055 13311
rect 7205 13277 7239 13311
rect 8401 13277 8435 13311
rect 9229 13277 9263 13311
rect 12265 13481 12299 13515
rect 13093 13481 13127 13515
rect 13461 13481 13495 13515
rect 13829 13481 13863 13515
rect 14289 13481 14323 13515
rect 14749 13481 14783 13515
rect 15117 13481 15151 13515
rect 15301 13481 15335 13515
rect 16957 13481 16991 13515
rect 19073 13481 19107 13515
rect 11069 13345 11103 13379
rect 11161 13277 11195 13311
rect 11345 13277 11379 13311
rect 10701 13209 10735 13243
rect 2145 13141 2179 13175
rect 7849 13141 7883 13175
rect 9505 13141 9539 13175
rect 13001 13345 13035 13379
rect 13921 13345 13955 13379
rect 14657 13345 14691 13379
rect 12541 13277 12575 13311
rect 13185 13277 13219 13311
rect 14013 13277 14047 13311
rect 14933 13277 14967 13311
rect 16497 13413 16531 13447
rect 19410 13413 19444 13447
rect 15669 13345 15703 13379
rect 17141 13345 17175 13379
rect 17693 13345 17727 13379
rect 17960 13345 17994 13379
rect 19165 13345 19199 13379
rect 20913 13345 20947 13379
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 16589 13277 16623 13311
rect 16681 13277 16715 13311
rect 12633 13209 12667 13243
rect 15117 13209 15151 13243
rect 16129 13209 16163 13243
rect 12265 13141 12299 13175
rect 20545 13141 20579 13175
rect 21097 13141 21131 13175
rect 1777 12937 1811 12971
rect 1961 12937 1995 12971
rect 5273 12937 5307 12971
rect 6837 12937 6871 12971
rect 7665 12937 7699 12971
rect 9505 12937 9539 12971
rect 10425 12937 10459 12971
rect 11253 12937 11287 12971
rect 13185 12937 13219 12971
rect 16405 12937 16439 12971
rect 18061 12937 18095 12971
rect 18889 12937 18923 12971
rect 19717 12937 19751 12971
rect 20545 12937 20579 12971
rect 4629 12869 4663 12903
rect 14657 12869 14691 12903
rect 2513 12801 2547 12835
rect 2973 12801 3007 12835
rect 3249 12801 3283 12835
rect 5733 12801 5767 12835
rect 5917 12801 5951 12835
rect 7481 12801 7515 12835
rect 8033 12801 8067 12835
rect 10057 12801 10091 12835
rect 10977 12801 11011 12835
rect 11805 12801 11839 12835
rect 13737 12801 13771 12835
rect 15301 12801 15335 12835
rect 16037 12801 16071 12835
rect 16957 12801 16991 12835
rect 18613 12801 18647 12835
rect 19441 12801 19475 12835
rect 20269 12801 20303 12835
rect 21097 12801 21131 12835
rect 1593 12733 1627 12767
rect 7205 12733 7239 12767
rect 7849 12733 7883 12767
rect 8289 12733 8323 12767
rect 9965 12733 9999 12767
rect 13645 12733 13679 12767
rect 19349 12733 19383 12767
rect 20085 12733 20119 12767
rect 21005 12733 21039 12767
rect 2421 12665 2455 12699
rect 3516 12665 3550 12699
rect 5641 12665 5675 12699
rect 7297 12665 7331 12699
rect 10793 12665 10827 12699
rect 10885 12665 10919 12699
rect 11621 12665 11655 12699
rect 12081 12665 12115 12699
rect 13553 12665 13587 12699
rect 14013 12665 14047 12699
rect 15025 12665 15059 12699
rect 15853 12665 15887 12699
rect 16865 12665 16899 12699
rect 20913 12665 20947 12699
rect 2329 12597 2363 12631
rect 9413 12597 9447 12631
rect 9873 12597 9907 12631
rect 11713 12597 11747 12631
rect 15117 12597 15151 12631
rect 15485 12597 15519 12631
rect 15945 12597 15979 12631
rect 16773 12597 16807 12631
rect 18429 12597 18463 12631
rect 18521 12597 18555 12631
rect 19257 12597 19291 12631
rect 20177 12597 20211 12631
rect 3249 12393 3283 12427
rect 8217 12393 8251 12427
rect 8585 12393 8619 12427
rect 9045 12393 9079 12427
rect 11529 12393 11563 12427
rect 13737 12393 13771 12427
rect 14381 12393 14415 12427
rect 16773 12393 16807 12427
rect 17233 12393 17267 12427
rect 18981 12393 19015 12427
rect 19073 12393 19107 12427
rect 3617 12325 3651 12359
rect 4721 12325 4755 12359
rect 11866 12325 11900 12359
rect 17141 12325 17175 12359
rect 17868 12325 17902 12359
rect 19616 12325 19650 12359
rect 1501 12257 1535 12291
rect 2136 12257 2170 12291
rect 3341 12257 3375 12291
rect 6368 12257 6402 12291
rect 8125 12257 8159 12291
rect 8953 12257 8987 12291
rect 10416 12257 10450 12291
rect 13921 12257 13955 12291
rect 14749 12257 14783 12291
rect 15568 12257 15602 12291
rect 17601 12257 17635 12291
rect 19349 12257 19383 12291
rect 21005 12257 21039 12291
rect 1869 12189 1903 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 6101 12189 6135 12223
rect 8309 12189 8343 12223
rect 9229 12189 9263 12223
rect 10149 12189 10183 12223
rect 11621 12189 11655 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 15301 12189 15335 12223
rect 17325 12189 17359 12223
rect 7481 12121 7515 12155
rect 16681 12121 16715 12155
rect 1685 12053 1719 12087
rect 4353 12053 4387 12087
rect 7757 12053 7791 12087
rect 13001 12053 13035 12087
rect 20729 12053 20763 12087
rect 21189 12053 21223 12087
rect 1593 11849 1627 11883
rect 5917 11849 5951 11883
rect 8309 11849 8343 11883
rect 9137 11849 9171 11883
rect 15669 11849 15703 11883
rect 17141 11849 17175 11883
rect 18061 11849 18095 11883
rect 8217 11781 8251 11815
rect 10241 11781 10275 11815
rect 1777 11713 1811 11747
rect 4261 11713 4295 11747
rect 4997 11713 5031 11747
rect 5089 11713 5123 11747
rect 6469 11713 6503 11747
rect 6837 11713 6871 11747
rect 8769 11713 8803 11747
rect 8861 11713 8895 11747
rect 9597 11713 9631 11747
rect 9689 11713 9723 11747
rect 10793 11713 10827 11747
rect 11529 11713 11563 11747
rect 11621 11713 11655 11747
rect 18613 11713 18647 11747
rect 19441 11713 19475 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 20821 11713 20855 11747
rect 1409 11645 1443 11679
rect 6285 11645 6319 11679
rect 7104 11645 7138 11679
rect 8677 11645 8711 11679
rect 10609 11645 10643 11679
rect 11437 11645 11471 11679
rect 12449 11645 12483 11679
rect 12716 11645 12750 11679
rect 14289 11645 14323 11679
rect 15761 11645 15795 11679
rect 16028 11645 16062 11679
rect 19349 11645 19383 11679
rect 20545 11645 20579 11679
rect 2044 11577 2078 11611
rect 14556 11577 14590 11611
rect 18429 11577 18463 11611
rect 20085 11577 20119 11611
rect 3157 11509 3191 11543
rect 3709 11509 3743 11543
rect 4077 11509 4111 11543
rect 4169 11509 4203 11543
rect 4537 11509 4571 11543
rect 4905 11509 4939 11543
rect 5641 11509 5675 11543
rect 6377 11509 6411 11543
rect 9505 11509 9539 11543
rect 10701 11509 10735 11543
rect 11069 11509 11103 11543
rect 13829 11509 13863 11543
rect 18521 11509 18555 11543
rect 18889 11509 18923 11543
rect 19257 11509 19291 11543
rect 19717 11509 19751 11543
rect 1685 11305 1719 11339
rect 2145 11305 2179 11339
rect 3893 11305 3927 11339
rect 4813 11305 4847 11339
rect 6469 11305 6503 11339
rect 14381 11305 14415 11339
rect 15301 11305 15335 11339
rect 16129 11305 16163 11339
rect 16589 11305 16623 11339
rect 17601 11305 17635 11339
rect 18429 11305 18463 11339
rect 21097 11305 21131 11339
rect 2053 11237 2087 11271
rect 6561 11237 6595 11271
rect 12900 11237 12934 11271
rect 14749 11237 14783 11271
rect 16497 11237 16531 11271
rect 18797 11237 18831 11271
rect 19616 11237 19650 11271
rect 2513 11169 2547 11203
rect 2780 11169 2814 11203
rect 5181 11169 5215 11203
rect 7481 11169 7515 11203
rect 7840 11169 7874 11203
rect 10517 11169 10551 11203
rect 12265 11169 12299 11203
rect 15669 11169 15703 11203
rect 17969 11169 18003 11203
rect 18061 11169 18095 11203
rect 19349 11169 19383 11203
rect 20913 11169 20947 11203
rect 2329 11101 2363 11135
rect 5273 11101 5307 11135
rect 5365 11101 5399 11135
rect 6653 11101 6687 11135
rect 7573 11101 7607 11135
rect 12633 11101 12667 11135
rect 14841 11101 14875 11135
rect 14933 11101 14967 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 16681 11101 16715 11135
rect 16957 11101 16991 11135
rect 17417 11101 17451 11135
rect 18153 11101 18187 11135
rect 18889 11101 18923 11135
rect 19073 11101 19107 11135
rect 6101 11033 6135 11067
rect 7297 11033 7331 11067
rect 8953 10965 8987 10999
rect 14013 10965 14047 10999
rect 20729 10965 20763 10999
rect 1593 10761 1627 10795
rect 3249 10761 3283 10795
rect 4905 10761 4939 10795
rect 9045 10761 9079 10795
rect 11345 10761 11379 10795
rect 12449 10761 12483 10795
rect 14657 10761 14691 10795
rect 16129 10761 16163 10795
rect 16957 10761 16991 10795
rect 19901 10761 19935 10795
rect 11253 10693 11287 10727
rect 2145 10625 2179 10659
rect 3065 10625 3099 10659
rect 3893 10625 3927 10659
rect 4629 10625 4663 10659
rect 5457 10625 5491 10659
rect 6285 10625 6319 10659
rect 7573 10625 7607 10659
rect 8861 10625 8895 10659
rect 9689 10625 9723 10659
rect 9873 10625 9907 10659
rect 11897 10625 11931 10659
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 13829 10625 13863 10659
rect 15301 10625 15335 10659
rect 16773 10625 16807 10659
rect 17509 10625 17543 10659
rect 20545 10625 20579 10659
rect 21005 10625 21039 10659
rect 3709 10557 3743 10591
rect 4445 10557 4479 10591
rect 5273 10557 5307 10591
rect 8677 10557 8711 10591
rect 11713 10557 11747 10591
rect 12817 10557 12851 10591
rect 14565 10557 14599 10591
rect 16497 10557 16531 10591
rect 17325 10557 17359 10591
rect 18521 10557 18555 10591
rect 20361 10557 20395 10591
rect 20821 10557 20855 10591
rect 1961 10489 1995 10523
rect 2881 10489 2915 10523
rect 3617 10489 3651 10523
rect 5365 10489 5399 10523
rect 10140 10489 10174 10523
rect 11805 10489 11839 10523
rect 13645 10489 13679 10523
rect 14105 10489 14139 10523
rect 15117 10489 15151 10523
rect 18766 10489 18800 10523
rect 2053 10421 2087 10455
rect 2421 10421 2455 10455
rect 2789 10421 2823 10455
rect 4077 10421 4111 10455
rect 4537 10421 4571 10455
rect 5733 10421 5767 10455
rect 6101 10421 6135 10455
rect 6193 10421 6227 10455
rect 7021 10421 7055 10455
rect 7389 10421 7423 10455
rect 7481 10421 7515 10455
rect 8217 10421 8251 10455
rect 8585 10421 8619 10455
rect 9413 10421 9447 10455
rect 9505 10421 9539 10455
rect 13277 10421 13311 10455
rect 13737 10421 13771 10455
rect 14381 10421 14415 10455
rect 15025 10421 15059 10455
rect 16589 10421 16623 10455
rect 17417 10421 17451 10455
rect 19993 10421 20027 10455
rect 20453 10421 20487 10455
rect 1593 10217 1627 10251
rect 2053 10217 2087 10251
rect 2421 10217 2455 10251
rect 3249 10217 3283 10251
rect 6929 10217 6963 10251
rect 9137 10217 9171 10251
rect 10425 10217 10459 10251
rect 11253 10217 11287 10251
rect 13921 10217 13955 10251
rect 14013 10217 14047 10251
rect 16681 10217 16715 10251
rect 18889 10217 18923 10251
rect 19625 10217 19659 10251
rect 2881 10149 2915 10183
rect 4344 10149 4378 10183
rect 10793 10149 10827 10183
rect 11713 10149 11747 10183
rect 13461 10149 13495 10183
rect 17776 10149 17810 10183
rect 1961 10081 1995 10115
rect 2789 10081 2823 10115
rect 6285 10081 6319 10115
rect 7297 10081 7331 10115
rect 8024 10081 8058 10115
rect 10885 10081 10919 10115
rect 11621 10081 11655 10115
rect 13001 10081 13035 10115
rect 2145 10013 2179 10047
rect 3065 10013 3099 10047
rect 4077 10013 4111 10047
rect 6377 10013 6411 10047
rect 6561 10013 6595 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 11069 10013 11103 10047
rect 11805 10013 11839 10047
rect 13093 10013 13127 10047
rect 13277 10013 13311 10047
rect 14749 10081 14783 10115
rect 15568 10081 15602 10115
rect 19993 10081 20027 10115
rect 14197 10013 14231 10047
rect 14841 10013 14875 10047
rect 15025 10013 15059 10047
rect 15301 10013 15335 10047
rect 17509 10013 17543 10047
rect 20085 10013 20119 10047
rect 20177 10013 20211 10047
rect 5917 9945 5951 9979
rect 13461 9945 13495 9979
rect 14381 9945 14415 9979
rect 5457 9877 5491 9911
rect 12633 9877 12667 9911
rect 13553 9877 13587 9911
rect 2145 9673 2179 9707
rect 4353 9673 4387 9707
rect 8217 9673 8251 9707
rect 20269 9673 20303 9707
rect 8585 9605 8619 9639
rect 11529 9605 11563 9639
rect 13921 9605 13955 9639
rect 15577 9605 15611 9639
rect 18061 9605 18095 9639
rect 19441 9605 19475 9639
rect 2789 9537 2823 9571
rect 6285 9537 6319 9571
rect 9137 9537 9171 9571
rect 10057 9537 10091 9571
rect 11345 9537 11379 9571
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 14565 9537 14599 9571
rect 15301 9537 15335 9571
rect 16037 9537 16071 9571
rect 16221 9537 16255 9571
rect 17049 9537 17083 9571
rect 18705 9537 18739 9571
rect 19993 9537 20027 9571
rect 20821 9537 20855 9571
rect 1777 9469 1811 9503
rect 2513 9469 2547 9503
rect 2973 9469 3007 9503
rect 4813 9469 4847 9503
rect 5080 9469 5114 9503
rect 6837 9469 6871 9503
rect 8493 9469 8527 9503
rect 9045 9469 9079 9503
rect 11161 9469 11195 9503
rect 11897 9469 11931 9503
rect 12449 9469 12483 9503
rect 15117 9469 15151 9503
rect 15209 9469 15243 9503
rect 18429 9469 18463 9503
rect 20637 9469 20671 9503
rect 20729 9469 20763 9503
rect 3218 9401 3252 9435
rect 7082 9401 7116 9435
rect 8953 9401 8987 9435
rect 9873 9401 9907 9435
rect 11069 9401 11103 9435
rect 12716 9401 12750 9435
rect 14381 9401 14415 9435
rect 15945 9401 15979 9435
rect 16865 9401 16899 9435
rect 1961 9333 1995 9367
rect 2605 9333 2639 9367
rect 6193 9333 6227 9367
rect 8309 9333 8343 9367
rect 9505 9333 9539 9367
rect 9965 9333 9999 9367
rect 10701 9333 10735 9367
rect 13829 9333 13863 9367
rect 14289 9333 14323 9367
rect 14749 9333 14783 9367
rect 16405 9333 16439 9367
rect 16773 9333 16807 9367
rect 18521 9333 18555 9367
rect 19809 9333 19843 9367
rect 19901 9333 19935 9367
rect 2421 9129 2455 9163
rect 5365 9129 5399 9163
rect 5733 9129 5767 9163
rect 6285 9129 6319 9163
rect 6745 9129 6779 9163
rect 7297 9129 7331 9163
rect 7757 9129 7791 9163
rect 8125 9129 8159 9163
rect 11069 9129 11103 9163
rect 13645 9129 13679 9163
rect 15393 9129 15427 9163
rect 15761 9129 15795 9163
rect 18061 9129 18095 9163
rect 18521 9129 18555 9163
rect 19993 9129 20027 9163
rect 2789 9061 2823 9095
rect 5825 9061 5859 9095
rect 8493 9061 8527 9095
rect 8585 9061 8619 9095
rect 11980 9061 12014 9095
rect 14381 9061 14415 9095
rect 16926 9061 16960 9095
rect 19533 9061 19567 9095
rect 2881 8993 2915 9027
rect 6653 8993 6687 9027
rect 7665 8993 7699 9027
rect 9956 8993 9990 9027
rect 13553 8993 13587 9027
rect 14473 8993 14507 9027
rect 15853 8993 15887 9027
rect 16405 8993 16439 9027
rect 19625 8993 19659 9027
rect 20361 8993 20395 9027
rect 3065 8925 3099 8959
rect 6009 8925 6043 8959
rect 6837 8925 6871 8959
rect 7849 8925 7883 8959
rect 8769 8925 8803 8959
rect 9689 8925 9723 8959
rect 11713 8925 11747 8959
rect 13829 8925 13863 8959
rect 14565 8925 14599 8959
rect 16037 8925 16071 8959
rect 16681 8925 16715 8959
rect 18613 8925 18647 8959
rect 18705 8925 18739 8959
rect 19717 8925 19751 8959
rect 20453 8925 20487 8959
rect 20545 8925 20579 8959
rect 16221 8857 16255 8891
rect 13093 8789 13127 8823
rect 13185 8789 13219 8823
rect 14013 8789 14047 8823
rect 18153 8789 18187 8823
rect 19165 8789 19199 8823
rect 1685 8585 1719 8619
rect 7665 8585 7699 8619
rect 11529 8585 11563 8619
rect 12633 8585 12667 8619
rect 14565 8585 14599 8619
rect 16957 8585 16991 8619
rect 18061 8585 18095 8619
rect 18889 8585 18923 8619
rect 2421 8517 2455 8551
rect 5457 8517 5491 8551
rect 10057 8517 10091 8551
rect 13737 8517 13771 8551
rect 16129 8517 16163 8551
rect 20269 8517 20303 8551
rect 2053 8449 2087 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3893 8449 3927 8483
rect 6009 8449 6043 8483
rect 7389 8449 7423 8483
rect 8217 8449 8251 8483
rect 13277 8449 13311 8483
rect 15117 8449 15151 8483
rect 16681 8449 16715 8483
rect 17509 8449 17543 8483
rect 18613 8449 18647 8483
rect 19533 8449 19567 8483
rect 19901 8449 19935 8483
rect 20821 8449 20855 8483
rect 1501 8381 1535 8415
rect 1869 8381 1903 8415
rect 3709 8381 3743 8415
rect 7297 8381 7331 8415
rect 8677 8381 8711 8415
rect 10156 8381 10190 8415
rect 10405 8381 10439 8415
rect 13093 8381 13127 8415
rect 13921 8381 13955 8415
rect 16589 8381 16623 8415
rect 17325 8381 17359 8415
rect 18429 8381 18463 8415
rect 19349 8381 19383 8415
rect 20729 8381 20763 8415
rect 3617 8313 3651 8347
rect 5825 8313 5859 8347
rect 7205 8313 7239 8347
rect 8033 8313 8067 8347
rect 8125 8313 8159 8347
rect 8944 8313 8978 8347
rect 14933 8313 14967 8347
rect 16497 8313 16531 8347
rect 19257 8313 19291 8347
rect 2789 8245 2823 8279
rect 3249 8245 3283 8279
rect 5917 8245 5951 8279
rect 6837 8245 6871 8279
rect 11621 8245 11655 8279
rect 13001 8245 13035 8279
rect 15025 8245 15059 8279
rect 17417 8245 17451 8279
rect 18521 8245 18555 8279
rect 20637 8245 20671 8279
rect 2973 8041 3007 8075
rect 3525 8041 3559 8075
rect 5549 8041 5583 8075
rect 6285 8041 6319 8075
rect 6653 8041 6687 8075
rect 7113 8041 7147 8075
rect 7481 8041 7515 8075
rect 8401 8041 8435 8075
rect 8769 8041 8803 8075
rect 9689 8041 9723 8075
rect 10885 8041 10919 8075
rect 14381 8041 14415 8075
rect 16773 8041 16807 8075
rect 18521 8041 18555 8075
rect 20545 8041 20579 8075
rect 4436 7973 4470 8007
rect 8309 7973 8343 8007
rect 12808 7973 12842 8007
rect 17141 7973 17175 8007
rect 18429 7973 18463 8007
rect 19432 7973 19466 8007
rect 1860 7905 1894 7939
rect 4169 7905 4203 7939
rect 5917 7905 5951 7939
rect 7573 7905 7607 7939
rect 9137 7905 9171 7939
rect 10057 7905 10091 7939
rect 10977 7905 11011 7939
rect 14749 7905 14783 7939
rect 15568 7905 15602 7939
rect 17233 7905 17267 7939
rect 19165 7905 19199 7939
rect 1593 7837 1627 7871
rect 3617 7837 3651 7871
rect 3801 7837 3835 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 7757 7837 7791 7871
rect 8585 7837 8619 7871
rect 9229 7837 9263 7871
rect 9413 7837 9447 7871
rect 10149 7837 10183 7871
rect 10333 7837 10367 7871
rect 11069 7837 11103 7871
rect 12541 7837 12575 7871
rect 14841 7837 14875 7871
rect 15025 7837 15059 7871
rect 15301 7837 15335 7871
rect 17325 7837 17359 7871
rect 18613 7837 18647 7871
rect 5733 7769 5767 7803
rect 18061 7769 18095 7803
rect 3157 7701 3191 7735
rect 7941 7701 7975 7735
rect 10517 7701 10551 7735
rect 13921 7701 13955 7735
rect 16681 7701 16715 7735
rect 2789 7497 2823 7531
rect 3709 7497 3743 7531
rect 12449 7497 12483 7531
rect 14749 7497 14783 7531
rect 19901 7497 19935 7531
rect 5917 7429 5951 7463
rect 7113 7429 7147 7463
rect 7941 7429 7975 7463
rect 8401 7429 8435 7463
rect 17049 7429 17083 7463
rect 19809 7429 19843 7463
rect 1593 7361 1627 7395
rect 2605 7361 2639 7395
rect 3249 7361 3283 7395
rect 3433 7361 3467 7395
rect 4261 7361 4295 7395
rect 4537 7361 4571 7395
rect 7665 7361 7699 7395
rect 9045 7361 9079 7395
rect 9873 7361 9907 7395
rect 10609 7361 10643 7395
rect 13645 7361 13679 7395
rect 14473 7361 14507 7395
rect 15301 7361 15335 7395
rect 17693 7361 17727 7395
rect 20453 7361 20487 7395
rect 1409 7293 1443 7327
rect 3157 7293 3191 7327
rect 7481 7293 7515 7327
rect 8125 7293 8159 7327
rect 10517 7293 10551 7327
rect 10885 7293 10919 7327
rect 12633 7293 12667 7327
rect 13553 7293 13587 7327
rect 14381 7293 14415 7327
rect 15577 7293 15611 7327
rect 15844 7293 15878 7327
rect 17509 7293 17543 7327
rect 18429 7293 18463 7327
rect 18696 7293 18730 7327
rect 4169 7225 4203 7259
rect 4782 7225 4816 7259
rect 10425 7225 10459 7259
rect 11152 7225 11186 7259
rect 12725 7225 12759 7259
rect 14289 7225 14323 7259
rect 15117 7225 15151 7259
rect 15209 7225 15243 7259
rect 17417 7225 17451 7259
rect 18061 7225 18095 7259
rect 20361 7225 20395 7259
rect 1961 7157 1995 7191
rect 2329 7157 2363 7191
rect 2421 7157 2455 7191
rect 4077 7157 4111 7191
rect 7021 7157 7055 7191
rect 7573 7157 7607 7191
rect 8769 7157 8803 7191
rect 8861 7157 8895 7191
rect 9229 7157 9263 7191
rect 9597 7157 9631 7191
rect 9689 7157 9723 7191
rect 10057 7157 10091 7191
rect 12265 7157 12299 7191
rect 13093 7157 13127 7191
rect 13461 7157 13495 7191
rect 13921 7157 13955 7191
rect 16957 7157 16991 7191
rect 20269 7157 20303 7191
rect 1685 6953 1719 6987
rect 3893 6953 3927 6987
rect 7113 6953 7147 6987
rect 8769 6953 8803 6987
rect 9137 6953 9171 6987
rect 9689 6953 9723 6987
rect 10057 6953 10091 6987
rect 12909 6953 12943 6987
rect 13737 6953 13771 6987
rect 15669 6953 15703 6987
rect 19717 6953 19751 6987
rect 19809 6953 19843 6987
rect 2053 6885 2087 6919
rect 10149 6885 10183 6919
rect 11590 6885 11624 6919
rect 14105 6885 14139 6919
rect 17417 6885 17451 6919
rect 2513 6817 2547 6851
rect 2780 6817 2814 6851
rect 4077 6817 4111 6851
rect 4813 6817 4847 6851
rect 5080 6817 5114 6851
rect 7021 6817 7055 6851
rect 7849 6817 7883 6851
rect 9229 6817 9263 6851
rect 13277 6817 13311 6851
rect 16129 6817 16163 6851
rect 18337 6817 18371 6851
rect 18604 6817 18638 6851
rect 20177 6817 20211 6851
rect 2145 6749 2179 6783
rect 2329 6749 2363 6783
rect 7205 6749 7239 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 9413 6749 9447 6783
rect 10241 6749 10275 6783
rect 11345 6749 11379 6783
rect 13369 6749 13403 6783
rect 13461 6749 13495 6783
rect 14197 6749 14231 6783
rect 14381 6749 14415 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 17509 6749 17543 6783
rect 17693 6749 17727 6783
rect 20269 6749 20303 6783
rect 20361 6749 20395 6783
rect 6653 6681 6687 6715
rect 7481 6681 7515 6715
rect 15301 6681 15335 6715
rect 6193 6613 6227 6647
rect 6561 6613 6595 6647
rect 10517 6613 10551 6647
rect 12725 6613 12759 6647
rect 17049 6613 17083 6647
rect 2973 6409 3007 6443
rect 12541 6409 12575 6443
rect 19441 6409 19475 6443
rect 2881 6341 2915 6375
rect 10517 6341 10551 6375
rect 3525 6273 3559 6307
rect 4353 6273 4387 6307
rect 5181 6273 5215 6307
rect 6101 6273 6135 6307
rect 6837 6273 6871 6307
rect 11161 6273 11195 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 13093 6273 13127 6307
rect 15853 6273 15887 6307
rect 19993 6273 20027 6307
rect 20821 6273 20855 6307
rect 1501 6205 1535 6239
rect 1768 6205 1802 6239
rect 3433 6205 3467 6239
rect 4997 6205 5031 6239
rect 5089 6205 5123 6239
rect 7104 6205 7138 6239
rect 8677 6205 8711 6239
rect 11897 6205 11931 6239
rect 13001 6205 13035 6239
rect 13921 6205 13955 6239
rect 14013 6205 14047 6239
rect 16120 6205 16154 6239
rect 18061 6205 18095 6239
rect 20729 6205 20763 6239
rect 3341 6137 3375 6171
rect 8922 6137 8956 6171
rect 10977 6137 11011 6171
rect 12909 6137 12943 6171
rect 14280 6137 14314 6171
rect 18328 6137 18362 6171
rect 3801 6069 3835 6103
rect 4169 6069 4203 6103
rect 4261 6069 4295 6103
rect 4629 6069 4663 6103
rect 5457 6069 5491 6103
rect 5825 6069 5859 6103
rect 5917 6069 5951 6103
rect 8217 6069 8251 6103
rect 10057 6069 10091 6103
rect 10885 6069 10919 6103
rect 11529 6069 11563 6103
rect 13921 6069 13955 6103
rect 15393 6069 15427 6103
rect 17233 6069 17267 6103
rect 20269 6069 20303 6103
rect 20637 6069 20671 6103
rect 2973 5865 3007 5899
rect 6561 5865 6595 5899
rect 8125 5865 8159 5899
rect 10149 5865 10183 5899
rect 10885 5865 10919 5899
rect 11897 5865 11931 5899
rect 12909 5865 12943 5899
rect 14749 5865 14783 5899
rect 15301 5865 15335 5899
rect 15761 5865 15795 5899
rect 18245 5865 18279 5899
rect 18613 5865 18647 5899
rect 19533 5865 19567 5899
rect 19993 5865 20027 5899
rect 20361 5865 20395 5899
rect 3433 5797 3467 5831
rect 4353 5797 4387 5831
rect 4905 5797 4939 5831
rect 5641 5797 5675 5831
rect 6469 5797 6503 5831
rect 7665 5797 7699 5831
rect 8493 5797 8527 5831
rect 19073 5797 19107 5831
rect 19625 5797 19659 5831
rect 1593 5729 1627 5763
rect 1860 5729 1894 5763
rect 3525 5729 3559 5763
rect 4813 5729 4847 5763
rect 7205 5729 7239 5763
rect 7757 5729 7791 5763
rect 8585 5729 8619 5763
rect 10057 5729 10091 5763
rect 13277 5729 13311 5763
rect 13369 5729 13403 5763
rect 14841 5729 14875 5763
rect 15669 5729 15703 5763
rect 17029 5729 17063 5763
rect 18705 5729 18739 5763
rect 3709 5661 3743 5695
rect 5089 5661 5123 5695
rect 5733 5661 5767 5695
rect 5917 5661 5951 5695
rect 6745 5661 6779 5695
rect 7941 5661 7975 5695
rect 8677 5661 8711 5695
rect 10241 5661 10275 5695
rect 10977 5661 11011 5695
rect 11069 5661 11103 5695
rect 11989 5661 12023 5695
rect 12081 5661 12115 5695
rect 13553 5661 13587 5695
rect 15025 5661 15059 5695
rect 15945 5661 15979 5695
rect 16773 5661 16807 5695
rect 18797 5661 18831 5695
rect 18153 5593 18187 5627
rect 19717 5661 19751 5695
rect 20453 5661 20487 5695
rect 20545 5661 20579 5695
rect 3065 5525 3099 5559
rect 4445 5525 4479 5559
rect 5273 5525 5307 5559
rect 6101 5525 6135 5559
rect 7297 5525 7331 5559
rect 9689 5525 9723 5559
rect 10517 5525 10551 5559
rect 11529 5525 11563 5559
rect 14381 5525 14415 5559
rect 19073 5525 19107 5559
rect 19165 5525 19199 5559
rect 2145 5321 2179 5355
rect 4629 5321 4663 5355
rect 8861 5321 8895 5355
rect 11805 5321 11839 5355
rect 14381 5321 14415 5355
rect 15209 5321 15243 5355
rect 18889 5321 18923 5355
rect 19717 5321 19751 5355
rect 18061 5253 18095 5287
rect 2697 5185 2731 5219
rect 5089 5185 5123 5219
rect 5181 5185 5215 5219
rect 6561 5185 6595 5219
rect 7481 5185 7515 5219
rect 9321 5185 9355 5219
rect 10149 5185 10183 5219
rect 14013 5185 14047 5219
rect 14197 5185 14231 5219
rect 15025 5185 15059 5219
rect 15853 5185 15887 5219
rect 17141 5185 17175 5219
rect 18613 5185 18647 5219
rect 19441 5185 19475 5219
rect 20177 5185 20211 5219
rect 20361 5185 20395 5219
rect 20821 5185 20855 5219
rect 2513 5117 2547 5151
rect 2605 5117 2639 5151
rect 3157 5117 3191 5151
rect 3424 5117 3458 5151
rect 4997 5117 5031 5151
rect 9965 5117 9999 5151
rect 10425 5117 10459 5151
rect 14749 5117 14783 5151
rect 15669 5117 15703 5151
rect 16865 5117 16899 5151
rect 20085 5117 20119 5151
rect 20545 5117 20579 5151
rect 6285 5049 6319 5083
rect 6837 5049 6871 5083
rect 7748 5049 7782 5083
rect 10692 5049 10726 5083
rect 19349 5049 19383 5083
rect 1869 4981 1903 5015
rect 4537 4981 4571 5015
rect 5917 4981 5951 5015
rect 6377 4981 6411 5015
rect 9597 4981 9631 5015
rect 10057 4981 10091 5015
rect 13369 4981 13403 5015
rect 13553 4981 13587 5015
rect 13921 4981 13955 5015
rect 14841 4981 14875 5015
rect 15577 4981 15611 5015
rect 16497 4981 16531 5015
rect 16957 4981 16991 5015
rect 18429 4981 18463 5015
rect 18521 4981 18555 5015
rect 19257 4981 19291 5015
rect 1869 4777 1903 4811
rect 2237 4777 2271 4811
rect 4905 4777 4939 4811
rect 5365 4777 5399 4811
rect 6193 4777 6227 4811
rect 7021 4777 7055 4811
rect 7113 4777 7147 4811
rect 7481 4777 7515 4811
rect 9229 4777 9263 4811
rect 10333 4777 10367 4811
rect 11621 4777 11655 4811
rect 12633 4777 12667 4811
rect 12725 4777 12759 4811
rect 15301 4777 15335 4811
rect 18521 4777 18555 4811
rect 20729 4777 20763 4811
rect 7849 4709 7883 4743
rect 9137 4709 9171 4743
rect 10241 4709 10275 4743
rect 15761 4709 15795 4743
rect 17316 4709 17350 4743
rect 3433 4641 3467 4675
rect 6285 4641 6319 4675
rect 10701 4641 10735 4675
rect 11529 4641 11563 4675
rect 13093 4641 13127 4675
rect 13360 4641 13394 4675
rect 15669 4641 15703 4675
rect 18889 4641 18923 4675
rect 19349 4641 19383 4675
rect 19616 4641 19650 4675
rect 2329 4573 2363 4607
rect 2513 4573 2547 4607
rect 3525 4573 3559 4607
rect 3709 4573 3743 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 6377 4573 6411 4607
rect 7205 4573 7239 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 9413 4573 9447 4607
rect 10241 4573 10275 4607
rect 10793 4573 10827 4607
rect 10977 4573 11011 4607
rect 11713 4573 11747 4607
rect 12909 4573 12943 4607
rect 15945 4573 15979 4607
rect 17049 4573 17083 4607
rect 18981 4573 19015 4607
rect 19073 4573 19107 4607
rect 18429 4505 18463 4539
rect 3065 4437 3099 4471
rect 4997 4437 5031 4471
rect 5825 4437 5859 4471
rect 6653 4437 6687 4471
rect 8769 4437 8803 4471
rect 11161 4437 11195 4471
rect 12265 4437 12299 4471
rect 14473 4437 14507 4471
rect 4261 4233 4295 4267
rect 19717 4233 19751 4267
rect 10517 4165 10551 4199
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 4905 4097 4939 4131
rect 5733 4097 5767 4131
rect 7481 4097 7515 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 8769 4097 8803 4131
rect 11069 4097 11103 4131
rect 11897 4097 11931 4131
rect 13185 4097 13219 4131
rect 13829 4097 13863 4131
rect 14013 4097 14047 4131
rect 14841 4097 14875 4131
rect 15025 4097 15059 4131
rect 17049 4097 17083 4131
rect 2421 4029 2455 4063
rect 3148 4029 3182 4063
rect 4813 4029 4847 4063
rect 7297 4029 7331 4063
rect 9036 4029 9070 4063
rect 11713 4029 11747 4063
rect 13737 4029 13771 4063
rect 16773 4029 16807 4063
rect 18337 4029 18371 4063
rect 18604 4029 18638 4063
rect 4721 3961 4755 3995
rect 5641 3961 5675 3995
rect 8125 3961 8159 3995
rect 10977 3961 11011 3995
rect 12909 3961 12943 3995
rect 14749 3961 14783 3995
rect 15209 3961 15243 3995
rect 2053 3893 2087 3927
rect 2513 3893 2547 3927
rect 4353 3893 4387 3927
rect 5181 3893 5215 3927
rect 5549 3893 5583 3927
rect 6929 3893 6963 3927
rect 7389 3893 7423 3927
rect 7757 3893 7791 3927
rect 10149 3893 10183 3927
rect 10885 3893 10919 3927
rect 11345 3893 11379 3927
rect 11805 3893 11839 3927
rect 12541 3893 12575 3927
rect 13001 3893 13035 3927
rect 13369 3893 13403 3927
rect 14381 3893 14415 3927
rect 16405 3893 16439 3927
rect 16865 3893 16899 3927
rect 18061 3893 18095 3927
rect 3525 3689 3559 3723
rect 4629 3689 4663 3723
rect 6377 3689 6411 3723
rect 7941 3689 7975 3723
rect 11069 3689 11103 3723
rect 11529 3689 11563 3723
rect 11897 3689 11931 3723
rect 13001 3689 13035 3723
rect 14841 3689 14875 3723
rect 15485 3689 15519 3723
rect 17601 3689 17635 3723
rect 18429 3689 18463 3723
rect 19717 3689 19751 3723
rect 4537 3621 4571 3655
rect 6736 3621 6770 3655
rect 9229 3621 9263 3655
rect 11989 3621 12023 3655
rect 13093 3621 13127 3655
rect 13728 3621 13762 3655
rect 15853 3621 15887 3655
rect 15945 3621 15979 3655
rect 17141 3621 17175 3655
rect 17233 3621 17267 3655
rect 18797 3621 18831 3655
rect 19625 3621 19659 3655
rect 2053 3553 2087 3587
rect 2320 3553 2354 3587
rect 5253 3553 5287 3587
rect 8309 3553 8343 3587
rect 9137 3553 9171 3587
rect 9689 3553 9723 3587
rect 9956 3553 9990 3587
rect 11161 3553 11195 3587
rect 16313 3553 16347 3587
rect 17969 3553 18003 3587
rect 18061 3553 18095 3587
rect 4813 3485 4847 3519
rect 4997 3485 5031 3519
rect 6469 3485 6503 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 9321 3485 9355 3519
rect 12173 3485 12207 3519
rect 13277 3485 13311 3519
rect 13461 3485 13495 3519
rect 16129 3485 16163 3519
rect 17325 3485 17359 3519
rect 18153 3485 18187 3519
rect 18889 3485 18923 3519
rect 18981 3485 19015 3519
rect 19809 3485 19843 3519
rect 19257 3417 19291 3451
rect 3433 3349 3467 3383
rect 4169 3349 4203 3383
rect 7849 3349 7883 3383
rect 8769 3349 8803 3383
rect 11345 3349 11379 3383
rect 12633 3349 12667 3383
rect 16497 3349 16531 3383
rect 16773 3349 16807 3383
rect 2237 3145 2271 3179
rect 6285 3145 6319 3179
rect 10333 3145 10367 3179
rect 13829 3145 13863 3179
rect 15025 3145 15059 3179
rect 17325 3145 17359 3179
rect 18061 3145 18095 3179
rect 4445 3077 4479 3111
rect 14105 3077 14139 3111
rect 17601 3077 17635 3111
rect 2697 3009 2731 3043
rect 2881 3009 2915 3043
rect 10977 3009 11011 3043
rect 12449 3009 12483 3043
rect 15485 3009 15519 3043
rect 15669 3009 15703 3043
rect 15945 3009 15979 3043
rect 18613 3009 18647 3043
rect 2605 2941 2639 2975
rect 3065 2941 3099 2975
rect 4905 2941 4939 2975
rect 7481 2941 7515 2975
rect 7748 2941 7782 2975
rect 8953 2941 8987 2975
rect 9220 2941 9254 2975
rect 11253 2941 11287 2975
rect 11805 2941 11839 2975
rect 13921 2941 13955 2975
rect 14381 2941 14415 2975
rect 17417 2941 17451 2975
rect 18429 2941 18463 2975
rect 18889 2941 18923 2975
rect 3310 2873 3344 2907
rect 5172 2873 5206 2907
rect 10793 2873 10827 2907
rect 11529 2873 11563 2907
rect 12081 2873 12115 2907
rect 12716 2873 12750 2907
rect 14657 2873 14691 2907
rect 16212 2873 16246 2907
rect 8861 2805 8895 2839
rect 10425 2805 10459 2839
rect 10885 2805 10919 2839
rect 15393 2805 15427 2839
rect 18521 2805 18555 2839
rect 19073 2805 19107 2839
rect 3157 2601 3191 2635
rect 5365 2601 5399 2635
rect 7481 2601 7515 2635
rect 8309 2601 8343 2635
rect 8769 2601 8803 2635
rect 9781 2601 9815 2635
rect 10149 2601 10183 2635
rect 10241 2601 10275 2635
rect 14841 2601 14875 2635
rect 16405 2601 16439 2635
rect 17141 2601 17175 2635
rect 18337 2601 18371 2635
rect 18797 2601 18831 2635
rect 19717 2601 19751 2635
rect 3617 2533 3651 2567
rect 7941 2533 7975 2567
rect 8677 2533 8711 2567
rect 10885 2533 10919 2567
rect 11437 2533 11471 2567
rect 3525 2465 3559 2499
rect 4905 2465 4939 2499
rect 5733 2465 5767 2499
rect 5825 2465 5859 2499
rect 7849 2465 7883 2499
rect 10609 2465 10643 2499
rect 11161 2465 11195 2499
rect 11897 2465 11931 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13578 2465 13612 2499
rect 13921 2465 13955 2499
rect 14289 2465 14323 2499
rect 14657 2465 14691 2499
rect 15025 2465 15059 2499
rect 15669 2465 15703 2499
rect 16221 2465 16255 2499
rect 16589 2465 16623 2499
rect 16957 2465 16991 2499
rect 17325 2465 17359 2499
rect 17693 2465 17727 2499
rect 18705 2465 18739 2499
rect 19165 2465 19199 2499
rect 19533 2465 19567 2499
rect 19901 2465 19935 2499
rect 3709 2397 3743 2431
rect 4997 2397 5031 2431
rect 5181 2397 5215 2431
rect 5917 2397 5951 2431
rect 8033 2397 8067 2431
rect 8861 2397 8895 2431
rect 10333 2397 10367 2431
rect 12909 2397 12943 2431
rect 15945 2397 15979 2431
rect 18981 2397 19015 2431
rect 4537 2329 4571 2363
rect 14473 2329 14507 2363
rect 17877 2329 17911 2363
rect 20085 2329 20119 2363
rect 12081 2261 12115 2295
rect 13369 2261 13403 2295
rect 13737 2261 13771 2295
rect 14105 2261 14139 2295
rect 15209 2261 15243 2295
rect 16773 2261 16807 2295
rect 17509 2261 17543 2295
rect 19349 2261 19383 2295
<< metal1 >>
rect 7006 20544 7012 20596
rect 7064 20584 7070 20596
rect 7558 20584 7564 20596
rect 7064 20556 7564 20584
rect 7064 20544 7070 20556
rect 7558 20544 7564 20556
rect 7616 20544 7622 20596
rect 4338 20340 4344 20392
rect 4396 20380 4402 20392
rect 9030 20380 9036 20392
rect 4396 20352 9036 20380
rect 4396 20340 4402 20352
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 7098 20272 7104 20324
rect 7156 20312 7162 20324
rect 8110 20312 8116 20324
rect 7156 20284 8116 20312
rect 7156 20272 7162 20284
rect 8110 20272 8116 20284
rect 8168 20272 8174 20324
rect 4062 20204 4068 20256
rect 4120 20244 4126 20256
rect 15194 20244 15200 20256
rect 4120 20216 15200 20244
rect 4120 20204 4126 20216
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 20622 20244 20628 20256
rect 19392 20216 20628 20244
rect 19392 20204 19398 20216
rect 20622 20204 20628 20216
rect 20680 20204 20686 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 4798 20000 4804 20052
rect 4856 20040 4862 20052
rect 9766 20040 9772 20052
rect 4856 20012 9772 20040
rect 4856 20000 4862 20012
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 13449 20043 13507 20049
rect 13449 20009 13461 20043
rect 13495 20040 13507 20043
rect 13814 20040 13820 20052
rect 13495 20012 13820 20040
rect 13495 20009 13507 20012
rect 13449 20003 13507 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 15657 20043 15715 20049
rect 15657 20009 15669 20043
rect 15703 20040 15715 20043
rect 15746 20040 15752 20052
rect 15703 20012 15752 20040
rect 15703 20009 15715 20012
rect 15657 20003 15715 20009
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 16025 20043 16083 20049
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 16114 20040 16120 20052
rect 16071 20012 16120 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 22186 20040 22192 20052
rect 19628 20012 22192 20040
rect 5166 19972 5172 19984
rect 3620 19944 5172 19972
rect 3620 19913 3648 19944
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 7193 19975 7251 19981
rect 7193 19941 7205 19975
rect 7239 19972 7251 19975
rect 10134 19972 10140 19984
rect 7239 19944 10140 19972
rect 7239 19941 7251 19944
rect 7193 19935 7251 19941
rect 10134 19932 10140 19944
rect 10192 19932 10198 19984
rect 19628 19981 19656 20012
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 19613 19975 19671 19981
rect 18800 19944 19564 19972
rect 3605 19907 3663 19913
rect 3605 19873 3617 19907
rect 3651 19873 3663 19907
rect 3605 19867 3663 19873
rect 4516 19907 4574 19913
rect 4516 19873 4528 19907
rect 4562 19904 4574 19907
rect 5534 19904 5540 19916
rect 4562 19876 5540 19904
rect 4562 19873 4574 19876
rect 4516 19867 4574 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 6917 19907 6975 19913
rect 6917 19904 6929 19907
rect 6880 19876 6929 19904
rect 6880 19864 6886 19876
rect 6917 19873 6929 19876
rect 6963 19873 6975 19907
rect 6917 19867 6975 19873
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 7929 19907 7987 19913
rect 7929 19904 7941 19907
rect 7340 19876 7941 19904
rect 7340 19864 7346 19876
rect 7929 19873 7941 19876
rect 7975 19873 7987 19907
rect 7929 19867 7987 19873
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19904 8079 19907
rect 8202 19904 8208 19916
rect 8067 19876 8208 19904
rect 8067 19873 8079 19876
rect 8021 19867 8079 19873
rect 8202 19864 8208 19876
rect 8260 19864 8266 19916
rect 13262 19904 13268 19916
rect 13223 19876 13268 19904
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 15838 19904 15844 19916
rect 15799 19876 15844 19904
rect 15473 19867 15531 19873
rect 4246 19836 4252 19848
rect 4207 19808 4252 19836
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 7800 19808 8125 19836
rect 7800 19796 7806 19808
rect 8113 19805 8125 19808
rect 8159 19805 8171 19839
rect 15488 19836 15516 19867
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18800 19904 18828 19944
rect 19536 19916 19564 19944
rect 19613 19941 19625 19975
rect 19659 19941 19671 19975
rect 19613 19935 19671 19941
rect 20717 19975 20775 19981
rect 20717 19941 20729 19975
rect 20763 19972 20775 19975
rect 21450 19972 21456 19984
rect 20763 19944 21456 19972
rect 20763 19941 20775 19944
rect 20717 19935 20775 19941
rect 21450 19932 21456 19944
rect 21508 19932 21514 19984
rect 19334 19904 19340 19916
rect 18371 19876 18828 19904
rect 19295 19876 19340 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 19518 19864 19524 19916
rect 19576 19904 19582 19916
rect 19794 19904 19800 19916
rect 19576 19876 19800 19904
rect 19576 19864 19582 19876
rect 19794 19864 19800 19876
rect 19852 19904 19858 19916
rect 19889 19907 19947 19913
rect 19889 19904 19901 19907
rect 19852 19876 19901 19904
rect 19852 19864 19858 19876
rect 19889 19873 19901 19876
rect 19935 19873 19947 19907
rect 20438 19904 20444 19916
rect 19889 19867 19947 19873
rect 19996 19876 20444 19904
rect 16298 19836 16304 19848
rect 15488 19808 16304 19836
rect 8113 19799 8171 19805
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 11606 19768 11612 19780
rect 5552 19740 11612 19768
rect 3789 19703 3847 19709
rect 3789 19669 3801 19703
rect 3835 19700 3847 19703
rect 5552 19700 5580 19740
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 3835 19672 5580 19700
rect 3835 19669 3847 19672
rect 3789 19663 3847 19669
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 5684 19672 5729 19700
rect 5684 19660 5690 19672
rect 5810 19660 5816 19712
rect 5868 19700 5874 19712
rect 7561 19703 7619 19709
rect 7561 19700 7573 19703
rect 5868 19672 7573 19700
rect 5868 19660 5874 19672
rect 7561 19669 7573 19672
rect 7607 19669 7619 19703
rect 7561 19663 7619 19669
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 18524 19700 18552 19799
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19996 19836 20024 19876
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 19208 19808 20024 19836
rect 20165 19839 20223 19845
rect 19208 19796 19214 19808
rect 20165 19805 20177 19839
rect 20211 19836 20223 19839
rect 21818 19836 21824 19848
rect 20211 19808 21824 19836
rect 20211 19805 20223 19808
rect 20165 19799 20223 19805
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 9824 19672 18552 19700
rect 9824 19660 9830 19672
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 4246 19456 4252 19508
rect 4304 19496 4310 19508
rect 5534 19496 5540 19508
rect 4304 19468 4660 19496
rect 4304 19456 4310 19468
rect 4632 19440 4660 19468
rect 4724 19468 5540 19496
rect 2792 19400 4568 19428
rect 198 19252 204 19304
rect 256 19292 262 19304
rect 2792 19292 2820 19400
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19360 3847 19363
rect 4246 19360 4252 19372
rect 3835 19332 4252 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 4246 19320 4252 19332
rect 4304 19320 4310 19372
rect 4540 19301 4568 19400
rect 4614 19388 4620 19440
rect 4672 19388 4678 19440
rect 4724 19369 4752 19468
rect 5534 19456 5540 19468
rect 5592 19496 5598 19508
rect 6273 19499 6331 19505
rect 6273 19496 6285 19499
rect 5592 19468 6285 19496
rect 5592 19456 5598 19468
rect 6273 19465 6285 19468
rect 6319 19465 6331 19499
rect 6273 19459 6331 19465
rect 9674 19388 9680 19440
rect 9732 19388 9738 19440
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19329 4767 19363
rect 9214 19360 9220 19372
rect 4709 19323 4767 19329
rect 6840 19332 7052 19360
rect 9175 19332 9220 19360
rect 4433 19295 4491 19301
rect 4433 19292 4445 19295
rect 256 19264 2820 19292
rect 2884 19264 4445 19292
rect 256 19252 262 19264
rect 566 19184 572 19236
rect 624 19224 630 19236
rect 2884 19224 2912 19264
rect 4433 19261 4445 19264
rect 4479 19261 4491 19295
rect 4433 19255 4491 19261
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 4798 19292 4804 19304
rect 4571 19264 4804 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 3513 19227 3571 19233
rect 3513 19224 3525 19227
rect 624 19196 2912 19224
rect 2976 19196 3525 19224
rect 624 19184 630 19196
rect 2976 19168 3004 19196
rect 3513 19193 3525 19196
rect 3559 19193 3571 19227
rect 3513 19187 3571 19193
rect 3605 19227 3663 19233
rect 3605 19193 3617 19227
rect 3651 19224 3663 19227
rect 4154 19224 4160 19236
rect 3651 19196 4160 19224
rect 3651 19193 3663 19196
rect 3605 19187 3663 19193
rect 4154 19184 4160 19196
rect 4212 19184 4218 19236
rect 4448 19224 4476 19255
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 4893 19295 4951 19301
rect 4893 19261 4905 19295
rect 4939 19292 4951 19295
rect 4982 19292 4988 19304
rect 4939 19264 4988 19292
rect 4939 19261 4951 19264
rect 4893 19255 4951 19261
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 5160 19227 5218 19233
rect 4448 19196 5120 19224
rect 2958 19116 2964 19168
rect 3016 19116 3022 19168
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 3418 19156 3424 19168
rect 3191 19128 3424 19156
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 4062 19156 4068 19168
rect 4023 19128 4068 19156
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 4982 19156 4988 19168
rect 4672 19128 4988 19156
rect 4672 19116 4678 19128
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 5092 19156 5120 19196
rect 5160 19193 5172 19227
rect 5206 19224 5218 19227
rect 6086 19224 6092 19236
rect 5206 19196 6092 19224
rect 5206 19193 5218 19196
rect 5160 19187 5218 19193
rect 6086 19184 6092 19196
rect 6144 19184 6150 19236
rect 5258 19156 5264 19168
rect 5092 19128 5264 19156
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 5442 19116 5448 19168
rect 5500 19156 5506 19168
rect 6840 19156 6868 19332
rect 6917 19295 6975 19301
rect 6917 19261 6929 19295
rect 6963 19261 6975 19295
rect 7024 19292 7052 19332
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 7024 19264 9597 19292
rect 6917 19255 6975 19261
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 9692 19292 9720 19388
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19360 9919 19363
rect 12805 19363 12863 19369
rect 9907 19332 10548 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 9950 19292 9956 19304
rect 9692 19264 9956 19292
rect 9585 19255 9643 19261
rect 5500 19128 6868 19156
rect 6932 19156 6960 19255
rect 9950 19252 9956 19264
rect 10008 19252 10014 19304
rect 10134 19292 10140 19304
rect 10095 19264 10140 19292
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 10520 19301 10548 19332
rect 12805 19329 12817 19363
rect 12851 19360 12863 19363
rect 13262 19360 13268 19372
rect 12851 19332 13268 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 13262 19320 13268 19332
rect 13320 19320 13326 19372
rect 15194 19320 15200 19372
rect 15252 19360 15258 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15252 19332 16129 19360
rect 15252 19320 15258 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 10505 19295 10563 19301
rect 10505 19261 10517 19295
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 10870 19252 10876 19304
rect 10928 19292 10934 19304
rect 11425 19295 11483 19301
rect 11425 19292 11437 19295
rect 10928 19264 11437 19292
rect 10928 19252 10934 19264
rect 11425 19261 11437 19264
rect 11471 19261 11483 19295
rect 11425 19255 11483 19261
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 11882 19292 11888 19304
rect 11839 19264 11888 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 11882 19252 11888 19264
rect 11940 19252 11946 19304
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19292 12587 19295
rect 12986 19292 12992 19304
rect 12575 19264 12992 19292
rect 12575 19261 12587 19264
rect 12529 19255 12587 19261
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19261 13139 19295
rect 13446 19292 13452 19304
rect 13407 19264 13452 19292
rect 13081 19255 13139 19261
rect 7184 19227 7242 19233
rect 7184 19193 7196 19227
rect 7230 19224 7242 19227
rect 8662 19224 8668 19236
rect 7230 19196 8668 19224
rect 7230 19193 7242 19196
rect 7184 19187 7242 19193
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 9033 19227 9091 19233
rect 9033 19224 9045 19227
rect 8812 19196 9045 19224
rect 8812 19184 8818 19196
rect 9033 19193 9045 19196
rect 9079 19193 9091 19227
rect 10778 19224 10784 19236
rect 9033 19187 9091 19193
rect 10336 19196 10784 19224
rect 7650 19156 7656 19168
rect 6932 19128 7656 19156
rect 5500 19116 5506 19128
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 8297 19159 8355 19165
rect 8297 19156 8309 19159
rect 7800 19128 8309 19156
rect 7800 19116 7806 19128
rect 8297 19125 8309 19128
rect 8343 19125 8355 19159
rect 8570 19156 8576 19168
rect 8531 19128 8576 19156
rect 8297 19119 8355 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 8941 19159 8999 19165
rect 8941 19125 8953 19159
rect 8987 19156 8999 19159
rect 9122 19156 9128 19168
rect 8987 19128 9128 19156
rect 8987 19125 8999 19128
rect 8941 19119 8999 19125
rect 9122 19116 9128 19128
rect 9180 19156 9186 19168
rect 9490 19156 9496 19168
rect 9180 19128 9496 19156
rect 9180 19116 9186 19128
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 10336 19165 10364 19196
rect 10778 19184 10784 19196
rect 10836 19184 10842 19236
rect 12342 19224 12348 19236
rect 11624 19196 12348 19224
rect 10321 19159 10379 19165
rect 10321 19125 10333 19159
rect 10367 19125 10379 19159
rect 10321 19119 10379 19125
rect 10689 19159 10747 19165
rect 10689 19125 10701 19159
rect 10735 19156 10747 19159
rect 11146 19156 11152 19168
rect 10735 19128 11152 19156
rect 10735 19125 10747 19128
rect 10689 19119 10747 19125
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11624 19165 11652 19196
rect 12342 19184 12348 19196
rect 12400 19184 12406 19236
rect 12802 19184 12808 19236
rect 12860 19224 12866 19236
rect 13096 19224 13124 19255
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 13814 19292 13820 19304
rect 13775 19264 13820 19292
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 14185 19295 14243 19301
rect 14185 19292 14197 19295
rect 13964 19264 14197 19292
rect 13964 19252 13970 19264
rect 14185 19261 14197 19264
rect 14231 19261 14243 19295
rect 14185 19255 14243 19261
rect 14366 19252 14372 19304
rect 14424 19292 14430 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14424 19264 14565 19292
rect 14424 19252 14430 19264
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14553 19255 14611 19261
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 12860 19196 13124 19224
rect 12860 19184 12866 19196
rect 13170 19184 13176 19236
rect 13228 19224 13234 19236
rect 13228 19196 13400 19224
rect 13228 19184 13234 19196
rect 11609 19159 11667 19165
rect 11609 19125 11621 19159
rect 11655 19125 11667 19159
rect 11974 19156 11980 19168
rect 11935 19128 11980 19156
rect 11609 19119 11667 19125
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12710 19116 12716 19168
rect 12768 19156 12774 19168
rect 13265 19159 13323 19165
rect 13265 19156 13277 19159
rect 12768 19128 13277 19156
rect 12768 19116 12774 19128
rect 13265 19125 13277 19128
rect 13311 19125 13323 19159
rect 13372 19156 13400 19196
rect 13538 19184 13544 19236
rect 13596 19224 13602 19236
rect 13596 19196 14044 19224
rect 13596 19184 13602 19196
rect 14016 19165 14044 19196
rect 14090 19184 14096 19236
rect 14148 19224 14154 19236
rect 14936 19224 14964 19255
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 15160 19264 15301 19292
rect 15160 19252 15166 19264
rect 15289 19261 15301 19264
rect 15335 19261 15347 19295
rect 15930 19292 15936 19304
rect 15891 19264 15936 19292
rect 15289 19255 15347 19261
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 16482 19292 16488 19304
rect 16443 19264 16488 19292
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19292 16911 19295
rect 16942 19292 16948 19304
rect 16899 19264 16948 19292
rect 16899 19261 16911 19264
rect 16853 19255 16911 19261
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19261 17463 19295
rect 17678 19292 17684 19304
rect 17639 19264 17684 19292
rect 17405 19255 17463 19261
rect 17126 19224 17132 19236
rect 14148 19196 14964 19224
rect 17087 19196 17132 19224
rect 14148 19184 14154 19196
rect 17126 19184 17132 19196
rect 17184 19184 17190 19236
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13372 19128 13645 19156
rect 13265 19119 13323 19125
rect 13633 19125 13645 19128
rect 13679 19125 13691 19159
rect 13633 19119 13691 19125
rect 14001 19159 14059 19165
rect 14001 19125 14013 19159
rect 14047 19125 14059 19159
rect 14001 19119 14059 19125
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 14369 19159 14427 19165
rect 14369 19156 14381 19159
rect 14240 19128 14381 19156
rect 14240 19116 14246 19128
rect 14369 19125 14381 19128
rect 14415 19125 14427 19159
rect 14369 19119 14427 19125
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14608 19128 14749 19156
rect 14608 19116 14614 19128
rect 14737 19125 14749 19128
rect 14783 19125 14795 19159
rect 14737 19119 14795 19125
rect 15010 19116 15016 19168
rect 15068 19156 15074 19168
rect 15105 19159 15163 19165
rect 15105 19156 15117 19159
rect 15068 19128 15117 19156
rect 15068 19116 15074 19128
rect 15105 19125 15117 19128
rect 15151 19125 15163 19159
rect 15105 19119 15163 19125
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 15473 19159 15531 19165
rect 15473 19156 15485 19159
rect 15436 19128 15485 19156
rect 15436 19116 15442 19128
rect 15473 19125 15485 19128
rect 15519 19125 15531 19159
rect 15473 19119 15531 19125
rect 16669 19159 16727 19165
rect 16669 19125 16681 19159
rect 16715 19156 16727 19159
rect 16850 19156 16856 19168
rect 16715 19128 16856 19156
rect 16715 19125 16727 19128
rect 16669 19119 16727 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 17420 19156 17448 19255
rect 17678 19252 17684 19264
rect 17736 19252 17742 19304
rect 18322 19292 18328 19304
rect 18235 19264 18328 19292
rect 18322 19252 18328 19264
rect 18380 19292 18386 19304
rect 18782 19292 18788 19304
rect 18380 19264 18788 19292
rect 18380 19252 18386 19264
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 19061 19295 19119 19301
rect 19061 19261 19073 19295
rect 19107 19292 19119 19295
rect 19886 19292 19892 19304
rect 19107 19264 19892 19292
rect 19107 19261 19119 19264
rect 19061 19255 19119 19261
rect 19886 19252 19892 19264
rect 19944 19252 19950 19304
rect 20438 19292 20444 19304
rect 20399 19264 20444 19292
rect 20438 19252 20444 19264
rect 20496 19252 20502 19304
rect 20714 19292 20720 19304
rect 20675 19264 20720 19292
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 18598 19224 18604 19236
rect 18559 19196 18604 19224
rect 18598 19184 18604 19196
rect 18656 19184 18662 19236
rect 19610 19184 19616 19236
rect 19668 19224 19674 19236
rect 19705 19227 19763 19233
rect 19705 19224 19717 19227
rect 19668 19196 19717 19224
rect 19668 19184 19674 19196
rect 19705 19193 19717 19196
rect 19751 19193 19763 19227
rect 19705 19187 19763 19193
rect 19334 19156 19340 19168
rect 17420 19128 19340 19156
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 3050 18952 3056 18964
rect 1728 18924 3056 18952
rect 1728 18912 1734 18924
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 3234 18952 3240 18964
rect 3195 18924 3240 18952
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 3786 18952 3792 18964
rect 3344 18924 3792 18952
rect 934 18844 940 18896
rect 992 18884 998 18896
rect 3344 18884 3372 18924
rect 3786 18912 3792 18924
rect 3844 18912 3850 18964
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 4120 18924 4537 18952
rect 4120 18912 4126 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 5442 18952 5448 18964
rect 5403 18924 5448 18952
rect 4525 18915 4583 18921
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5810 18952 5816 18964
rect 5771 18924 5816 18952
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 5994 18912 6000 18964
rect 6052 18952 6058 18964
rect 9401 18955 9459 18961
rect 9401 18952 9413 18955
rect 6052 18924 9413 18952
rect 6052 18912 6058 18924
rect 9401 18921 9413 18924
rect 9447 18921 9459 18955
rect 9401 18915 9459 18921
rect 9490 18912 9496 18964
rect 9548 18952 9554 18964
rect 11698 18952 11704 18964
rect 9548 18924 11704 18952
rect 9548 18912 9554 18924
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 13446 18952 13452 18964
rect 11808 18924 13452 18952
rect 992 18856 3372 18884
rect 992 18844 998 18856
rect 3418 18844 3424 18896
rect 3476 18884 3482 18896
rect 5166 18884 5172 18896
rect 3476 18856 4936 18884
rect 5127 18856 5172 18884
rect 3476 18844 3482 18856
rect 2406 18776 2412 18828
rect 2464 18816 2470 18828
rect 3145 18819 3203 18825
rect 3145 18816 3157 18819
rect 2464 18788 3157 18816
rect 2464 18776 2470 18788
rect 3145 18785 3157 18788
rect 3191 18816 3203 18819
rect 4062 18816 4068 18828
rect 3191 18788 4068 18816
rect 3191 18785 3203 18788
rect 3145 18779 3203 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 4908 18825 4936 18856
rect 5166 18844 5172 18856
rect 5224 18844 5230 18896
rect 5258 18844 5264 18896
rect 5316 18884 5322 18896
rect 8754 18884 8760 18896
rect 5316 18856 8760 18884
rect 5316 18844 5322 18856
rect 8754 18844 8760 18856
rect 8812 18844 8818 18896
rect 8846 18844 8852 18896
rect 8904 18884 8910 18896
rect 10870 18884 10876 18896
rect 8904 18856 10640 18884
rect 10831 18856 10876 18884
rect 8904 18844 8910 18856
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4893 18819 4951 18825
rect 4479 18788 4844 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 2038 18708 2044 18760
rect 2096 18748 2102 18760
rect 3418 18757 3424 18760
rect 3375 18751 3424 18757
rect 2096 18720 3188 18748
rect 2096 18708 2102 18720
rect 2866 18640 2872 18692
rect 2924 18680 2930 18692
rect 3160 18680 3188 18720
rect 3375 18717 3387 18751
rect 3421 18717 3424 18751
rect 3375 18711 3424 18717
rect 3418 18708 3424 18711
rect 3476 18708 3482 18760
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 4448 18748 4476 18779
rect 3844 18720 4476 18748
rect 4709 18751 4767 18757
rect 3844 18708 3850 18720
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4816 18748 4844 18788
rect 4893 18785 4905 18819
rect 4939 18785 4951 18819
rect 4893 18779 4951 18785
rect 4982 18776 4988 18828
rect 5040 18816 5046 18828
rect 5350 18816 5356 18828
rect 5040 18788 5356 18816
rect 5040 18776 5046 18788
rect 5350 18776 5356 18788
rect 5408 18816 5414 18828
rect 6273 18819 6331 18825
rect 6273 18816 6285 18819
rect 5408 18788 6285 18816
rect 5408 18776 5414 18788
rect 6273 18785 6285 18788
rect 6319 18785 6331 18819
rect 6273 18779 6331 18785
rect 6540 18819 6598 18825
rect 6540 18785 6552 18819
rect 6586 18816 6598 18819
rect 7834 18816 7840 18828
rect 6586 18788 7840 18816
rect 6586 18785 6598 18788
rect 6540 18779 6598 18785
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 8196 18819 8254 18825
rect 8196 18785 8208 18819
rect 8242 18816 8254 18819
rect 9214 18816 9220 18828
rect 8242 18788 9220 18816
rect 8242 18785 8254 18788
rect 8196 18779 8254 18785
rect 9214 18776 9220 18788
rect 9272 18776 9278 18828
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10502 18816 10508 18828
rect 10091 18788 10508 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 10612 18825 10640 18856
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11808 18884 11836 18924
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 16761 18955 16819 18961
rect 16761 18921 16773 18955
rect 16807 18952 16819 18955
rect 17310 18952 17316 18964
rect 16807 18924 17316 18952
rect 16807 18921 16819 18924
rect 16761 18915 16819 18921
rect 17310 18912 17316 18924
rect 17368 18912 17374 18964
rect 19150 18912 19156 18964
rect 19208 18912 19214 18964
rect 19518 18952 19524 18964
rect 19352 18924 19524 18952
rect 11072 18856 11836 18884
rect 10597 18819 10655 18825
rect 10597 18785 10609 18819
rect 10643 18785 10655 18819
rect 10597 18779 10655 18785
rect 10686 18776 10692 18828
rect 10744 18816 10750 18828
rect 11072 18816 11100 18856
rect 12158 18844 12164 18896
rect 12216 18884 12222 18896
rect 13906 18884 13912 18896
rect 12216 18856 13912 18884
rect 12216 18844 12222 18856
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 14553 18887 14611 18893
rect 14553 18853 14565 18887
rect 14599 18884 14611 18887
rect 15102 18884 15108 18896
rect 14599 18856 15108 18884
rect 14599 18853 14611 18856
rect 14553 18847 14611 18853
rect 15102 18844 15108 18856
rect 15160 18844 15166 18896
rect 15565 18887 15623 18893
rect 15565 18853 15577 18887
rect 15611 18884 15623 18887
rect 16482 18884 16488 18896
rect 15611 18856 16488 18884
rect 15611 18853 15623 18856
rect 15565 18847 15623 18853
rect 16482 18844 16488 18856
rect 16540 18844 16546 18896
rect 19168 18884 19196 18912
rect 18524 18856 19196 18884
rect 11606 18825 11612 18828
rect 11600 18816 11612 18825
rect 10744 18788 11100 18816
rect 11567 18788 11612 18816
rect 10744 18776 10750 18788
rect 11600 18779 11612 18788
rect 11606 18776 11612 18779
rect 11664 18776 11670 18828
rect 13072 18819 13130 18825
rect 13072 18816 13084 18819
rect 12728 18788 13084 18816
rect 5258 18748 5264 18760
rect 4816 18720 5264 18748
rect 4709 18711 4767 18717
rect 3234 18680 3240 18692
rect 2924 18652 3004 18680
rect 3160 18652 3240 18680
rect 2924 18640 2930 18652
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 2976 18612 3004 18652
rect 3234 18640 3240 18652
rect 3292 18640 3298 18692
rect 3970 18640 3976 18692
rect 4028 18680 4034 18692
rect 4724 18680 4752 18711
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 5902 18748 5908 18760
rect 5863 18720 5908 18748
rect 5902 18708 5908 18720
rect 5960 18708 5966 18760
rect 6086 18748 6092 18760
rect 5999 18720 6092 18748
rect 6086 18708 6092 18720
rect 6144 18708 6150 18760
rect 7650 18708 7656 18760
rect 7708 18748 7714 18760
rect 7929 18751 7987 18757
rect 7929 18748 7941 18751
rect 7708 18720 7941 18748
rect 7708 18708 7714 18720
rect 7929 18717 7941 18720
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18748 9459 18751
rect 9582 18748 9588 18760
rect 9447 18720 9588 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9582 18708 9588 18720
rect 9640 18748 9646 18760
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 9640 18720 10149 18748
rect 9640 18708 9646 18720
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 11333 18751 11391 18757
rect 11333 18717 11345 18751
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 4982 18680 4988 18692
rect 4028 18652 4988 18680
rect 4028 18640 4034 18652
rect 4982 18640 4988 18652
rect 5040 18680 5046 18692
rect 5626 18680 5632 18692
rect 5040 18652 5632 18680
rect 5040 18640 5046 18652
rect 5626 18640 5632 18652
rect 5684 18640 5690 18692
rect 4065 18615 4123 18621
rect 4065 18612 4077 18615
rect 2832 18584 2877 18612
rect 2976 18584 4077 18612
rect 2832 18572 2838 18584
rect 4065 18581 4077 18584
rect 4111 18581 4123 18615
rect 6104 18612 6132 18708
rect 9214 18640 9220 18692
rect 9272 18680 9278 18692
rect 10244 18680 10272 18711
rect 9272 18652 10272 18680
rect 9272 18640 9278 18652
rect 7653 18615 7711 18621
rect 7653 18612 7665 18615
rect 6104 18584 7665 18612
rect 4065 18575 4123 18581
rect 7653 18581 7665 18584
rect 7699 18581 7711 18615
rect 7653 18575 7711 18581
rect 8662 18572 8668 18624
rect 8720 18612 8726 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 8720 18584 9321 18612
rect 8720 18572 8726 18584
rect 9309 18581 9321 18584
rect 9355 18581 9367 18615
rect 9309 18575 9367 18581
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 9456 18584 9689 18612
rect 9456 18572 9462 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 9677 18575 9735 18581
rect 10778 18572 10784 18624
rect 10836 18612 10842 18624
rect 11348 18612 11376 18711
rect 12728 18689 12756 18788
rect 13072 18785 13084 18788
rect 13118 18816 13130 18819
rect 13814 18816 13820 18828
rect 13118 18788 13820 18816
rect 13118 18785 13130 18788
rect 13072 18779 13130 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 14274 18816 14280 18828
rect 14235 18788 14280 18816
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 15010 18776 15016 18828
rect 15068 18816 15074 18828
rect 15289 18819 15347 18825
rect 15289 18816 15301 18819
rect 15068 18788 15301 18816
rect 15068 18776 15074 18788
rect 15289 18785 15301 18788
rect 15335 18785 15347 18819
rect 15289 18779 15347 18785
rect 16577 18819 16635 18825
rect 16577 18785 16589 18819
rect 16623 18816 16635 18819
rect 16758 18816 16764 18828
rect 16623 18788 16764 18816
rect 16623 18785 16635 18788
rect 16577 18779 16635 18785
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 17957 18819 18015 18825
rect 17957 18785 17969 18819
rect 18003 18816 18015 18819
rect 18322 18816 18328 18828
rect 18003 18788 18328 18816
rect 18003 18785 18015 18788
rect 17957 18779 18015 18785
rect 18322 18776 18328 18788
rect 18380 18776 18386 18828
rect 18524 18825 18552 18856
rect 18509 18819 18567 18825
rect 18509 18785 18521 18819
rect 18555 18785 18567 18819
rect 19153 18819 19211 18825
rect 19153 18816 19165 18819
rect 18509 18779 18567 18785
rect 18800 18788 19165 18816
rect 12805 18751 12863 18757
rect 12805 18717 12817 18751
rect 12851 18717 12863 18751
rect 18138 18748 18144 18760
rect 18099 18720 18144 18748
rect 12805 18711 12863 18717
rect 12713 18683 12771 18689
rect 12713 18649 12725 18683
rect 12759 18649 12771 18683
rect 12713 18643 12771 18649
rect 12820 18612 12848 18711
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18690 18748 18696 18760
rect 18651 18720 18696 18748
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 16942 18640 16948 18692
rect 17000 18680 17006 18692
rect 18800 18680 18828 18788
rect 19153 18785 19165 18788
rect 19199 18816 19211 18819
rect 19352 18816 19380 18924
rect 19518 18912 19524 18924
rect 19576 18952 19582 18964
rect 21082 18952 21088 18964
rect 19576 18924 21088 18952
rect 19576 18912 19582 18924
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 20530 18884 20536 18896
rect 20491 18856 20536 18884
rect 20530 18844 20536 18856
rect 20588 18844 20594 18896
rect 19199 18788 19380 18816
rect 19199 18785 19211 18788
rect 19153 18779 19211 18785
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 19484 18788 19717 18816
rect 19484 18776 19490 18788
rect 19705 18785 19717 18788
rect 19751 18785 19763 18819
rect 19705 18779 19763 18785
rect 19794 18776 19800 18828
rect 19852 18816 19858 18828
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 19852 18788 20269 18816
rect 19852 18776 19858 18788
rect 20257 18785 20269 18788
rect 20303 18785 20315 18819
rect 20257 18779 20315 18785
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 19024 18720 19349 18748
rect 19024 18708 19030 18720
rect 19337 18717 19349 18720
rect 19383 18717 19395 18751
rect 19337 18711 19395 18717
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18717 19947 18751
rect 19889 18711 19947 18717
rect 17000 18652 18828 18680
rect 17000 18640 17006 18652
rect 19058 18640 19064 18692
rect 19116 18680 19122 18692
rect 19904 18680 19932 18711
rect 19116 18652 19932 18680
rect 19116 18640 19122 18652
rect 13446 18612 13452 18624
rect 10836 18584 13452 18612
rect 10836 18572 10842 18584
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 13780 18584 14197 18612
rect 13780 18572 13786 18584
rect 14185 18581 14197 18584
rect 14231 18581 14243 18615
rect 14185 18575 14243 18581
rect 15930 18572 15936 18624
rect 15988 18612 15994 18624
rect 20346 18612 20352 18624
rect 15988 18584 20352 18612
rect 15988 18572 15994 18584
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 2133 18411 2191 18417
rect 2133 18377 2145 18411
rect 2179 18408 2191 18411
rect 4433 18411 4491 18417
rect 4433 18408 4445 18411
rect 2179 18380 2820 18408
rect 2179 18377 2191 18380
rect 2133 18371 2191 18377
rect 1946 18340 1952 18352
rect 1907 18312 1952 18340
rect 1946 18300 1952 18312
rect 2004 18300 2010 18352
rect 2130 18232 2136 18284
rect 2188 18272 2194 18284
rect 2685 18275 2743 18281
rect 2685 18272 2697 18275
rect 2188 18244 2697 18272
rect 2188 18232 2194 18244
rect 2685 18241 2697 18244
rect 2731 18241 2743 18275
rect 2792 18272 2820 18380
rect 2884 18380 4445 18408
rect 2884 18352 2912 18380
rect 4433 18377 4445 18380
rect 4479 18377 4491 18411
rect 4433 18371 4491 18377
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 7285 18411 7343 18417
rect 7285 18408 7297 18411
rect 5960 18380 7297 18408
rect 5960 18368 5966 18380
rect 7285 18377 7297 18380
rect 7331 18377 7343 18411
rect 7285 18371 7343 18377
rect 9217 18411 9275 18417
rect 9217 18377 9229 18411
rect 9263 18408 9275 18411
rect 11146 18408 11152 18420
rect 9263 18380 11152 18408
rect 9263 18377 9275 18380
rect 9217 18371 9275 18377
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 12483 18380 13124 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 2866 18300 2872 18352
rect 2924 18300 2930 18352
rect 4246 18300 4252 18352
rect 4304 18340 4310 18352
rect 4341 18343 4399 18349
rect 4341 18340 4353 18343
rect 4304 18312 4353 18340
rect 4304 18300 4310 18312
rect 4341 18309 4353 18312
rect 4387 18309 4399 18343
rect 4341 18303 4399 18309
rect 4448 18312 10272 18340
rect 2792 18244 3096 18272
rect 2685 18235 2743 18241
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 1765 18167 1823 18173
rect 2501 18207 2559 18213
rect 2501 18173 2513 18207
rect 2547 18204 2559 18207
rect 2866 18204 2872 18216
rect 2547 18176 2872 18204
rect 2547 18173 2559 18176
rect 2501 18167 2559 18173
rect 1780 18136 1808 18167
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18173 3019 18207
rect 3068 18204 3096 18244
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4448 18272 4476 18312
rect 4893 18275 4951 18281
rect 4893 18272 4905 18275
rect 4120 18244 4476 18272
rect 4816 18244 4905 18272
rect 4120 18232 4126 18244
rect 4430 18204 4436 18216
rect 3068 18176 4436 18204
rect 2961 18167 3019 18173
rect 1780 18108 2268 18136
rect 2240 18068 2268 18108
rect 2406 18096 2412 18148
rect 2464 18136 2470 18148
rect 2593 18139 2651 18145
rect 2593 18136 2605 18139
rect 2464 18108 2605 18136
rect 2464 18096 2470 18108
rect 2593 18105 2605 18108
rect 2639 18105 2651 18139
rect 2593 18099 2651 18105
rect 2682 18096 2688 18148
rect 2740 18136 2746 18148
rect 2976 18136 3004 18167
rect 4430 18164 4436 18176
rect 4488 18164 4494 18216
rect 3234 18145 3240 18148
rect 3228 18136 3240 18145
rect 2740 18108 3004 18136
rect 3195 18108 3240 18136
rect 2740 18096 2746 18108
rect 3228 18099 3240 18108
rect 3234 18096 3240 18099
rect 3292 18096 3298 18148
rect 3694 18096 3700 18148
rect 3752 18136 3758 18148
rect 4706 18136 4712 18148
rect 3752 18108 4712 18136
rect 3752 18096 3758 18108
rect 4706 18096 4712 18108
rect 4764 18136 4770 18148
rect 4816 18136 4844 18244
rect 4893 18241 4905 18244
rect 4939 18241 4951 18275
rect 4893 18235 4951 18241
rect 4982 18232 4988 18284
rect 5040 18272 5046 18284
rect 5040 18244 5085 18272
rect 5040 18232 5046 18244
rect 5718 18204 5724 18216
rect 4764 18108 4844 18136
rect 5000 18176 5724 18204
rect 4764 18096 4770 18108
rect 2866 18068 2872 18080
rect 2240 18040 2872 18068
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 3050 18028 3056 18080
rect 3108 18068 3114 18080
rect 4801 18071 4859 18077
rect 4801 18068 4813 18071
rect 3108 18040 4813 18068
rect 3108 18028 3114 18040
rect 4801 18037 4813 18040
rect 4847 18068 4859 18071
rect 5000 18068 5028 18176
rect 5718 18164 5724 18176
rect 5776 18204 5782 18216
rect 6089 18207 6147 18213
rect 6089 18204 6101 18207
rect 5776 18176 6101 18204
rect 5776 18164 5782 18176
rect 6089 18173 6101 18176
rect 6135 18173 6147 18207
rect 6089 18167 6147 18173
rect 5997 18139 6055 18145
rect 5997 18105 6009 18139
rect 6043 18136 6055 18139
rect 6196 18136 6224 18312
rect 6273 18275 6331 18281
rect 6273 18241 6285 18275
rect 6319 18272 6331 18275
rect 6454 18272 6460 18284
rect 6319 18244 6460 18272
rect 6319 18241 6331 18244
rect 6273 18235 6331 18241
rect 6454 18232 6460 18244
rect 6512 18232 6518 18284
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8570 18272 8576 18284
rect 8531 18244 8576 18272
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 8662 18232 8668 18284
rect 8720 18272 8726 18284
rect 9858 18272 9864 18284
rect 8720 18244 8765 18272
rect 9819 18244 9864 18272
rect 8720 18232 8726 18244
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10244 18272 10272 18312
rect 11238 18300 11244 18352
rect 11296 18340 11302 18352
rect 12986 18340 12992 18352
rect 11296 18312 12992 18340
rect 11296 18300 11302 18312
rect 12986 18300 12992 18312
rect 13044 18300 13050 18352
rect 13096 18340 13124 18380
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 13265 18411 13323 18417
rect 13265 18408 13277 18411
rect 13228 18380 13277 18408
rect 13228 18368 13234 18380
rect 13265 18377 13277 18380
rect 13311 18377 13323 18411
rect 13265 18371 13323 18377
rect 17221 18411 17279 18417
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 17586 18408 17592 18420
rect 17267 18380 17592 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 22554 18340 22560 18352
rect 13096 18312 13400 18340
rect 10244 18244 10364 18272
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18204 8539 18207
rect 9398 18204 9404 18216
rect 8527 18176 9404 18204
rect 8527 18173 8539 18176
rect 8481 18167 8539 18173
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9582 18204 9588 18216
rect 9543 18176 9588 18204
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 9732 18176 10241 18204
rect 9732 18164 9738 18176
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 6043 18108 6224 18136
rect 7653 18139 7711 18145
rect 6043 18105 6055 18108
rect 5997 18099 6055 18105
rect 7653 18105 7665 18139
rect 7699 18136 7711 18139
rect 9766 18136 9772 18148
rect 7699 18108 9772 18136
rect 7699 18105 7711 18108
rect 7653 18099 7711 18105
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 5626 18068 5632 18080
rect 4847 18040 5028 18068
rect 5587 18040 5632 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 7745 18071 7803 18077
rect 7745 18037 7757 18071
rect 7791 18068 7803 18071
rect 8113 18071 8171 18077
rect 8113 18068 8125 18071
rect 7791 18040 8125 18068
rect 7791 18037 7803 18040
rect 7745 18031 7803 18037
rect 8113 18037 8125 18040
rect 8159 18037 8171 18071
rect 8113 18031 8171 18037
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 9677 18071 9735 18077
rect 9677 18068 9689 18071
rect 8812 18040 9689 18068
rect 8812 18028 8818 18040
rect 9677 18037 9689 18040
rect 9723 18037 9735 18071
rect 10336 18068 10364 18244
rect 11606 18232 11612 18284
rect 11664 18272 11670 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 11664 18244 13093 18272
rect 11664 18232 11670 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 11112 18176 12909 18204
rect 11112 18164 11118 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 13372 18204 13400 18312
rect 19628 18312 22560 18340
rect 13814 18272 13820 18284
rect 13775 18244 13820 18272
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 19628 18281 19656 18312
rect 22554 18300 22560 18312
rect 22612 18300 22618 18352
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20717 18275 20775 18281
rect 20312 18244 20484 18272
rect 20312 18232 20318 18244
rect 13725 18207 13783 18213
rect 13725 18204 13737 18207
rect 13372 18176 13737 18204
rect 12897 18167 12955 18173
rect 13725 18173 13737 18176
rect 13771 18173 13783 18207
rect 13725 18167 13783 18173
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18204 17095 18207
rect 17494 18204 17500 18216
rect 17083 18176 17500 18204
rect 17083 18173 17095 18176
rect 17037 18167 17095 18173
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 19518 18204 19524 18216
rect 19383 18176 19524 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 19518 18164 19524 18176
rect 19576 18164 19582 18216
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18204 19947 18207
rect 20346 18204 20352 18216
rect 19935 18176 20352 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 20346 18164 20352 18176
rect 20404 18164 20410 18216
rect 20456 18213 20484 18244
rect 20717 18241 20729 18275
rect 20763 18272 20775 18275
rect 20806 18272 20812 18284
rect 20763 18244 20812 18272
rect 20763 18241 20775 18244
rect 20717 18235 20775 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 20441 18207 20499 18213
rect 20441 18173 20453 18207
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 10496 18139 10554 18145
rect 10496 18105 10508 18139
rect 10542 18136 10554 18139
rect 10962 18136 10968 18148
rect 10542 18108 10968 18136
rect 10542 18105 10554 18108
rect 10496 18099 10554 18105
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 12250 18136 12256 18148
rect 11072 18108 12256 18136
rect 11072 18068 11100 18108
rect 12250 18096 12256 18108
rect 12308 18096 12314 18148
rect 12986 18096 12992 18148
rect 13044 18136 13050 18148
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 13044 18108 13645 18136
rect 13044 18096 13050 18108
rect 13633 18105 13645 18108
rect 13679 18105 13691 18139
rect 13633 18099 13691 18105
rect 19978 18096 19984 18148
rect 20036 18136 20042 18148
rect 20165 18139 20223 18145
rect 20165 18136 20177 18139
rect 20036 18108 20177 18136
rect 20036 18096 20042 18108
rect 20165 18105 20177 18108
rect 20211 18105 20223 18139
rect 20165 18099 20223 18105
rect 10336 18040 11100 18068
rect 9677 18031 9735 18037
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11606 18068 11612 18080
rect 11480 18040 11612 18068
rect 11480 18028 11486 18040
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 11790 18028 11796 18080
rect 11848 18068 11854 18080
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 11848 18040 12817 18068
rect 11848 18028 11854 18040
rect 12805 18037 12817 18040
rect 12851 18037 12863 18071
rect 12805 18031 12863 18037
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 5442 17864 5448 17876
rect 4948 17836 5448 17864
rect 4948 17824 4954 17836
rect 5442 17824 5448 17836
rect 5500 17864 5506 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 5500 17836 6469 17864
rect 5500 17824 5506 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 6457 17827 6515 17833
rect 7193 17867 7251 17873
rect 7193 17833 7205 17867
rect 7239 17864 7251 17867
rect 7282 17864 7288 17876
rect 7239 17836 7288 17864
rect 7239 17833 7251 17836
rect 7193 17827 7251 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 8021 17867 8079 17873
rect 8021 17833 8033 17867
rect 8067 17864 8079 17867
rect 8202 17864 8208 17876
rect 8067 17836 8208 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 10965 17867 11023 17873
rect 10965 17833 10977 17867
rect 11011 17864 11023 17867
rect 11054 17864 11060 17876
rect 11011 17836 11060 17864
rect 11011 17833 11023 17836
rect 10965 17827 11023 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 11425 17867 11483 17873
rect 11425 17864 11437 17867
rect 11204 17836 11437 17864
rect 11204 17824 11210 17836
rect 11425 17833 11437 17836
rect 11471 17833 11483 17867
rect 11425 17827 11483 17833
rect 11606 17824 11612 17876
rect 11664 17864 11670 17876
rect 11882 17864 11888 17876
rect 11664 17836 11888 17864
rect 11664 17824 11670 17836
rect 11882 17824 11888 17836
rect 11940 17824 11946 17876
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12308 17836 13001 17864
rect 12308 17824 12314 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 21082 17864 21088 17876
rect 21043 17836 21088 17864
rect 12989 17827 13047 17833
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 2130 17805 2136 17808
rect 2124 17796 2136 17805
rect 2091 17768 2136 17796
rect 2124 17759 2136 17768
rect 2130 17756 2136 17759
rect 2188 17756 2194 17808
rect 2866 17756 2872 17808
rect 2924 17796 2930 17808
rect 4062 17796 4068 17808
rect 2924 17768 4068 17796
rect 2924 17756 2930 17768
rect 4062 17756 4068 17768
rect 4120 17756 4126 17808
rect 4246 17756 4252 17808
rect 4304 17796 4310 17808
rect 4770 17799 4828 17805
rect 4770 17796 4782 17799
rect 4304 17768 4782 17796
rect 4304 17756 4310 17768
rect 4770 17765 4782 17768
rect 4816 17765 4828 17799
rect 4770 17759 4828 17765
rect 5258 17756 5264 17808
rect 5316 17796 5322 17808
rect 6365 17799 6423 17805
rect 6365 17796 6377 17799
rect 5316 17768 6377 17796
rect 5316 17756 5322 17768
rect 6365 17765 6377 17768
rect 6411 17796 6423 17799
rect 9674 17796 9680 17808
rect 6411 17768 9680 17796
rect 6411 17765 6423 17768
rect 6365 17759 6423 17765
rect 9674 17756 9680 17768
rect 9732 17756 9738 17808
rect 9858 17756 9864 17808
rect 9916 17796 9922 17808
rect 11974 17796 11980 17808
rect 9916 17768 11980 17796
rect 9916 17756 9922 17768
rect 11974 17756 11980 17768
rect 12032 17796 12038 17808
rect 12032 17768 12296 17796
rect 12032 17756 12038 17768
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17697 1547 17731
rect 1489 17691 1547 17697
rect 1857 17731 1915 17737
rect 1857 17697 1869 17731
rect 1903 17728 1915 17731
rect 2406 17728 2412 17740
rect 1903 17700 2412 17728
rect 1903 17697 1915 17700
rect 1857 17691 1915 17697
rect 1504 17592 1532 17691
rect 2406 17688 2412 17700
rect 2464 17728 2470 17740
rect 2682 17728 2688 17740
rect 2464 17700 2688 17728
rect 2464 17688 2470 17700
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 7561 17731 7619 17737
rect 3068 17700 6224 17728
rect 1504 17564 1900 17592
rect 1872 17524 1900 17564
rect 3068 17524 3096 17700
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4522 17660 4528 17672
rect 4120 17632 4528 17660
rect 4120 17620 4126 17632
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 5534 17552 5540 17604
rect 5592 17592 5598 17604
rect 6086 17592 6092 17604
rect 5592 17564 6092 17592
rect 5592 17552 5598 17564
rect 6086 17552 6092 17564
rect 6144 17552 6150 17604
rect 3234 17524 3240 17536
rect 1872 17496 3096 17524
rect 3147 17496 3240 17524
rect 3234 17484 3240 17496
rect 3292 17524 3298 17536
rect 5166 17524 5172 17536
rect 3292 17496 5172 17524
rect 3292 17484 3298 17496
rect 5166 17484 5172 17496
rect 5224 17484 5230 17536
rect 5902 17524 5908 17536
rect 5863 17496 5908 17524
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 6196 17524 6224 17700
rect 7561 17697 7573 17731
rect 7607 17728 7619 17731
rect 8110 17728 8116 17740
rect 7607 17700 8116 17728
rect 7607 17697 7619 17700
rect 7561 17691 7619 17697
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17728 8447 17731
rect 8570 17728 8576 17740
rect 8435 17700 8576 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 11146 17728 11152 17740
rect 10551 17700 11152 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 12158 17728 12164 17740
rect 11379 17700 12020 17728
rect 12119 17700 12164 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 6454 17620 6460 17672
rect 6512 17660 6518 17672
rect 6549 17663 6607 17669
rect 6549 17660 6561 17663
rect 6512 17632 6561 17660
rect 6512 17620 6518 17632
rect 6549 17629 6561 17632
rect 6595 17629 6607 17663
rect 6549 17623 6607 17629
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17660 7711 17663
rect 7742 17660 7748 17672
rect 7699 17632 7748 17660
rect 7699 17629 7711 17632
rect 7653 17623 7711 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17629 7895 17663
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 7837 17623 7895 17629
rect 7852 17592 7880 17623
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8662 17660 8668 17672
rect 8623 17632 8668 17660
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 11422 17660 11428 17672
rect 10827 17632 11428 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 11517 17663 11575 17669
rect 11517 17629 11529 17663
rect 11563 17629 11575 17663
rect 11992 17660 12020 17700
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 12268 17728 12296 17768
rect 12342 17756 12348 17808
rect 12400 17796 12406 17808
rect 13081 17799 13139 17805
rect 13081 17796 13093 17799
rect 12400 17768 13093 17796
rect 12400 17756 12406 17768
rect 13081 17765 13093 17768
rect 13127 17765 13139 17799
rect 13081 17759 13139 17765
rect 18690 17756 18696 17808
rect 18748 17796 18754 17808
rect 18748 17768 20944 17796
rect 18748 17756 18754 17768
rect 13722 17737 13728 17740
rect 13716 17728 13728 17737
rect 12268 17700 12388 17728
rect 12066 17660 12072 17672
rect 11992 17632 12072 17660
rect 11517 17623 11575 17629
rect 8680 17592 8708 17620
rect 7852 17564 8708 17592
rect 10137 17595 10195 17601
rect 10137 17561 10149 17595
rect 10183 17592 10195 17595
rect 11238 17592 11244 17604
rect 10183 17564 11244 17592
rect 10183 17561 10195 17564
rect 10137 17555 10195 17561
rect 11238 17552 11244 17564
rect 11296 17552 11302 17604
rect 8754 17524 8760 17536
rect 6052 17496 6097 17524
rect 6196 17496 8760 17524
rect 6052 17484 6058 17496
rect 8754 17484 8760 17496
rect 8812 17524 8818 17536
rect 10870 17524 10876 17536
rect 8812 17496 10876 17524
rect 8812 17484 8818 17496
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11532 17524 11560 17623
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12250 17660 12256 17672
rect 12211 17632 12256 17660
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 12360 17669 12388 17700
rect 13280 17700 13728 17728
rect 13280 17669 13308 17700
rect 13716 17691 13728 17700
rect 13722 17688 13728 17691
rect 13780 17688 13786 17740
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 20916 17737 20944 17768
rect 20257 17731 20315 17737
rect 20257 17728 20269 17731
rect 19852 17700 20269 17728
rect 19852 17688 19858 17700
rect 20257 17697 20269 17700
rect 20303 17697 20315 17731
rect 20257 17691 20315 17697
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17629 13323 17663
rect 13446 17660 13452 17672
rect 13407 17632 13452 17660
rect 13265 17623 13323 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17660 20591 17663
rect 21358 17660 21364 17672
rect 20579 17632 21364 17660
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 20898 17592 20904 17604
rect 14608 17564 20904 17592
rect 14608 17552 14614 17564
rect 20898 17552 20904 17564
rect 20956 17552 20962 17604
rect 11020 17496 11560 17524
rect 11793 17527 11851 17533
rect 11020 17484 11026 17496
rect 11793 17493 11805 17527
rect 11839 17524 11851 17527
rect 11882 17524 11888 17536
rect 11839 17496 11888 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 12618 17524 12624 17536
rect 12579 17496 12624 17524
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 14829 17527 14887 17533
rect 14829 17524 14841 17527
rect 14516 17496 14841 17524
rect 14516 17484 14522 17496
rect 14829 17493 14841 17496
rect 14875 17493 14887 17527
rect 14829 17487 14887 17493
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4617 17323 4675 17329
rect 4617 17320 4629 17323
rect 4212 17292 4629 17320
rect 4212 17280 4218 17292
rect 4617 17289 4629 17292
rect 4663 17289 4675 17323
rect 4617 17283 4675 17289
rect 4798 17280 4804 17332
rect 4856 17320 4862 17332
rect 6822 17320 6828 17332
rect 4856 17292 6224 17320
rect 6783 17292 6828 17320
rect 4856 17280 4862 17292
rect 2133 17255 2191 17261
rect 2133 17221 2145 17255
rect 2179 17252 2191 17255
rect 3326 17252 3332 17264
rect 2179 17224 3332 17252
rect 2179 17221 2191 17224
rect 2133 17215 2191 17221
rect 3326 17212 3332 17224
rect 3384 17212 3390 17264
rect 3418 17212 3424 17264
rect 3476 17252 3482 17264
rect 3476 17224 3556 17252
rect 3476 17212 3482 17224
rect 2222 17144 2228 17196
rect 2280 17184 2286 17196
rect 3528 17193 3556 17224
rect 3878 17212 3884 17264
rect 3936 17252 3942 17264
rect 5258 17252 5264 17264
rect 3936 17224 5264 17252
rect 3936 17212 3942 17224
rect 5258 17212 5264 17224
rect 5316 17212 5322 17264
rect 5534 17212 5540 17264
rect 5592 17252 5598 17264
rect 6196 17252 6224 17292
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 8389 17323 8447 17329
rect 8389 17289 8401 17323
rect 8435 17320 8447 17323
rect 8478 17320 8484 17332
rect 8435 17292 8484 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 10686 17320 10692 17332
rect 8588 17292 10692 17320
rect 8588 17252 8616 17292
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 10962 17320 10968 17332
rect 10923 17292 10968 17320
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 11425 17323 11483 17329
rect 11425 17289 11437 17323
rect 11471 17320 11483 17323
rect 11790 17320 11796 17332
rect 11471 17292 11796 17320
rect 11471 17289 11483 17292
rect 11425 17283 11483 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12299 17292 12747 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 5592 17224 6132 17252
rect 6196 17224 8616 17252
rect 5592 17212 5598 17224
rect 2685 17187 2743 17193
rect 2685 17184 2697 17187
rect 2280 17156 2697 17184
rect 2280 17144 2286 17156
rect 2685 17153 2697 17156
rect 2731 17184 2743 17187
rect 3513 17187 3571 17193
rect 2731 17156 3464 17184
rect 2731 17153 2743 17156
rect 2685 17147 2743 17153
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 2774 17116 2780 17128
rect 2639 17088 2780 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 3436 17116 3464 17156
rect 3513 17153 3525 17187
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 3694 17144 3700 17196
rect 3752 17184 3758 17196
rect 4341 17187 4399 17193
rect 4341 17184 4353 17187
rect 3752 17156 4353 17184
rect 3752 17144 3758 17156
rect 4341 17153 4353 17156
rect 4387 17153 4399 17187
rect 5166 17184 5172 17196
rect 5127 17156 5172 17184
rect 4341 17147 4399 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5994 17184 6000 17196
rect 5955 17156 6000 17184
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 6104 17193 6132 17224
rect 8938 17212 8944 17264
rect 8996 17252 9002 17264
rect 9490 17252 9496 17264
rect 8996 17224 9496 17252
rect 8996 17212 9002 17224
rect 9490 17212 9496 17224
rect 9548 17212 9554 17264
rect 10980 17252 11008 17280
rect 11514 17252 11520 17264
rect 10980 17224 11520 17252
rect 11514 17212 11520 17224
rect 11572 17252 11578 17264
rect 12437 17255 12495 17261
rect 11572 17224 12020 17252
rect 11572 17212 11578 17224
rect 6089 17187 6147 17193
rect 6089 17153 6101 17187
rect 6135 17153 6147 17187
rect 7466 17184 7472 17196
rect 7427 17156 7472 17184
rect 6089 17147 6147 17153
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 8110 17184 8116 17196
rect 8071 17156 8116 17184
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 9033 17187 9091 17193
rect 9033 17153 9045 17187
rect 9079 17184 9091 17187
rect 9214 17184 9220 17196
rect 9079 17156 9220 17184
rect 9079 17153 9091 17156
rect 9033 17147 9091 17153
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9582 17184 9588 17196
rect 9543 17156 9588 17184
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 11882 17184 11888 17196
rect 11843 17156 11888 17184
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 11992 17193 12020 17224
rect 12437 17221 12449 17255
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 3712 17116 3740 17144
rect 3436 17088 3740 17116
rect 4080 17088 4660 17116
rect 2501 17051 2559 17057
rect 2501 17017 2513 17051
rect 2547 17048 2559 17051
rect 2547 17020 3004 17048
rect 2547 17017 2559 17020
rect 2501 17011 2559 17017
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 2682 16980 2688 16992
rect 1912 16952 2688 16980
rect 1912 16940 1918 16952
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 2976 16989 3004 17020
rect 3050 17008 3056 17060
rect 3108 17048 3114 17060
rect 3421 17051 3479 17057
rect 3421 17048 3433 17051
rect 3108 17020 3433 17048
rect 3108 17008 3114 17020
rect 3421 17017 3433 17020
rect 3467 17048 3479 17051
rect 4080 17048 4108 17088
rect 3467 17020 4108 17048
rect 4157 17051 4215 17057
rect 3467 17017 3479 17020
rect 3421 17011 3479 17017
rect 4157 17017 4169 17051
rect 4203 17048 4215 17051
rect 4522 17048 4528 17060
rect 4203 17020 4528 17048
rect 4203 17017 4215 17020
rect 4157 17011 4215 17017
rect 4522 17008 4528 17020
rect 4580 17008 4586 17060
rect 2961 16983 3019 16989
rect 2961 16949 2973 16983
rect 3007 16949 3019 16983
rect 3326 16980 3332 16992
rect 3287 16952 3332 16980
rect 2961 16943 3019 16949
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 3786 16980 3792 16992
rect 3747 16952 3792 16980
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 4246 16980 4252 16992
rect 4207 16952 4252 16980
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 4632 16980 4660 17088
rect 4890 17076 4896 17128
rect 4948 17116 4954 17128
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4948 17088 4997 17116
rect 4948 17076 4954 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5626 17076 5632 17128
rect 5684 17116 5690 17128
rect 9858 17125 9864 17128
rect 5905 17119 5963 17125
rect 5905 17116 5917 17119
rect 5684 17088 5917 17116
rect 5684 17076 5690 17088
rect 5905 17085 5917 17088
rect 5951 17085 5963 17119
rect 9852 17116 9864 17125
rect 5905 17079 5963 17085
rect 6104 17088 9444 17116
rect 9819 17088 9864 17116
rect 4706 17008 4712 17060
rect 4764 17048 4770 17060
rect 5077 17051 5135 17057
rect 5077 17048 5089 17051
rect 4764 17020 5089 17048
rect 4764 17008 4770 17020
rect 5077 17017 5089 17020
rect 5123 17017 5135 17051
rect 6104 17048 6132 17088
rect 5077 17011 5135 17017
rect 5460 17020 6132 17048
rect 5460 16980 5488 17020
rect 6178 17008 6184 17060
rect 6236 17048 6242 17060
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 6236 17020 7297 17048
rect 6236 17008 6242 17020
rect 7285 17017 7297 17020
rect 7331 17017 7343 17051
rect 9416 17048 9444 17088
rect 9852 17079 9864 17088
rect 9858 17076 9864 17079
rect 9916 17076 9922 17128
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11698 17116 11704 17128
rect 11195 17088 11704 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 11698 17076 11704 17088
rect 11756 17076 11762 17128
rect 12452 17116 12480 17215
rect 12719 17116 12747 17292
rect 12986 17280 12992 17332
rect 13044 17320 13050 17332
rect 15838 17320 15844 17332
rect 13044 17292 15844 17320
rect 13044 17280 13050 17292
rect 15838 17280 15844 17292
rect 15896 17280 15902 17332
rect 19886 17320 19892 17332
rect 19847 17292 19892 17320
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 20254 17320 20260 17332
rect 20215 17292 20260 17320
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 21174 17320 21180 17332
rect 21135 17292 21180 17320
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 12894 17184 12900 17196
rect 12855 17156 12900 17184
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13078 17184 13084 17196
rect 12991 17156 13084 17184
rect 13078 17144 13084 17156
rect 13136 17184 13142 17196
rect 13136 17156 13400 17184
rect 13136 17144 13142 17156
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 11808 17088 12204 17116
rect 12452 17088 12664 17116
rect 12719 17088 12817 17116
rect 10502 17048 10508 17060
rect 9416 17020 10508 17048
rect 7285 17011 7343 17017
rect 10502 17008 10508 17020
rect 10560 17048 10566 17060
rect 11808 17057 11836 17088
rect 11793 17051 11851 17057
rect 10560 17020 11560 17048
rect 10560 17008 10566 17020
rect 4632 16952 5488 16980
rect 5537 16983 5595 16989
rect 5537 16949 5549 16983
rect 5583 16980 5595 16983
rect 6638 16980 6644 16992
rect 5583 16952 6644 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7193 16983 7251 16989
rect 7193 16980 7205 16983
rect 6972 16952 7205 16980
rect 6972 16940 6978 16952
rect 7193 16949 7205 16952
rect 7239 16949 7251 16983
rect 8754 16980 8760 16992
rect 8715 16952 8760 16980
rect 7193 16943 7251 16949
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 8849 16983 8907 16989
rect 8849 16949 8861 16983
rect 8895 16980 8907 16983
rect 8938 16980 8944 16992
rect 8895 16952 8944 16980
rect 8895 16949 8907 16952
rect 8849 16943 8907 16949
rect 8938 16940 8944 16952
rect 8996 16980 9002 16992
rect 11422 16980 11428 16992
rect 8996 16952 11428 16980
rect 8996 16940 9002 16952
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 11532 16980 11560 17020
rect 11793 17017 11805 17051
rect 11839 17017 11851 17051
rect 12176 17048 12204 17088
rect 12526 17048 12532 17060
rect 12176 17020 12532 17048
rect 11793 17011 11851 17017
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12253 16983 12311 16989
rect 12253 16980 12265 16983
rect 11532 16952 12265 16980
rect 12253 16949 12265 16952
rect 12299 16949 12311 16983
rect 12253 16943 12311 16949
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12636 16980 12664 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 13262 17116 13268 17128
rect 13223 17088 13268 17116
rect 12805 17079 12863 17085
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 13372 17116 13400 17156
rect 14292 17156 14872 17184
rect 14292 17116 14320 17156
rect 13372 17088 14320 17116
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17085 14795 17119
rect 14844 17116 14872 17156
rect 19426 17144 19432 17196
rect 19484 17184 19490 17196
rect 19484 17156 20484 17184
rect 19484 17144 19490 17156
rect 16666 17116 16672 17128
rect 14844 17088 16672 17116
rect 14737 17079 14795 17085
rect 13532 17051 13590 17057
rect 13532 17017 13544 17051
rect 13578 17048 13590 17051
rect 14458 17048 14464 17060
rect 13578 17020 14464 17048
rect 13578 17017 13590 17020
rect 13532 17011 13590 17017
rect 14458 17008 14464 17020
rect 14516 17008 14522 17060
rect 12492 16952 12664 16980
rect 12492 16940 12498 16952
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 14274 16980 14280 16992
rect 12952 16952 14280 16980
rect 12952 16940 12958 16952
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 14645 16983 14703 16989
rect 14645 16980 14657 16983
rect 14608 16952 14657 16980
rect 14608 16940 14614 16952
rect 14645 16949 14657 16952
rect 14691 16949 14703 16983
rect 14752 16980 14780 17079
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 14826 17008 14832 17060
rect 14884 17048 14890 17060
rect 14982 17051 15040 17057
rect 14982 17048 14994 17051
rect 14884 17020 14994 17048
rect 14884 17008 14890 17020
rect 14982 17017 14994 17020
rect 15028 17017 15040 17051
rect 14982 17011 15040 17017
rect 19426 17008 19432 17060
rect 19484 17048 19490 17060
rect 19720 17048 19748 17079
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 20456 17125 20484 17156
rect 20073 17119 20131 17125
rect 20073 17116 20085 17119
rect 19852 17088 20085 17116
rect 19852 17076 19858 17088
rect 20073 17085 20085 17088
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17085 20499 17119
rect 20441 17079 20499 17085
rect 20622 17076 20628 17128
rect 20680 17116 20686 17128
rect 20993 17119 21051 17125
rect 20993 17116 21005 17119
rect 20680 17088 21005 17116
rect 20680 17076 20686 17088
rect 20993 17085 21005 17088
rect 21039 17085 21051 17119
rect 20993 17079 21051 17085
rect 19484 17020 19748 17048
rect 20717 17051 20775 17057
rect 19484 17008 19490 17020
rect 20717 17017 20729 17051
rect 20763 17048 20775 17051
rect 21266 17048 21272 17060
rect 20763 17020 21272 17048
rect 20763 17017 20775 17020
rect 20717 17011 20775 17017
rect 21266 17008 21272 17020
rect 21324 17008 21330 17060
rect 15194 16980 15200 16992
rect 14752 16952 15200 16980
rect 14645 16943 14703 16949
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 16114 16980 16120 16992
rect 16075 16952 16120 16980
rect 16114 16940 16120 16952
rect 16172 16940 16178 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 1765 16779 1823 16785
rect 1765 16745 1777 16779
rect 1811 16776 1823 16779
rect 1854 16776 1860 16788
rect 1811 16748 1860 16776
rect 1811 16745 1823 16748
rect 1765 16739 1823 16745
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2133 16779 2191 16785
rect 2133 16745 2145 16779
rect 2179 16776 2191 16779
rect 2593 16779 2651 16785
rect 2593 16776 2605 16779
rect 2179 16748 2605 16776
rect 2179 16745 2191 16748
rect 2133 16739 2191 16745
rect 2593 16745 2605 16748
rect 2639 16745 2651 16779
rect 3602 16776 3608 16788
rect 3563 16748 3608 16776
rect 2593 16739 2651 16745
rect 3602 16736 3608 16748
rect 3660 16736 3666 16788
rect 4522 16776 4528 16788
rect 4483 16748 4528 16776
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 5718 16776 5724 16788
rect 5679 16748 5724 16776
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 6178 16776 6184 16788
rect 6139 16748 6184 16776
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 6638 16776 6644 16788
rect 6599 16748 6644 16776
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 8665 16779 8723 16785
rect 8665 16745 8677 16779
rect 8711 16776 8723 16779
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 8711 16748 10057 16776
rect 8711 16745 8723 16748
rect 8665 16739 8723 16745
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 10045 16739 10103 16745
rect 10594 16736 10600 16788
rect 10652 16776 10658 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 10652 16748 10885 16776
rect 10652 16736 10658 16748
rect 10873 16745 10885 16748
rect 10919 16745 10931 16779
rect 11330 16776 11336 16788
rect 10873 16739 10931 16745
rect 10980 16748 11336 16776
rect 2225 16711 2283 16717
rect 2225 16677 2237 16711
rect 2271 16708 2283 16711
rect 3786 16708 3792 16720
rect 2271 16680 3792 16708
rect 2271 16677 2283 16680
rect 2225 16671 2283 16677
rect 3786 16668 3792 16680
rect 3844 16668 3850 16720
rect 4893 16711 4951 16717
rect 4893 16677 4905 16711
rect 4939 16708 4951 16711
rect 4982 16708 4988 16720
rect 4939 16680 4988 16708
rect 4939 16677 4951 16680
rect 4893 16671 4951 16677
rect 4982 16668 4988 16680
rect 5040 16668 5046 16720
rect 7650 16708 7656 16720
rect 7208 16680 7656 16708
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2682 16640 2688 16652
rect 1443 16612 2688 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2682 16600 2688 16612
rect 2740 16600 2746 16652
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2832 16612 2973 16640
rect 2832 16600 2838 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3421 16643 3479 16649
rect 3421 16609 3433 16643
rect 3467 16640 3479 16643
rect 3467 16612 5396 16640
rect 3467 16609 3479 16612
rect 3421 16603 3479 16609
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 3050 16572 3056 16584
rect 2455 16544 2912 16572
rect 3011 16544 3056 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2884 16504 2912 16544
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 3694 16572 3700 16584
rect 3283 16544 3700 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 3694 16532 3700 16544
rect 3752 16532 3758 16584
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 4985 16575 5043 16581
rect 4985 16572 4997 16575
rect 4856 16544 4997 16572
rect 4856 16532 4862 16544
rect 4985 16541 4997 16544
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 5077 16575 5135 16581
rect 5077 16541 5089 16575
rect 5123 16541 5135 16575
rect 5368 16572 5396 16612
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 5813 16643 5871 16649
rect 5813 16640 5825 16643
rect 5500 16612 5825 16640
rect 5500 16600 5506 16612
rect 5813 16609 5825 16612
rect 5859 16609 5871 16643
rect 6546 16640 6552 16652
rect 6507 16612 6552 16640
rect 5813 16603 5871 16609
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 7208 16649 7236 16680
rect 7650 16668 7656 16680
rect 7708 16668 7714 16720
rect 9033 16711 9091 16717
rect 9033 16677 9045 16711
rect 9079 16708 9091 16711
rect 10980 16708 11008 16748
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 11701 16779 11759 16785
rect 11701 16776 11713 16779
rect 11615 16748 11713 16776
rect 9079 16680 11008 16708
rect 9079 16677 9091 16680
rect 9033 16671 9091 16677
rect 11146 16668 11152 16720
rect 11204 16708 11210 16720
rect 11615 16708 11643 16748
rect 11701 16745 11713 16748
rect 11747 16745 11759 16779
rect 11701 16739 11759 16745
rect 11790 16736 11796 16788
rect 11848 16776 11854 16788
rect 12069 16779 12127 16785
rect 12069 16776 12081 16779
rect 11848 16748 12081 16776
rect 11848 16736 11854 16748
rect 12069 16745 12081 16748
rect 12115 16745 12127 16779
rect 12069 16739 12127 16745
rect 12621 16779 12679 16785
rect 12621 16745 12633 16779
rect 12667 16776 12679 16779
rect 12894 16776 12900 16788
rect 12667 16748 12900 16776
rect 12667 16745 12679 16748
rect 12621 16739 12679 16745
rect 12894 16736 12900 16748
rect 12952 16736 12958 16788
rect 13081 16779 13139 16785
rect 13081 16745 13093 16779
rect 13127 16776 13139 16779
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 13127 16748 13461 16776
rect 13127 16745 13139 16748
rect 13081 16739 13139 16745
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13449 16739 13507 16745
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 14737 16779 14795 16785
rect 14737 16776 14749 16779
rect 13596 16748 14749 16776
rect 13596 16736 13602 16748
rect 14737 16745 14749 16748
rect 14783 16745 14795 16779
rect 14737 16739 14795 16745
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 16945 16779 17003 16785
rect 16945 16776 16957 16779
rect 16632 16748 16957 16776
rect 16632 16736 16638 16748
rect 16945 16745 16957 16748
rect 16991 16745 17003 16779
rect 21082 16776 21088 16788
rect 21043 16748 21088 16776
rect 16945 16739 17003 16745
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 11204 16680 11643 16708
rect 12989 16711 13047 16717
rect 11204 16668 11210 16680
rect 12989 16677 13001 16711
rect 13035 16708 13047 16711
rect 14274 16708 14280 16720
rect 13035 16680 14280 16708
rect 13035 16677 13047 16680
rect 12989 16671 13047 16677
rect 14274 16668 14280 16680
rect 14332 16668 14338 16720
rect 15534 16711 15592 16717
rect 15534 16708 15546 16711
rect 14936 16680 15546 16708
rect 7466 16649 7472 16652
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16609 7251 16643
rect 7460 16640 7472 16649
rect 7379 16612 7472 16640
rect 7193 16603 7251 16609
rect 7460 16603 7472 16612
rect 7524 16640 7530 16652
rect 8202 16640 8208 16652
rect 7524 16612 8208 16640
rect 7466 16600 7472 16603
rect 7524 16600 7530 16612
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 9766 16640 9772 16652
rect 9692 16612 9772 16640
rect 5626 16572 5632 16584
rect 5368 16544 5632 16572
rect 5077 16535 5135 16541
rect 3142 16504 3148 16516
rect 2884 16476 3148 16504
rect 3142 16464 3148 16476
rect 3200 16464 3206 16516
rect 3418 16464 3424 16516
rect 3476 16504 3482 16516
rect 4890 16504 4896 16516
rect 3476 16476 4896 16504
rect 3476 16464 3482 16476
rect 4890 16464 4896 16476
rect 4948 16504 4954 16516
rect 5092 16504 5120 16535
rect 5626 16532 5632 16544
rect 5684 16532 5690 16584
rect 5902 16572 5908 16584
rect 5863 16544 5908 16572
rect 5902 16532 5908 16544
rect 5960 16532 5966 16584
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 6733 16575 6791 16581
rect 6733 16572 6745 16575
rect 6696 16544 6745 16572
rect 6696 16532 6702 16544
rect 6733 16541 6745 16544
rect 6779 16541 6791 16575
rect 9122 16572 9128 16584
rect 9083 16544 9128 16572
rect 6733 16535 6791 16541
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 9272 16544 9317 16572
rect 9272 16532 9278 16544
rect 4948 16476 5120 16504
rect 4948 16464 4954 16476
rect 5350 16436 5356 16448
rect 5311 16408 5356 16436
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 5920 16436 5948 16532
rect 8573 16507 8631 16513
rect 8573 16473 8585 16507
rect 8619 16504 8631 16507
rect 9232 16504 9260 16532
rect 9398 16504 9404 16516
rect 8619 16476 9404 16504
rect 8619 16473 8631 16476
rect 8573 16467 8631 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 9692 16513 9720 16612
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 11241 16643 11299 16649
rect 11241 16640 11253 16643
rect 10744 16612 11253 16640
rect 10744 16600 10750 16612
rect 11241 16609 11253 16612
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16640 11391 16643
rect 11790 16640 11796 16652
rect 11379 16612 11796 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 12161 16643 12219 16649
rect 12161 16609 12173 16643
rect 12207 16640 12219 16643
rect 12526 16640 12532 16652
rect 12207 16612 12532 16640
rect 12207 16609 12219 16612
rect 12161 16603 12219 16609
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 13814 16640 13820 16652
rect 13775 16612 13820 16640
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 14642 16640 14648 16652
rect 14603 16612 14648 16640
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 10134 16572 10140 16584
rect 10095 16544 10140 16572
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 11514 16572 11520 16584
rect 10367 16544 10548 16572
rect 11475 16544 11520 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 9677 16507 9735 16513
rect 9677 16473 9689 16507
rect 9723 16473 9735 16507
rect 9677 16467 9735 16473
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 10410 16504 10416 16516
rect 9824 16476 10416 16504
rect 9824 16464 9830 16476
rect 10410 16464 10416 16476
rect 10468 16464 10474 16516
rect 8110 16436 8116 16448
rect 5920 16408 8116 16436
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 10520 16436 10548 16544
rect 11514 16532 11520 16544
rect 11572 16572 11578 16584
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11572 16544 12265 16572
rect 11572 16532 11578 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16541 13231 16575
rect 13173 16535 13231 16541
rect 13188 16504 13216 16535
rect 13262 16532 13268 16584
rect 13320 16572 13326 16584
rect 13909 16575 13967 16581
rect 13909 16572 13921 16575
rect 13320 16544 13921 16572
rect 13320 16532 13326 16544
rect 13909 16541 13921 16544
rect 13955 16541 13967 16575
rect 13909 16535 13967 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14550 16572 14556 16584
rect 14139 16544 14556 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 14550 16532 14556 16544
rect 14608 16572 14614 16584
rect 14829 16575 14887 16581
rect 14829 16572 14841 16575
rect 14608 16544 14841 16572
rect 14608 16532 14614 16544
rect 14829 16541 14841 16544
rect 14875 16541 14887 16575
rect 14829 16535 14887 16541
rect 14936 16504 14964 16680
rect 15534 16677 15546 16680
rect 15580 16708 15592 16711
rect 16114 16708 16120 16720
rect 15580 16680 16120 16708
rect 15580 16677 15592 16680
rect 15534 16671 15592 16677
rect 16114 16668 16120 16680
rect 16172 16668 16178 16720
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15252 16612 15301 16640
rect 15252 16600 15258 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16640 16819 16643
rect 17218 16640 17224 16652
rect 16807 16612 17224 16640
rect 16807 16609 16819 16612
rect 16761 16603 16819 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 20257 16643 20315 16649
rect 20257 16640 20269 16643
rect 19576 16612 20269 16640
rect 19576 16600 19582 16612
rect 20257 16609 20269 16612
rect 20303 16609 20315 16643
rect 20257 16603 20315 16609
rect 20533 16643 20591 16649
rect 20533 16609 20545 16643
rect 20579 16640 20591 16643
rect 20806 16640 20812 16652
rect 20579 16612 20812 16640
rect 20579 16609 20591 16612
rect 20533 16603 20591 16609
rect 20806 16600 20812 16612
rect 20864 16600 20870 16652
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 20956 16612 21001 16640
rect 20956 16600 20962 16612
rect 16666 16504 16672 16516
rect 13188 16476 14964 16504
rect 16627 16476 16672 16504
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 8720 16408 10548 16436
rect 8720 16396 8726 16408
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 13630 16436 13636 16448
rect 10928 16408 13636 16436
rect 10928 16396 10934 16408
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14274 16436 14280 16448
rect 14235 16408 14280 16436
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 3694 16232 3700 16244
rect 3655 16204 3700 16232
rect 3694 16192 3700 16204
rect 3752 16192 3758 16244
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4433 16235 4491 16241
rect 4433 16232 4445 16235
rect 4304 16204 4445 16232
rect 4304 16192 4310 16204
rect 4433 16201 4445 16204
rect 4479 16201 4491 16235
rect 4433 16195 4491 16201
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 6362 16232 6368 16244
rect 5224 16204 6368 16232
rect 5224 16192 5230 16204
rect 6362 16192 6368 16204
rect 6420 16232 6426 16244
rect 8202 16232 8208 16244
rect 6420 16204 7788 16232
rect 8163 16204 8208 16232
rect 6420 16192 6426 16204
rect 1946 16164 1952 16176
rect 1907 16136 1952 16164
rect 1946 16124 1952 16136
rect 2004 16124 2010 16176
rect 7760 16164 7788 16204
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 10134 16232 10140 16244
rect 8895 16204 10140 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10888 16204 11928 16232
rect 10888 16164 10916 16204
rect 7760 16136 10916 16164
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 4985 16099 5043 16105
rect 4985 16096 4997 16099
rect 4948 16068 4997 16096
rect 4948 16056 4954 16068
rect 4985 16065 4997 16068
rect 5031 16065 5043 16099
rect 9398 16096 9404 16108
rect 9359 16068 9404 16096
rect 4985 16059 5043 16065
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10192 16068 10517 16096
rect 10192 16056 10198 16068
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10836 16068 10885 16096
rect 10836 16056 10842 16068
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 11900 16096 11928 16204
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 12253 16235 12311 16241
rect 12253 16232 12265 16235
rect 12032 16204 12265 16232
rect 12032 16192 12038 16204
rect 12253 16201 12265 16204
rect 12299 16201 12311 16235
rect 12253 16195 12311 16201
rect 13081 16235 13139 16241
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13262 16232 13268 16244
rect 13127 16204 13268 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 13872 16204 13921 16232
rect 13872 16192 13878 16204
rect 13909 16201 13921 16204
rect 13955 16201 13967 16235
rect 13909 16195 13967 16201
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 14737 16235 14795 16241
rect 14737 16232 14749 16235
rect 14700 16204 14749 16232
rect 14700 16192 14706 16204
rect 14737 16201 14749 16204
rect 14783 16201 14795 16235
rect 14737 16195 14795 16201
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18233 16235 18291 16241
rect 18233 16232 18245 16235
rect 18012 16204 18245 16232
rect 18012 16192 18018 16204
rect 18233 16201 18245 16204
rect 18279 16201 18291 16235
rect 20346 16232 20352 16244
rect 20307 16204 20352 16232
rect 18233 16195 18291 16201
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 13354 16124 13360 16176
rect 13412 16164 13418 16176
rect 14090 16164 14096 16176
rect 13412 16136 14096 16164
rect 13412 16124 13418 16136
rect 14090 16124 14096 16136
rect 14148 16124 14154 16176
rect 19518 16164 19524 16176
rect 15396 16136 19524 16164
rect 11900 16068 12572 16096
rect 10873 16059 10931 16065
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 2222 16028 2228 16040
rect 1811 16000 2228 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 15997 2375 16031
rect 2317 15991 2375 15997
rect 2584 16031 2642 16037
rect 2584 15997 2596 16031
rect 2630 16028 2642 16031
rect 3418 16028 3424 16040
rect 2630 16000 3424 16028
rect 2630 15997 2642 16000
rect 2584 15991 2642 15997
rect 2332 15960 2360 15991
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 4062 16028 4068 16040
rect 3896 16000 4068 16028
rect 3896 15972 3924 16000
rect 4062 15988 4068 16000
rect 4120 16028 4126 16040
rect 5261 16031 5319 16037
rect 5261 16028 5273 16031
rect 4120 16000 5273 16028
rect 4120 15988 4126 16000
rect 5261 15997 5273 16000
rect 5307 15997 5319 16031
rect 5261 15991 5319 15997
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7650 16028 7656 16040
rect 6871 16000 7656 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 8662 15988 8668 16040
rect 8720 16028 8726 16040
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 8720 16000 9229 16028
rect 8720 15988 8726 16000
rect 9217 15997 9229 16000
rect 9263 15997 9275 16031
rect 10888 16028 10916 16059
rect 12250 16028 12256 16040
rect 10888 16000 12256 16028
rect 9217 15991 9275 15997
rect 12250 15988 12256 16000
rect 12308 15988 12314 16040
rect 12544 16028 12572 16068
rect 12618 16056 12624 16108
rect 12676 16096 12682 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 12676 16068 13553 16096
rect 12676 16056 12682 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 14182 16096 14188 16108
rect 13771 16068 14188 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 14182 16056 14188 16068
rect 14240 16096 14246 16108
rect 14458 16096 14464 16108
rect 14240 16068 14464 16096
rect 14240 16056 14246 16068
rect 14458 16056 14464 16068
rect 14516 16096 14522 16108
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 14516 16068 15301 16096
rect 14516 16056 14522 16068
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15289 16059 15347 16065
rect 13998 16028 14004 16040
rect 12544 16000 14004 16028
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 15197 16031 15255 16037
rect 15197 16028 15209 16031
rect 14108 16000 15209 16028
rect 2406 15960 2412 15972
rect 2319 15932 2412 15960
rect 2406 15920 2412 15932
rect 2464 15960 2470 15972
rect 3878 15960 3884 15972
rect 2464 15932 3884 15960
rect 2464 15920 2470 15932
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 5534 15969 5540 15972
rect 4341 15963 4399 15969
rect 4341 15929 4353 15963
rect 4387 15960 4399 15963
rect 5528 15960 5540 15969
rect 4387 15932 4936 15960
rect 5495 15932 5540 15960
rect 4387 15929 4399 15932
rect 4341 15923 4399 15929
rect 4908 15904 4936 15932
rect 5528 15923 5540 15932
rect 5534 15920 5540 15923
rect 5592 15920 5598 15972
rect 11146 15969 11152 15972
rect 7070 15963 7128 15969
rect 7070 15960 7082 15963
rect 6840 15932 7082 15960
rect 2682 15852 2688 15904
rect 2740 15892 2746 15904
rect 3510 15892 3516 15904
rect 2740 15864 3516 15892
rect 2740 15852 2746 15864
rect 3510 15852 3516 15864
rect 3568 15892 3574 15904
rect 4801 15895 4859 15901
rect 4801 15892 4813 15895
rect 3568 15864 4813 15892
rect 3568 15852 3574 15864
rect 4801 15861 4813 15864
rect 4847 15861 4859 15895
rect 4801 15855 4859 15861
rect 4890 15852 4896 15904
rect 4948 15892 4954 15904
rect 6638 15892 6644 15904
rect 4948 15864 4993 15892
rect 6599 15864 6644 15892
rect 4948 15852 4954 15864
rect 6638 15852 6644 15864
rect 6696 15892 6702 15904
rect 6840 15892 6868 15932
rect 7070 15929 7082 15932
rect 7116 15929 7128 15963
rect 9309 15963 9367 15969
rect 9309 15960 9321 15963
rect 7070 15923 7128 15929
rect 8680 15932 9321 15960
rect 6696 15864 6868 15892
rect 6696 15852 6702 15864
rect 8570 15852 8576 15904
rect 8628 15892 8634 15904
rect 8680 15901 8708 15932
rect 9309 15929 9321 15932
rect 9355 15929 9367 15963
rect 9309 15923 9367 15929
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 11140 15960 11152 15969
rect 10367 15932 11008 15960
rect 11107 15932 11152 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8628 15864 8677 15892
rect 8628 15852 8634 15864
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 9950 15892 9956 15904
rect 9911 15864 9956 15892
rect 8665 15855 8723 15861
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10980 15892 11008 15932
rect 11140 15923 11152 15932
rect 11146 15920 11152 15923
rect 11204 15920 11210 15972
rect 14108 15960 14136 16000
rect 15197 15997 15209 16000
rect 15243 16028 15255 16031
rect 15396 16028 15424 16136
rect 19518 16124 19524 16136
rect 19576 16124 19582 16176
rect 16482 16056 16488 16108
rect 16540 16096 16546 16108
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16540 16068 16957 16096
rect 16540 16056 16546 16068
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17126 16056 17132 16108
rect 17184 16096 17190 16108
rect 19797 16099 19855 16105
rect 17184 16068 19564 16096
rect 17184 16056 17190 16068
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 15243 16000 15424 16028
rect 16224 16000 18061 16028
rect 15243 15997 15255 16000
rect 15197 15991 15255 15997
rect 14274 15960 14280 15972
rect 12544 15932 14136 15960
rect 14187 15932 14280 15960
rect 12544 15904 12572 15932
rect 14274 15920 14280 15932
rect 14332 15960 14338 15972
rect 16224 15960 16252 16000
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 19426 16028 19432 16040
rect 18095 16000 19432 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 19426 15988 19432 16000
rect 19484 15988 19490 16040
rect 19536 16037 19564 16068
rect 19797 16065 19809 16099
rect 19843 16096 19855 16099
rect 20622 16096 20628 16108
rect 19843 16068 20628 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 19521 16031 19579 16037
rect 19521 15997 19533 16031
rect 19567 15997 19579 16031
rect 20162 16028 20168 16040
rect 20123 16000 20168 16028
rect 19521 15991 19579 15997
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20898 16028 20904 16040
rect 20859 16000 20904 16028
rect 20533 15991 20591 15997
rect 14332 15932 16252 15960
rect 16761 15963 16819 15969
rect 14332 15920 14338 15932
rect 16761 15929 16773 15963
rect 16807 15960 16819 15963
rect 18598 15960 18604 15972
rect 16807 15932 18604 15960
rect 16807 15929 16819 15932
rect 16761 15923 16819 15929
rect 18598 15920 18604 15932
rect 18656 15920 18662 15972
rect 19334 15920 19340 15972
rect 19392 15960 19398 15972
rect 20548 15960 20576 15991
rect 20898 15988 20904 16000
rect 20956 15988 20962 16040
rect 19392 15932 20576 15960
rect 19392 15920 19398 15932
rect 11054 15892 11060 15904
rect 10468 15864 10513 15892
rect 10980 15864 11060 15892
rect 10468 15852 10474 15864
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 12526 15852 12532 15904
rect 12584 15852 12590 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 13412 15864 13461 15892
rect 13412 15852 13418 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 14366 15852 14372 15904
rect 14424 15892 14430 15904
rect 15102 15892 15108 15904
rect 14424 15864 14469 15892
rect 15063 15864 15108 15892
rect 14424 15852 14430 15864
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 16390 15892 16396 15904
rect 16351 15864 16396 15892
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17221 15895 17279 15901
rect 16908 15864 16953 15892
rect 16908 15852 16914 15864
rect 17221 15861 17233 15895
rect 17267 15892 17279 15895
rect 17954 15892 17960 15904
rect 17267 15864 17960 15892
rect 17267 15861 17279 15864
rect 17221 15855 17279 15861
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 20680 15864 21097 15892
rect 20680 15852 20686 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21085 15855 21143 15861
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 2041 15691 2099 15697
rect 2041 15657 2053 15691
rect 2087 15688 2099 15691
rect 2774 15688 2780 15700
rect 2087 15660 2780 15688
rect 2087 15657 2099 15660
rect 2041 15651 2099 15657
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 3050 15688 3056 15700
rect 2915 15660 3056 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 3329 15691 3387 15697
rect 3329 15657 3341 15691
rect 3375 15688 3387 15691
rect 5166 15688 5172 15700
rect 3375 15660 5172 15688
rect 3375 15657 3387 15660
rect 3329 15651 3387 15657
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 6825 15691 6883 15697
rect 6825 15688 6837 15691
rect 6604 15660 6837 15688
rect 6604 15648 6610 15660
rect 6825 15657 6837 15660
rect 6871 15657 6883 15691
rect 6825 15651 6883 15657
rect 8757 15691 8815 15697
rect 8757 15657 8769 15691
rect 8803 15688 8815 15691
rect 8846 15688 8852 15700
rect 8803 15660 8852 15688
rect 8803 15657 8815 15660
rect 8757 15651 8815 15657
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 9125 15691 9183 15697
rect 9125 15657 9137 15691
rect 9171 15688 9183 15691
rect 9950 15688 9956 15700
rect 9171 15660 9956 15688
rect 9171 15657 9183 15660
rect 9125 15651 9183 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 12066 15688 12072 15700
rect 12027 15660 12072 15688
rect 12066 15648 12072 15660
rect 12124 15648 12130 15700
rect 12437 15691 12495 15697
rect 12437 15657 12449 15691
rect 12483 15688 12495 15691
rect 12802 15688 12808 15700
rect 12483 15660 12808 15688
rect 12483 15657 12495 15660
rect 12437 15651 12495 15657
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13354 15688 13360 15700
rect 13315 15660 13360 15688
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 13630 15648 13636 15700
rect 13688 15688 13694 15700
rect 13725 15691 13783 15697
rect 13725 15688 13737 15691
rect 13688 15660 13737 15688
rect 13688 15648 13694 15660
rect 13725 15657 13737 15660
rect 13771 15657 13783 15691
rect 13725 15651 13783 15657
rect 14185 15691 14243 15697
rect 14185 15657 14197 15691
rect 14231 15688 14243 15691
rect 14366 15688 14372 15700
rect 14231 15660 14372 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 15160 15660 15301 15688
rect 15160 15648 15166 15660
rect 15289 15657 15301 15660
rect 15335 15657 15347 15691
rect 15289 15651 15347 15657
rect 16390 15648 16396 15700
rect 16448 15688 16454 15700
rect 18049 15691 18107 15697
rect 18049 15688 18061 15691
rect 16448 15660 18061 15688
rect 16448 15648 16454 15660
rect 18049 15657 18061 15660
rect 18095 15657 18107 15691
rect 18049 15651 18107 15657
rect 18141 15691 18199 15697
rect 18141 15657 18153 15691
rect 18187 15688 18199 15691
rect 18506 15688 18512 15700
rect 18187 15660 18512 15688
rect 18187 15657 18199 15660
rect 18141 15651 18199 15657
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 20254 15688 20260 15700
rect 20215 15660 20260 15688
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 1762 15620 1768 15632
rect 1723 15592 1768 15620
rect 1762 15580 1768 15592
rect 1820 15580 1826 15632
rect 2409 15623 2467 15629
rect 2409 15589 2421 15623
rect 2455 15620 2467 15623
rect 3697 15623 3755 15629
rect 3697 15620 3709 15623
rect 2455 15592 3709 15620
rect 2455 15589 2467 15592
rect 2409 15583 2467 15589
rect 3697 15589 3709 15592
rect 3743 15589 3755 15623
rect 3697 15583 3755 15589
rect 6365 15623 6423 15629
rect 6365 15589 6377 15623
rect 6411 15620 6423 15623
rect 8018 15620 8024 15632
rect 6411 15592 8024 15620
rect 6411 15589 6423 15592
rect 6365 15583 6423 15589
rect 8018 15580 8024 15592
rect 8076 15580 8082 15632
rect 11974 15580 11980 15632
rect 12032 15620 12038 15632
rect 12032 15592 12664 15620
rect 12032 15580 12038 15592
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 2130 15552 2136 15564
rect 1535 15524 2136 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 2130 15512 2136 15524
rect 2188 15512 2194 15564
rect 3237 15555 3295 15561
rect 3237 15552 3249 15555
rect 2240 15524 3249 15552
rect 1302 15444 1308 15496
rect 1360 15484 1366 15496
rect 2240 15484 2268 15524
rect 3237 15521 3249 15524
rect 3283 15521 3295 15555
rect 3237 15515 3295 15521
rect 4700 15555 4758 15561
rect 4700 15521 4712 15555
rect 4746 15552 4758 15555
rect 6546 15552 6552 15564
rect 4746 15524 6552 15552
rect 4746 15521 4758 15524
rect 4700 15515 4758 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 7190 15552 7196 15564
rect 7151 15524 7196 15552
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 9122 15552 9128 15564
rect 7331 15524 9128 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 9217 15555 9275 15561
rect 9217 15521 9229 15555
rect 9263 15552 9275 15555
rect 9950 15552 9956 15564
rect 9263 15524 9956 15552
rect 9263 15521 9275 15524
rect 9217 15515 9275 15521
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 10134 15561 10140 15564
rect 10128 15552 10140 15561
rect 10095 15524 10140 15552
rect 10128 15515 10140 15524
rect 10134 15512 10140 15515
rect 10192 15512 10198 15564
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12434 15552 12440 15564
rect 12216 15524 12440 15552
rect 12216 15512 12222 15524
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 1360 15456 2268 15484
rect 1360 15444 1366 15456
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2464 15456 2513 15484
rect 2464 15444 2470 15456
rect 2501 15453 2513 15456
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 3418 15484 3424 15496
rect 2731 15456 3424 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 3878 15444 3884 15496
rect 3936 15484 3942 15496
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 3936 15456 4445 15484
rect 3936 15444 3942 15456
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 4433 15447 4491 15453
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6638 15484 6644 15496
rect 6599 15456 6644 15484
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 7466 15484 7472 15496
rect 7427 15456 7472 15484
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15484 7711 15487
rect 8386 15484 8392 15496
rect 7699 15456 8392 15484
rect 7699 15453 7711 15456
rect 7653 15447 7711 15453
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 5997 15419 6055 15425
rect 5997 15385 6009 15419
rect 6043 15416 6055 15419
rect 6914 15416 6920 15428
rect 6043 15388 6920 15416
rect 6043 15385 6055 15388
rect 5997 15379 6055 15385
rect 6914 15376 6920 15388
rect 6972 15376 6978 15428
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 5813 15351 5871 15357
rect 5813 15348 5825 15351
rect 5592 15320 5825 15348
rect 5592 15308 5598 15320
rect 5813 15317 5825 15320
rect 5859 15348 5871 15351
rect 7466 15348 7472 15360
rect 5859 15320 7472 15348
rect 5859 15317 5871 15320
rect 5813 15311 5871 15317
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 9416 15348 9444 15447
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 9861 15487 9919 15493
rect 9861 15484 9873 15487
rect 9640 15456 9873 15484
rect 9640 15444 9646 15456
rect 9861 15453 9873 15456
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 12066 15444 12072 15496
rect 12124 15484 12130 15496
rect 12636 15493 12664 15592
rect 12894 15580 12900 15632
rect 12952 15620 12958 15632
rect 12952 15592 13952 15620
rect 12952 15580 12958 15592
rect 13924 15552 13952 15592
rect 13998 15580 14004 15632
rect 14056 15620 14062 15632
rect 19150 15620 19156 15632
rect 14056 15592 19156 15620
rect 14056 15580 14062 15592
rect 19150 15580 19156 15592
rect 19208 15620 19214 15632
rect 19208 15592 20944 15620
rect 19208 15580 19214 15592
rect 14550 15552 14556 15564
rect 13924 15524 14556 15552
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 16482 15561 16488 15564
rect 16476 15552 16488 15561
rect 16443 15524 16488 15552
rect 16476 15515 16488 15524
rect 16482 15512 16488 15515
rect 16540 15512 16546 15564
rect 18509 15555 18567 15561
rect 18509 15521 18521 15555
rect 18555 15552 18567 15555
rect 18966 15552 18972 15564
rect 18555 15524 18972 15552
rect 18555 15521 18567 15524
rect 18509 15515 18567 15521
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 20070 15552 20076 15564
rect 20031 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 20916 15561 20944 15592
rect 20441 15555 20499 15561
rect 20441 15521 20453 15555
rect 20487 15521 20499 15555
rect 20441 15515 20499 15521
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 12124 15456 12541 15484
rect 12124 15444 12130 15456
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15453 12679 15487
rect 13630 15484 13636 15496
rect 12621 15447 12679 15453
rect 12811 15456 13636 15484
rect 10870 15376 10876 15428
rect 10928 15416 10934 15428
rect 12811 15416 12839 15456
rect 13630 15444 13636 15456
rect 13688 15484 13694 15496
rect 13817 15487 13875 15493
rect 13817 15484 13829 15487
rect 13688 15456 13829 15484
rect 13688 15444 13694 15456
rect 13817 15453 13829 15456
rect 13863 15453 13875 15487
rect 13817 15447 13875 15453
rect 14001 15487 14059 15493
rect 14001 15453 14013 15487
rect 14047 15453 14059 15487
rect 14001 15447 14059 15453
rect 10928 15388 12839 15416
rect 10928 15376 10934 15388
rect 13722 15376 13728 15428
rect 13780 15416 13786 15428
rect 14016 15416 14044 15447
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14516 15456 14657 15484
rect 14516 15444 14522 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14752 15416 14780 15447
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 15252 15456 16221 15484
rect 15252 15444 15258 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15453 18291 15487
rect 18782 15484 18788 15496
rect 18743 15456 18788 15484
rect 18233 15447 18291 15453
rect 17586 15416 17592 15428
rect 13780 15388 14780 15416
rect 17499 15388 17592 15416
rect 13780 15376 13786 15388
rect 17586 15376 17592 15388
rect 17644 15416 17650 15428
rect 18248 15416 18276 15447
rect 18782 15444 18788 15456
rect 18840 15444 18846 15496
rect 19886 15444 19892 15496
rect 19944 15484 19950 15496
rect 20456 15484 20484 15515
rect 19944 15456 20484 15484
rect 19944 15444 19950 15456
rect 17644 15388 18276 15416
rect 17644 15376 17650 15388
rect 11146 15348 11152 15360
rect 9416 15320 11152 15348
rect 11146 15308 11152 15320
rect 11204 15348 11210 15360
rect 11241 15351 11299 15357
rect 11241 15348 11253 15351
rect 11204 15320 11253 15348
rect 11204 15308 11210 15320
rect 11241 15317 11253 15320
rect 11287 15317 11299 15351
rect 11241 15311 11299 15317
rect 17681 15351 17739 15357
rect 17681 15317 17693 15351
rect 17727 15348 17739 15351
rect 19242 15348 19248 15360
rect 17727 15320 19248 15348
rect 17727 15317 17739 15320
rect 17681 15311 17739 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 20438 15308 20444 15360
rect 20496 15348 20502 15360
rect 20625 15351 20683 15357
rect 20625 15348 20637 15351
rect 20496 15320 20637 15348
rect 20496 15308 20502 15320
rect 20625 15317 20637 15320
rect 20671 15317 20683 15351
rect 21082 15348 21088 15360
rect 21043 15320 21088 15348
rect 20625 15311 20683 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 1578 15144 1584 15156
rect 1539 15116 1584 15144
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 2685 15147 2743 15153
rect 2685 15113 2697 15147
rect 2731 15144 2743 15147
rect 2774 15144 2780 15156
rect 2731 15116 2780 15144
rect 2731 15113 2743 15116
rect 2685 15107 2743 15113
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 3053 15147 3111 15153
rect 3053 15144 3065 15147
rect 2924 15116 3065 15144
rect 2924 15104 2930 15116
rect 3053 15113 3065 15116
rect 3099 15113 3111 15147
rect 7190 15144 7196 15156
rect 7151 15116 7196 15144
rect 3053 15107 3111 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 8018 15144 8024 15156
rect 7979 15116 8024 15144
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 10008 15116 11529 15144
rect 10008 15104 10014 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 12636 15116 15148 15144
rect 3786 15076 3792 15088
rect 2148 15048 3792 15076
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 2038 14940 2044 14952
rect 1811 14912 2044 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 1412 14872 1440 14903
rect 2038 14900 2044 14912
rect 2096 14900 2102 14952
rect 2148 14949 2176 15048
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 6178 15076 6184 15088
rect 3896 15048 6184 15076
rect 3896 15008 3924 15048
rect 6178 15036 6184 15048
rect 6236 15036 6242 15088
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 10229 15079 10287 15085
rect 7524 15048 8616 15076
rect 7524 15036 7530 15048
rect 4062 15008 4068 15020
rect 2240 14980 3924 15008
rect 4023 14980 4068 15008
rect 2133 14943 2191 14949
rect 2133 14909 2145 14943
rect 2179 14909 2191 14943
rect 2133 14903 2191 14909
rect 2240 14872 2268 14980
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4798 15008 4804 15020
rect 4759 14980 4804 15008
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 5902 15008 5908 15020
rect 5863 14980 5908 15008
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 6696 14980 7757 15008
rect 6696 14968 6702 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 8478 15008 8484 15020
rect 8439 14980 8484 15008
rect 7745 14971 7803 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8588 15017 8616 15048
rect 10229 15045 10241 15079
rect 10275 15045 10287 15079
rect 10229 15039 10287 15045
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 14977 8631 15011
rect 8846 15008 8852 15020
rect 8807 14980 8852 15008
rect 8573 14971 8631 14977
rect 8846 14968 8852 14980
rect 8904 14968 8910 15020
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10244 15008 10272 15039
rect 10686 15036 10692 15088
rect 10744 15076 10750 15088
rect 12636 15076 12664 15116
rect 10744 15048 12664 15076
rect 12713 15079 12771 15085
rect 10744 15036 10750 15048
rect 12713 15045 12725 15079
rect 12759 15076 12771 15079
rect 15010 15076 15016 15088
rect 12759 15048 15016 15076
rect 12759 15045 12771 15048
rect 12713 15039 12771 15045
rect 15010 15036 15016 15048
rect 15068 15036 15074 15088
rect 11333 15011 11391 15017
rect 10192 14980 11008 15008
rect 10192 14968 10198 14980
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14909 2559 14943
rect 2866 14940 2872 14952
rect 2827 14912 2872 14940
rect 2501 14903 2559 14909
rect 1412 14844 2268 14872
rect 2516 14872 2544 14903
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 4540 14912 5396 14940
rect 4540 14872 4568 14912
rect 2516 14844 4568 14872
rect 4617 14875 4675 14881
rect 4617 14841 4629 14875
rect 4663 14872 4675 14875
rect 4890 14872 4896 14884
rect 4663 14844 4896 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 4890 14832 4896 14844
rect 4948 14832 4954 14884
rect 5368 14872 5396 14912
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7340 14912 7573 14940
rect 7340 14900 7346 14912
rect 7561 14909 7573 14912
rect 7607 14909 7619 14943
rect 7561 14903 7619 14909
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7926 14940 7932 14952
rect 7699 14912 7932 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8386 14940 8392 14952
rect 8347 14912 8392 14940
rect 8386 14900 8392 14912
rect 8444 14900 8450 14952
rect 10870 14940 10876 14952
rect 8772 14912 10876 14940
rect 8772 14872 8800 14912
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 10980 14940 11008 14980
rect 11333 14977 11345 15011
rect 11379 15008 11391 15011
rect 11422 15008 11428 15020
rect 11379 14980 11428 15008
rect 11379 14977 11391 14980
rect 11333 14971 11391 14977
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15008 13415 15011
rect 13906 15008 13912 15020
rect 13403 14980 13912 15008
rect 13403 14977 13415 14980
rect 13357 14971 13415 14977
rect 12084 14940 12112 14971
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 14182 15008 14188 15020
rect 14143 14980 14188 15008
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 10980 14912 12112 14940
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 13688 14912 14688 14940
rect 13688 14900 13694 14912
rect 5368 14844 8800 14872
rect 9116 14875 9174 14881
rect 9116 14841 9128 14875
rect 9162 14872 9174 14875
rect 9306 14872 9312 14884
rect 9162 14844 9312 14872
rect 9162 14841 9174 14844
rect 9116 14835 9174 14841
rect 9306 14832 9312 14844
rect 9364 14832 9370 14884
rect 13081 14875 13139 14881
rect 13081 14841 13093 14875
rect 13127 14872 13139 14875
rect 14274 14872 14280 14884
rect 13127 14844 14280 14872
rect 13127 14841 13139 14844
rect 13081 14835 13139 14841
rect 14274 14832 14280 14844
rect 14332 14832 14338 14884
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2314 14804 2320 14816
rect 2275 14776 2320 14804
rect 2314 14764 2320 14776
rect 2372 14764 2378 14816
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3421 14807 3479 14813
rect 3421 14804 3433 14807
rect 3016 14776 3433 14804
rect 3016 14764 3022 14776
rect 3421 14773 3433 14776
rect 3467 14773 3479 14807
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 3421 14767 3479 14773
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 3881 14807 3939 14813
rect 3881 14773 3893 14807
rect 3927 14804 3939 14807
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 3927 14776 4261 14804
rect 3927 14773 3939 14776
rect 3881 14767 3939 14773
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 4249 14767 4307 14773
rect 4709 14807 4767 14813
rect 4709 14773 4721 14807
rect 4755 14804 4767 14807
rect 5353 14807 5411 14813
rect 5353 14804 5365 14807
rect 4755 14776 5365 14804
rect 4755 14773 4767 14776
rect 4709 14767 4767 14773
rect 5353 14773 5365 14776
rect 5399 14773 5411 14807
rect 5718 14804 5724 14816
rect 5679 14776 5724 14804
rect 5353 14767 5411 14773
rect 5718 14764 5724 14776
rect 5776 14764 5782 14816
rect 5813 14807 5871 14813
rect 5813 14773 5825 14807
rect 5859 14804 5871 14807
rect 5994 14804 6000 14816
rect 5859 14776 6000 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6270 14764 6276 14816
rect 6328 14804 6334 14816
rect 8478 14804 8484 14816
rect 6328 14776 8484 14804
rect 6328 14764 6334 14776
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 10778 14804 10784 14816
rect 10735 14776 10784 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11057 14807 11115 14813
rect 11057 14804 11069 14807
rect 11020 14776 11069 14804
rect 11020 14764 11026 14776
rect 11057 14773 11069 14776
rect 11103 14773 11115 14807
rect 11057 14767 11115 14773
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11882 14804 11888 14816
rect 11204 14776 11249 14804
rect 11843 14776 11888 14804
rect 11204 14764 11210 14776
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 13170 14804 13176 14816
rect 12032 14776 12077 14804
rect 13131 14776 13176 14804
rect 12032 14764 12038 14776
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13541 14807 13599 14813
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 13722 14804 13728 14816
rect 13587 14776 13728 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 13909 14807 13967 14813
rect 13909 14804 13921 14807
rect 13872 14776 13921 14804
rect 13872 14764 13878 14776
rect 13909 14773 13921 14776
rect 13955 14773 13967 14807
rect 13909 14767 13967 14773
rect 14001 14807 14059 14813
rect 14001 14773 14013 14807
rect 14047 14804 14059 14807
rect 14550 14804 14556 14816
rect 14047 14776 14556 14804
rect 14047 14773 14059 14776
rect 14001 14767 14059 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 14660 14804 14688 14912
rect 15120 14872 15148 15116
rect 16850 15104 16856 15156
rect 16908 15144 16914 15156
rect 17037 15147 17095 15153
rect 17037 15144 17049 15147
rect 16908 15116 17049 15144
rect 16908 15104 16914 15116
rect 17037 15113 17049 15116
rect 17083 15113 17095 15147
rect 17037 15107 17095 15113
rect 18049 15147 18107 15153
rect 18049 15113 18061 15147
rect 18095 15144 18107 15147
rect 18598 15144 18604 15156
rect 18095 15116 18604 15144
rect 18095 15113 18107 15116
rect 18049 15107 18107 15113
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 19702 15144 19708 15156
rect 19659 15116 19708 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 19702 15104 19708 15116
rect 19760 15104 19766 15156
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 16724 15048 18736 15076
rect 16724 15036 16730 15048
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15565 15011 15623 15017
rect 15565 15008 15577 15011
rect 15252 14980 15577 15008
rect 15252 14968 15258 14980
rect 15565 14977 15577 14980
rect 15611 14977 15623 15011
rect 17681 15011 17739 15017
rect 17681 15008 17693 15011
rect 15565 14971 15623 14977
rect 16592 14980 17693 15008
rect 15832 14943 15890 14949
rect 15832 14909 15844 14943
rect 15878 14940 15890 14943
rect 16390 14940 16396 14952
rect 15878 14912 16396 14940
rect 15878 14909 15890 14912
rect 15832 14903 15890 14909
rect 16390 14900 16396 14912
rect 16448 14940 16454 14952
rect 16592 14940 16620 14980
rect 17681 14977 17693 14980
rect 17727 15008 17739 15011
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 17727 14980 18613 15008
rect 17727 14977 17739 14980
rect 17681 14971 17739 14977
rect 18601 14977 18613 14980
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 17494 14940 17500 14952
rect 16448 14912 16620 14940
rect 17455 14912 17500 14940
rect 16448 14900 16454 14912
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 18012 14912 18429 14940
rect 18012 14900 18018 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18708 14940 18736 15048
rect 18874 15036 18880 15088
rect 18932 15076 18938 15088
rect 18932 15048 20484 15076
rect 18932 15036 18938 15048
rect 18782 14968 18788 15020
rect 18840 15008 18846 15020
rect 20456 15008 20484 15048
rect 20530 15036 20536 15088
rect 20588 15076 20594 15088
rect 21085 15079 21143 15085
rect 21085 15076 21097 15079
rect 20588 15048 21097 15076
rect 20588 15036 20594 15048
rect 21085 15045 21097 15048
rect 21131 15045 21143 15079
rect 21085 15039 21143 15045
rect 18840 14980 20208 15008
rect 20456 14980 20944 15008
rect 18840 14968 18846 14980
rect 20180 14949 20208 14980
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 18708 14912 19441 14940
rect 18417 14903 18475 14909
rect 19429 14909 19441 14912
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14940 20591 14943
rect 20714 14940 20720 14952
rect 20579 14912 20720 14940
rect 20579 14909 20591 14912
rect 20533 14903 20591 14909
rect 17405 14875 17463 14881
rect 17405 14872 17417 14875
rect 15120 14844 17417 14872
rect 17405 14841 17417 14844
rect 17451 14872 17463 14875
rect 19812 14872 19840 14903
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 20916 14949 20944 14980
rect 20901 14943 20959 14949
rect 20901 14909 20913 14943
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 17451 14844 19840 14872
rect 17451 14841 17463 14844
rect 17405 14835 17463 14841
rect 20254 14832 20260 14884
rect 20312 14872 20318 14884
rect 20312 14844 20760 14872
rect 20312 14832 20318 14844
rect 15930 14804 15936 14816
rect 14660 14776 15936 14804
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 16022 14764 16028 14816
rect 16080 14804 16086 14816
rect 16482 14804 16488 14816
rect 16080 14776 16488 14804
rect 16080 14764 16086 14776
rect 16482 14764 16488 14776
rect 16540 14804 16546 14816
rect 16945 14807 17003 14813
rect 16945 14804 16957 14807
rect 16540 14776 16957 14804
rect 16540 14764 16546 14776
rect 16945 14773 16957 14776
rect 16991 14773 17003 14807
rect 16945 14767 17003 14773
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 18509 14807 18567 14813
rect 18509 14804 18521 14807
rect 18472 14776 18521 14804
rect 18472 14764 18478 14776
rect 18509 14773 18521 14776
rect 18555 14804 18567 14807
rect 18690 14804 18696 14816
rect 18555 14776 18696 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 19702 14764 19708 14816
rect 19760 14804 19766 14816
rect 19981 14807 20039 14813
rect 19981 14804 19993 14807
rect 19760 14776 19993 14804
rect 19760 14764 19766 14776
rect 19981 14773 19993 14776
rect 20027 14773 20039 14807
rect 20346 14804 20352 14816
rect 20307 14776 20352 14804
rect 19981 14767 20039 14773
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 20732 14813 20760 14844
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14773 20775 14807
rect 20717 14767 20775 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 3786 14600 3792 14612
rect 3191 14572 3792 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 4120 14572 5457 14600
rect 4120 14560 4126 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5994 14600 6000 14612
rect 5955 14572 6000 14600
rect 5445 14563 5503 14569
rect 2225 14535 2283 14541
rect 2225 14501 2237 14535
rect 2271 14532 2283 14535
rect 2866 14532 2872 14544
rect 2271 14504 2872 14532
rect 2271 14501 2283 14504
rect 2225 14495 2283 14501
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 4332 14535 4390 14541
rect 4332 14532 4344 14535
rect 3896 14504 4344 14532
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14433 1639 14467
rect 1581 14427 1639 14433
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2501 14467 2559 14473
rect 1995 14436 2360 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 1596 14328 1624 14427
rect 2332 14396 2360 14436
rect 2501 14433 2513 14467
rect 2547 14464 2559 14467
rect 3050 14464 3056 14476
rect 2547 14436 3056 14464
rect 2547 14433 2559 14436
rect 2501 14427 2559 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3510 14464 3516 14476
rect 3471 14436 3516 14464
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 3234 14396 3240 14408
rect 2332 14368 3240 14396
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3602 14396 3608 14408
rect 3563 14368 3608 14396
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 3789 14399 3847 14405
rect 3789 14365 3801 14399
rect 3835 14396 3847 14399
rect 3896 14396 3924 14504
rect 4332 14501 4344 14504
rect 4378 14532 4390 14535
rect 4798 14532 4804 14544
rect 4378 14504 4804 14532
rect 4378 14501 4390 14504
rect 4332 14495 4390 14501
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 5460 14532 5488 14563
rect 5994 14560 6000 14572
rect 6052 14560 6058 14612
rect 6454 14560 6460 14612
rect 6512 14600 6518 14612
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6512 14572 6837 14600
rect 6512 14560 6518 14572
rect 6825 14569 6837 14572
rect 6871 14569 6883 14603
rect 6825 14563 6883 14569
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7650 14600 7656 14612
rect 7248 14572 7656 14600
rect 7248 14560 7254 14572
rect 7650 14560 7656 14572
rect 7708 14600 7714 14612
rect 8846 14600 8852 14612
rect 7708 14572 8852 14600
rect 7708 14560 7714 14572
rect 6365 14535 6423 14541
rect 5460 14504 6316 14532
rect 6288 14464 6316 14504
rect 6365 14501 6377 14535
rect 6411 14532 6423 14535
rect 6730 14532 6736 14544
rect 6411 14504 6736 14532
rect 6411 14501 6423 14504
rect 6365 14495 6423 14501
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 7098 14464 7104 14476
rect 3835 14368 3924 14396
rect 3988 14436 6132 14464
rect 6288 14436 7104 14464
rect 3835 14365 3847 14368
rect 3789 14359 3847 14365
rect 3988 14328 4016 14436
rect 6104 14408 6132 14436
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 7193 14467 7251 14473
rect 7193 14433 7205 14467
rect 7239 14464 7251 14467
rect 7239 14436 7604 14464
rect 7239 14433 7251 14436
rect 7193 14427 7251 14433
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4120 14368 4165 14396
rect 4120 14356 4126 14368
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6328 14368 6469 14396
rect 6328 14356 6334 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 7282 14396 7288 14408
rect 6604 14368 6649 14396
rect 7243 14368 7288 14396
rect 6604 14356 6610 14368
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7466 14396 7472 14408
rect 7427 14368 7472 14396
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 1596 14300 4016 14328
rect 7576 14328 7604 14436
rect 7650 14424 7656 14476
rect 7708 14464 7714 14476
rect 7837 14467 7895 14473
rect 7837 14464 7849 14467
rect 7708 14436 7849 14464
rect 7708 14424 7714 14436
rect 7837 14433 7849 14436
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 7936 14467 7994 14473
rect 7936 14433 7948 14467
rect 7982 14464 7994 14467
rect 8027 14464 8055 14572
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10321 14603 10379 14609
rect 10321 14569 10333 14603
rect 10367 14600 10379 14603
rect 10781 14603 10839 14609
rect 10781 14600 10793 14603
rect 10367 14572 10793 14600
rect 10367 14569 10379 14572
rect 10321 14563 10379 14569
rect 10781 14569 10793 14572
rect 10827 14569 10839 14603
rect 10781 14563 10839 14569
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 11112 14572 11621 14600
rect 11112 14560 11118 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 13906 14600 13912 14612
rect 13867 14572 13912 14600
rect 11609 14563 11667 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 14182 14600 14188 14612
rect 14056 14572 14188 14600
rect 14056 14560 14062 14572
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 14829 14603 14887 14609
rect 14829 14569 14841 14603
rect 14875 14600 14887 14603
rect 15749 14603 15807 14609
rect 15749 14600 15761 14603
rect 14875 14572 15761 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 15749 14569 15761 14572
rect 15795 14569 15807 14603
rect 15749 14563 15807 14569
rect 15930 14560 15936 14612
rect 15988 14600 15994 14612
rect 16482 14600 16488 14612
rect 15988 14572 16488 14600
rect 15988 14560 15994 14572
rect 16482 14560 16488 14572
rect 16540 14600 16546 14612
rect 16540 14572 20944 14600
rect 16540 14560 16546 14572
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 13630 14532 13636 14544
rect 8168 14504 13636 14532
rect 8168 14492 8174 14504
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 17488 14535 17546 14541
rect 17488 14501 17500 14535
rect 17534 14532 17546 14535
rect 17586 14532 17592 14544
rect 17534 14504 17592 14532
rect 17534 14501 17546 14504
rect 17488 14495 17546 14501
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 17678 14492 17684 14544
rect 17736 14532 17742 14544
rect 19334 14532 19340 14544
rect 17736 14504 19340 14532
rect 17736 14492 17742 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 19886 14532 19892 14544
rect 19847 14504 19892 14532
rect 19886 14492 19892 14504
rect 19944 14492 19950 14544
rect 20070 14492 20076 14544
rect 20128 14532 20134 14544
rect 20441 14535 20499 14541
rect 20441 14532 20453 14535
rect 20128 14504 20453 14532
rect 20128 14492 20134 14504
rect 20441 14501 20453 14504
rect 20487 14501 20499 14535
rect 20441 14495 20499 14501
rect 8202 14473 8208 14476
rect 8196 14464 8208 14473
rect 7982 14436 8055 14464
rect 8163 14436 8208 14464
rect 7982 14433 7994 14436
rect 7936 14427 7994 14433
rect 8196 14427 8208 14436
rect 8260 14464 8266 14476
rect 11149 14467 11207 14473
rect 8260 14436 11008 14464
rect 8202 14424 8208 14427
rect 8260 14424 8266 14436
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 9456 14368 10425 14396
rect 9456 14356 9462 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 10643 14368 10732 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 7926 14328 7932 14340
rect 7576 14300 7932 14328
rect 7926 14288 7932 14300
rect 7984 14288 7990 14340
rect 9306 14328 9312 14340
rect 9219 14300 9312 14328
rect 9306 14288 9312 14300
rect 9364 14328 9370 14340
rect 9364 14300 10088 14328
rect 9364 14288 9370 14300
rect 10060 14272 10088 14300
rect 1762 14260 1768 14272
rect 1723 14232 1768 14260
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 2685 14263 2743 14269
rect 2685 14229 2697 14263
rect 2731 14260 2743 14263
rect 2774 14260 2780 14272
rect 2731 14232 2780 14260
rect 2731 14229 2743 14232
rect 2685 14223 2743 14229
rect 2774 14220 2780 14232
rect 2832 14220 2838 14272
rect 3050 14220 3056 14272
rect 3108 14260 3114 14272
rect 3326 14260 3332 14272
rect 3108 14232 3332 14260
rect 3108 14220 3114 14232
rect 3326 14220 3332 14232
rect 3384 14260 3390 14272
rect 5166 14260 5172 14272
rect 3384 14232 5172 14260
rect 3384 14220 3390 14232
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 8846 14260 8852 14272
rect 7800 14232 8852 14260
rect 7800 14220 7806 14232
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 9398 14260 9404 14272
rect 9088 14232 9404 14260
rect 9088 14220 9094 14232
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10704 14260 10732 14368
rect 10980 14328 11008 14436
rect 11149 14433 11161 14467
rect 11195 14464 11207 14467
rect 11195 14436 11560 14464
rect 11195 14433 11207 14436
rect 11149 14427 11207 14433
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 11112 14368 11253 14396
rect 11112 14356 11118 14368
rect 11241 14365 11253 14368
rect 11287 14365 11299 14399
rect 11241 14359 11299 14365
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11532 14396 11560 14436
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11664 14436 11989 14464
rect 11664 14424 11670 14436
rect 11977 14433 11989 14436
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 12308 14436 12541 14464
rect 12308 14424 12314 14436
rect 12529 14433 12541 14436
rect 12575 14433 12587 14467
rect 12529 14427 12587 14433
rect 12796 14467 12854 14473
rect 12796 14433 12808 14467
rect 12842 14464 12854 14467
rect 13814 14464 13820 14476
rect 12842 14436 13820 14464
rect 12842 14433 12854 14436
rect 12796 14427 12854 14433
rect 11698 14396 11704 14408
rect 11388 14368 11481 14396
rect 11532 14368 11704 14396
rect 11388 14356 11394 14368
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12069 14399 12127 14405
rect 12069 14396 12081 14399
rect 11992 14368 12081 14396
rect 11348 14328 11376 14356
rect 11992 14340 12020 14368
rect 12069 14365 12081 14368
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 10980 14300 11376 14328
rect 11974 14288 11980 14340
rect 12032 14288 12038 14340
rect 10962 14260 10968 14272
rect 10100 14232 10968 14260
rect 10100 14220 10106 14232
rect 10962 14220 10968 14232
rect 11020 14260 11026 14272
rect 12176 14260 12204 14359
rect 11020 14232 12204 14260
rect 12544 14260 12572 14427
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 13998 14424 14004 14476
rect 14056 14464 14062 14476
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 14056 14436 14197 14464
rect 14056 14424 14062 14436
rect 14185 14433 14197 14436
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14464 14795 14467
rect 15562 14464 15568 14476
rect 14783 14436 15568 14464
rect 14783 14433 14795 14436
rect 14737 14427 14795 14433
rect 15562 14424 15568 14436
rect 15620 14424 15626 14476
rect 16114 14464 16120 14476
rect 16075 14436 16120 14464
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 18506 14464 18512 14476
rect 16316 14436 18512 14464
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 16022 14396 16028 14408
rect 15059 14368 16028 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16206 14396 16212 14408
rect 16167 14368 16212 14396
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 14369 14331 14427 14337
rect 14369 14297 14381 14331
rect 14415 14328 14427 14331
rect 16316 14328 16344 14436
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 20916 14473 20944 14572
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 19300 14436 19625 14464
rect 19300 14424 19306 14436
rect 19613 14433 19625 14436
rect 19659 14433 19671 14467
rect 19613 14427 19671 14433
rect 20165 14467 20223 14473
rect 20165 14433 20177 14467
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 16574 14396 16580 14408
rect 16439 14368 16580 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17221 14399 17279 14405
rect 17221 14396 17233 14399
rect 17000 14368 17233 14396
rect 17000 14356 17006 14368
rect 17221 14365 17233 14368
rect 17267 14365 17279 14399
rect 17221 14359 17279 14365
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 20180 14396 20208 14427
rect 19944 14368 20208 14396
rect 19944 14356 19950 14368
rect 14415 14300 16344 14328
rect 14415 14297 14427 14300
rect 14369 14291 14427 14297
rect 14001 14263 14059 14269
rect 14001 14260 14013 14263
rect 12544 14232 14013 14260
rect 11020 14220 11026 14232
rect 14001 14229 14013 14232
rect 14047 14229 14059 14263
rect 14001 14223 14059 14229
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 18601 14263 18659 14269
rect 18601 14260 18613 14263
rect 17920 14232 18613 14260
rect 17920 14220 17926 14232
rect 18601 14229 18613 14232
rect 18647 14229 18659 14263
rect 18601 14223 18659 14229
rect 21085 14263 21143 14269
rect 21085 14229 21097 14263
rect 21131 14260 21143 14263
rect 21174 14260 21180 14272
rect 21131 14232 21180 14260
rect 21131 14229 21143 14232
rect 21085 14223 21143 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4798 14056 4804 14068
rect 4203 14028 4804 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 5902 14056 5908 14068
rect 5500 14028 5908 14056
rect 5500 14016 5506 14028
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6086 14016 6092 14068
rect 6144 14056 6150 14068
rect 9493 14059 9551 14065
rect 6144 14028 9444 14056
rect 6144 14016 6150 14028
rect 5997 13991 6055 13997
rect 5997 13957 6009 13991
rect 6043 13988 6055 13991
rect 6362 13988 6368 14000
rect 6043 13960 6368 13988
rect 6043 13957 6055 13960
rect 5997 13951 6055 13957
rect 1964 13892 2912 13920
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13852 1639 13855
rect 1854 13852 1860 13864
rect 1627 13824 1860 13852
rect 1627 13821 1639 13824
rect 1581 13815 1639 13821
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 1964 13861 1992 13892
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13821 2007 13855
rect 1949 13815 2007 13821
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 2096 13824 2237 13852
rect 2096 13812 2102 13824
rect 2225 13821 2237 13824
rect 2271 13821 2283 13855
rect 2225 13815 2283 13821
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2884 13852 2912 13892
rect 3804 13892 4660 13920
rect 3804 13852 3832 13892
rect 2884 13824 3832 13852
rect 2777 13815 2835 13821
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 1765 13719 1823 13725
rect 1765 13716 1777 13719
rect 1728 13688 1777 13716
rect 1728 13676 1734 13688
rect 1765 13685 1777 13688
rect 1811 13685 1823 13719
rect 2792 13716 2820 13815
rect 3878 13812 3884 13864
rect 3936 13852 3942 13864
rect 4062 13852 4068 13864
rect 3936 13824 4068 13852
rect 3936 13812 3942 13824
rect 4062 13812 4068 13824
rect 4120 13852 4126 13864
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 4120 13824 4537 13852
rect 4120 13812 4126 13824
rect 4525 13821 4537 13824
rect 4571 13821 4583 13855
rect 4632 13852 4660 13892
rect 5810 13852 5816 13864
rect 4632 13824 5816 13852
rect 4525 13815 4583 13821
rect 3044 13787 3102 13793
rect 3044 13753 3056 13787
rect 3090 13784 3102 13787
rect 3694 13784 3700 13796
rect 3090 13756 3700 13784
rect 3090 13753 3102 13756
rect 3044 13747 3102 13753
rect 3694 13744 3700 13756
rect 3752 13744 3758 13796
rect 3878 13716 3884 13728
rect 2792 13688 3884 13716
rect 1765 13679 1823 13685
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 4540 13716 4568 13815
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 4792 13787 4850 13793
rect 4792 13753 4804 13787
rect 4838 13784 4850 13787
rect 5534 13784 5540 13796
rect 4838 13756 5540 13784
rect 4838 13753 4850 13756
rect 4792 13747 4850 13753
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 6012 13716 6040 13951
rect 6362 13948 6368 13960
rect 6420 13948 6426 14000
rect 9416 13988 9444 14028
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 10410 14056 10416 14068
rect 9539 14028 10416 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 11054 14056 11060 14068
rect 10704 14028 11060 14056
rect 10704 13988 10732 14028
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 13170 14056 13176 14068
rect 11563 14028 13176 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 16574 14056 16580 14068
rect 16448 14028 16580 14056
rect 16448 14016 16454 14028
rect 16574 14016 16580 14028
rect 16632 14056 16638 14068
rect 16761 14059 16819 14065
rect 16761 14056 16773 14059
rect 16632 14028 16773 14056
rect 16632 14016 16638 14028
rect 16761 14025 16773 14028
rect 16807 14025 16819 14059
rect 16761 14019 16819 14025
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 19705 14059 19763 14065
rect 18095 14028 19564 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 11882 13988 11888 14000
rect 9416 13960 10732 13988
rect 10796 13960 11888 13988
rect 10042 13920 10048 13932
rect 10003 13892 10048 13920
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10410 13880 10416 13932
rect 10468 13920 10474 13932
rect 10796 13920 10824 13960
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 13906 13948 13912 14000
rect 13964 13948 13970 14000
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 18506 13988 18512 14000
rect 17083 13960 18512 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 10962 13920 10968 13932
rect 10468 13892 10824 13920
rect 10923 13892 10968 13920
rect 10468 13880 10474 13892
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11606 13920 11612 13932
rect 11195 13892 11612 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 13924 13920 13952 13948
rect 12207 13892 12572 13920
rect 13924 13892 14044 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 6181 13855 6239 13861
rect 6181 13821 6193 13855
rect 6227 13821 6239 13855
rect 6181 13815 6239 13821
rect 6196 13784 6224 13815
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 7098 13861 7104 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6788 13824 6837 13852
rect 6788 13812 6794 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 7092 13852 7104 13861
rect 7059 13824 7104 13852
rect 6825 13815 6883 13821
rect 7092 13815 7104 13824
rect 7098 13812 7104 13815
rect 7156 13812 7162 13864
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 10226 13852 10232 13864
rect 9999 13824 10232 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 10870 13852 10876 13864
rect 10744 13824 10876 13852
rect 10744 13812 10750 13824
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 12066 13852 12072 13864
rect 11756 13824 12072 13852
rect 11756 13812 11762 13824
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12308 13824 12449 13852
rect 12308 13812 12314 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12544 13852 12572 13892
rect 13814 13852 13820 13864
rect 12544 13824 13820 13852
rect 12437 13815 12495 13821
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13821 13967 13855
rect 14016 13852 14044 13892
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 15381 13923 15439 13929
rect 15381 13920 15393 13923
rect 15252 13892 15393 13920
rect 15252 13880 15258 13892
rect 15381 13889 15393 13892
rect 15427 13889 15439 13923
rect 17681 13923 17739 13929
rect 15381 13883 15439 13889
rect 16408 13892 17632 13920
rect 14165 13855 14223 13861
rect 14165 13852 14177 13855
rect 14016 13824 14177 13852
rect 13909 13815 13967 13821
rect 14165 13821 14177 13824
rect 14211 13821 14223 13855
rect 14165 13815 14223 13821
rect 7650 13784 7656 13796
rect 6196 13756 7656 13784
rect 7650 13744 7656 13756
rect 7708 13744 7714 13796
rect 9861 13787 9919 13793
rect 7760 13756 8524 13784
rect 4540 13688 6040 13716
rect 6270 13676 6276 13728
rect 6328 13716 6334 13728
rect 7760 13716 7788 13756
rect 8202 13716 8208 13728
rect 6328 13688 7788 13716
rect 8163 13688 8208 13716
rect 6328 13676 6334 13688
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8496 13716 8524 13756
rect 9861 13753 9873 13787
rect 9907 13784 9919 13787
rect 10042 13784 10048 13796
rect 9907 13756 10048 13784
rect 9907 13753 9919 13756
rect 9861 13747 9919 13753
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 11146 13784 11152 13796
rect 10244 13756 11152 13784
rect 10244 13716 10272 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 11977 13787 12035 13793
rect 11977 13753 11989 13787
rect 12023 13784 12035 13787
rect 12158 13784 12164 13796
rect 12023 13756 12164 13784
rect 12023 13753 12035 13756
rect 11977 13747 12035 13753
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 12704 13787 12762 13793
rect 12704 13753 12716 13787
rect 12750 13784 12762 13787
rect 13078 13784 13084 13796
rect 12750 13756 13084 13784
rect 12750 13753 12762 13756
rect 12704 13747 12762 13753
rect 13078 13744 13084 13756
rect 13136 13784 13142 13796
rect 13722 13784 13728 13796
rect 13136 13756 13728 13784
rect 13136 13744 13142 13756
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 13924 13784 13952 13815
rect 15212 13784 15240 13880
rect 15654 13861 15660 13864
rect 15648 13815 15660 13861
rect 15712 13852 15718 13864
rect 15712 13824 15748 13852
rect 15654 13812 15660 13815
rect 15712 13812 15718 13824
rect 16022 13812 16028 13864
rect 16080 13852 16086 13864
rect 16408 13852 16436 13892
rect 16080 13824 16436 13852
rect 17604 13852 17632 13892
rect 17681 13889 17693 13923
rect 17727 13920 17739 13923
rect 17862 13920 17868 13932
rect 17727 13892 17868 13920
rect 17727 13889 17739 13892
rect 17681 13883 17739 13889
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18472 13892 18613 13920
rect 18472 13880 18478 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 19058 13880 19064 13932
rect 19116 13920 19122 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19116 13892 19441 13920
rect 19116 13880 19122 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19536 13920 19564 14028
rect 19705 14025 19717 14059
rect 19751 14056 19763 14059
rect 19886 14056 19892 14068
rect 19751 14028 19892 14056
rect 19751 14025 19763 14028
rect 19705 14019 19763 14025
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 19536 13892 20177 13920
rect 19429 13883 19487 13889
rect 20165 13889 20177 13892
rect 20211 13889 20223 13923
rect 20165 13883 20223 13889
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13920 20407 13923
rect 20438 13920 20444 13932
rect 20395 13892 20444 13920
rect 20395 13889 20407 13892
rect 20349 13883 20407 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20714 13920 20720 13932
rect 20675 13892 20720 13920
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 18322 13852 18328 13864
rect 17604 13824 18328 13852
rect 16080 13812 16086 13824
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 20533 13855 20591 13861
rect 18984 13824 20116 13852
rect 16942 13784 16948 13796
rect 13924 13756 16948 13784
rect 16942 13744 16948 13756
rect 17000 13744 17006 13796
rect 17402 13744 17408 13796
rect 17460 13784 17466 13796
rect 18417 13787 18475 13793
rect 17460 13756 17505 13784
rect 17460 13744 17466 13756
rect 18417 13753 18429 13787
rect 18463 13784 18475 13787
rect 18690 13784 18696 13796
rect 18463 13756 18696 13784
rect 18463 13753 18475 13756
rect 18417 13747 18475 13753
rect 18690 13744 18696 13756
rect 18748 13744 18754 13796
rect 8496 13688 10272 13716
rect 10321 13719 10379 13725
rect 10321 13685 10333 13719
rect 10367 13716 10379 13719
rect 10410 13716 10416 13728
rect 10367 13688 10416 13716
rect 10367 13685 10379 13688
rect 10321 13679 10379 13685
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 10686 13716 10692 13728
rect 10647 13688 10692 13716
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 11164 13716 11192 13744
rect 11698 13716 11704 13728
rect 10836 13688 10881 13716
rect 11164 13688 11704 13716
rect 10836 13676 10842 13688
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 11885 13719 11943 13725
rect 11885 13685 11897 13719
rect 11931 13716 11943 13719
rect 13446 13716 13452 13728
rect 11931 13688 13452 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 13814 13716 13820 13728
rect 13727 13688 13820 13716
rect 13814 13676 13820 13688
rect 13872 13716 13878 13728
rect 15010 13716 15016 13728
rect 13872 13688 15016 13716
rect 13872 13676 13878 13688
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 15289 13719 15347 13725
rect 15289 13685 15301 13719
rect 15335 13716 15347 13719
rect 17310 13716 17316 13728
rect 15335 13688 17316 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 17494 13716 17500 13728
rect 17455 13688 17500 13716
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 18877 13719 18935 13725
rect 18564 13688 18609 13716
rect 18564 13676 18570 13688
rect 18877 13685 18889 13719
rect 18923 13716 18935 13719
rect 18984 13716 19012 13824
rect 19245 13787 19303 13793
rect 19245 13753 19257 13787
rect 19291 13784 19303 13787
rect 19978 13784 19984 13796
rect 19291 13756 19984 13784
rect 19291 13753 19303 13756
rect 19245 13747 19303 13753
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 20088 13793 20116 13824
rect 20533 13821 20545 13855
rect 20579 13852 20591 13855
rect 20622 13852 20628 13864
rect 20579 13824 20628 13852
rect 20579 13821 20591 13824
rect 20533 13815 20591 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 20073 13787 20131 13793
rect 20073 13753 20085 13787
rect 20119 13753 20131 13787
rect 20073 13747 20131 13753
rect 19334 13716 19340 13728
rect 18923 13688 19012 13716
rect 19295 13688 19340 13716
rect 18923 13685 18935 13688
rect 18877 13679 18935 13685
rect 19334 13676 19340 13688
rect 19392 13676 19398 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 20346 13716 20352 13728
rect 19576 13688 20352 13716
rect 19576 13676 19582 13688
rect 20346 13676 20352 13688
rect 20404 13676 20410 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2866 13512 2872 13524
rect 1596 13484 2872 13512
rect 1596 13385 1624 13484
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 2961 13515 3019 13521
rect 2961 13481 2973 13515
rect 3007 13512 3019 13515
rect 3510 13512 3516 13524
rect 3007 13484 3516 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3602 13472 3608 13524
rect 3660 13512 3666 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3660 13484 4077 13512
rect 3660 13472 3666 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4890 13512 4896 13524
rect 4851 13484 4896 13512
rect 4065 13475 4123 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 5868 13484 6561 13512
rect 5868 13472 5874 13484
rect 6549 13481 6561 13484
rect 6595 13481 6607 13515
rect 6549 13475 6607 13481
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8665 13515 8723 13521
rect 8665 13512 8677 13515
rect 8343 13484 8677 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8665 13481 8677 13484
rect 8711 13481 8723 13515
rect 8665 13475 8723 13481
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8812 13484 9045 13512
rect 8812 13472 8818 13484
rect 9033 13481 9045 13484
rect 9079 13512 9091 13515
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 9079 13484 9505 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 9493 13475 9551 13481
rect 9692 13484 12265 13512
rect 1854 13444 1860 13456
rect 1815 13416 1860 13444
rect 1854 13404 1860 13416
rect 1912 13404 1918 13456
rect 4525 13447 4583 13453
rect 4525 13413 4537 13447
rect 4571 13444 4583 13447
rect 4571 13416 8340 13444
rect 4571 13413 4583 13416
rect 4525 13407 4583 13413
rect 1581 13379 1639 13385
rect 1581 13345 1593 13379
rect 1627 13345 1639 13379
rect 1581 13339 1639 13345
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2004 13348 2513 13376
rect 2004 13336 2010 13348
rect 2501 13345 2513 13348
rect 2547 13345 2559 13379
rect 2501 13339 2559 13345
rect 2958 13336 2964 13388
rect 3016 13376 3022 13388
rect 3329 13379 3387 13385
rect 3329 13376 3341 13379
rect 3016 13348 3341 13376
rect 3016 13336 3022 13348
rect 3329 13345 3341 13348
rect 3375 13345 3387 13379
rect 3329 13339 3387 13345
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4706 13376 4712 13388
rect 4479 13348 4712 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 5261 13379 5319 13385
rect 5261 13345 5273 13379
rect 5307 13376 5319 13379
rect 6086 13376 6092 13388
rect 5307 13348 5948 13376
rect 6047 13348 6092 13376
rect 5307 13345 5319 13348
rect 5261 13339 5319 13345
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2593 13311 2651 13317
rect 2593 13308 2605 13311
rect 1912 13280 2605 13308
rect 1912 13268 1918 13280
rect 2593 13277 2605 13280
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3421 13311 3479 13317
rect 2832 13280 2877 13308
rect 2832 13268 2838 13280
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 5350 13308 5356 13320
rect 5311 13280 5356 13308
rect 4617 13271 4675 13277
rect 2498 13200 2504 13252
rect 2556 13240 2562 13252
rect 3436 13240 3464 13271
rect 3620 13240 3648 13271
rect 3694 13240 3700 13252
rect 2556 13212 3464 13240
rect 3607 13212 3700 13240
rect 2556 13200 2562 13212
rect 3694 13200 3700 13212
rect 3752 13240 3758 13252
rect 4632 13240 4660 13271
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 5920 13308 5948 13348
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 6227 13348 6684 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 6270 13308 6276 13320
rect 5500 13280 5545 13308
rect 5920 13280 6276 13308
rect 5500 13268 5506 13280
rect 5460 13240 5488 13268
rect 6104 13252 6132 13280
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13308 6423 13311
rect 6546 13308 6552 13320
rect 6411 13280 6552 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 3752 13212 5488 13240
rect 3752 13200 3758 13212
rect 6086 13200 6092 13252
rect 6144 13200 6150 13252
rect 6656 13240 6684 13348
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 6880 13348 6929 13376
rect 6880 13336 6886 13348
rect 6917 13345 6929 13348
rect 6963 13345 6975 13379
rect 8202 13376 8208 13388
rect 8163 13348 8208 13376
rect 6917 13339 6975 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8312 13376 8340 13416
rect 8386 13404 8392 13456
rect 8444 13444 8450 13456
rect 9125 13447 9183 13453
rect 9125 13444 9137 13447
rect 8444 13416 9137 13444
rect 8444 13404 8450 13416
rect 9125 13413 9137 13416
rect 9171 13444 9183 13447
rect 9692 13444 9720 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 12253 13475 12311 13481
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13262 13512 13268 13524
rect 13127 13484 13268 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 13446 13512 13452 13524
rect 13407 13484 13452 13512
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 14090 13512 14096 13524
rect 13863 13484 14096 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 14274 13512 14280 13524
rect 14235 13484 14280 13512
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 14737 13515 14795 13521
rect 14737 13481 14749 13515
rect 14783 13512 14795 13515
rect 15105 13515 15163 13521
rect 15105 13512 15117 13515
rect 14783 13484 15117 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 15105 13481 15117 13484
rect 15151 13481 15163 13515
rect 15105 13475 15163 13481
rect 15289 13515 15347 13521
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 16206 13512 16212 13524
rect 15335 13484 16212 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 16206 13472 16212 13484
rect 16264 13472 16270 13524
rect 16942 13512 16948 13524
rect 16903 13484 16948 13512
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 18414 13472 18420 13524
rect 18472 13512 18478 13524
rect 19058 13512 19064 13524
rect 18472 13484 19064 13512
rect 18472 13472 18478 13484
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20898 13512 20904 13524
rect 20128 13484 20904 13512
rect 20128 13472 20134 13484
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 9171 13416 9720 13444
rect 9171 13413 9183 13416
rect 9125 13407 9183 13413
rect 10870 13404 10876 13456
rect 10928 13444 10934 13456
rect 12802 13444 12808 13456
rect 10928 13416 12808 13444
rect 10928 13404 10934 13416
rect 12802 13404 12808 13416
rect 12860 13404 12866 13456
rect 16485 13447 16543 13453
rect 16485 13444 16497 13447
rect 13464 13416 16497 13444
rect 13464 13388 13492 13416
rect 16485 13413 16497 13416
rect 16531 13413 16543 13447
rect 16960 13444 16988 13472
rect 17586 13444 17592 13456
rect 16960 13416 17592 13444
rect 16485 13407 16543 13413
rect 17586 13404 17592 13416
rect 17644 13444 17650 13456
rect 19076 13444 19104 13472
rect 19398 13447 19456 13453
rect 19398 13444 19410 13447
rect 17644 13416 19012 13444
rect 19076 13416 19410 13444
rect 17644 13404 17650 13416
rect 11054 13376 11060 13388
rect 8312 13348 9628 13376
rect 11015 13348 11060 13376
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 7742 13308 7748 13320
rect 7239 13280 7748 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 6914 13240 6920 13252
rect 6656 13212 6920 13240
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 7024 13240 7052 13271
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 8386 13308 8392 13320
rect 8347 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 9214 13308 9220 13320
rect 9175 13280 9220 13308
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 8294 13240 8300 13252
rect 7024 13212 8300 13240
rect 8294 13200 8300 13212
rect 8352 13200 8358 13252
rect 9600 13240 9628 13348
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13376 13047 13379
rect 13354 13376 13360 13388
rect 13035 13348 13360 13376
rect 13035 13345 13047 13348
rect 12989 13339 13047 13345
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10468 13280 11161 13308
rect 10468 13268 10474 13280
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 11333 13311 11391 13317
rect 11333 13277 11345 13311
rect 11379 13308 11391 13311
rect 11606 13308 11612 13320
rect 11379 13280 11612 13308
rect 11379 13277 11391 13280
rect 11333 13271 11391 13277
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 13004 13308 13032 13339
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 13446 13336 13452 13388
rect 13504 13336 13510 13388
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 13909 13379 13967 13385
rect 13909 13376 13921 13379
rect 13872 13348 13921 13376
rect 13872 13336 13878 13348
rect 13909 13345 13921 13348
rect 13955 13345 13967 13379
rect 14642 13376 14648 13388
rect 14603 13348 14648 13376
rect 13909 13339 13967 13345
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 15654 13376 15660 13388
rect 14752 13348 15148 13376
rect 15615 13348 15660 13376
rect 12575 13280 13032 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13136 13280 13185 13308
rect 13136 13268 13142 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 13630 13308 13636 13320
rect 13320 13280 13636 13308
rect 13320 13268 13326 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 14001 13311 14059 13317
rect 14001 13308 14013 13311
rect 13780 13280 14013 13308
rect 13780 13268 13786 13280
rect 14001 13277 14013 13280
rect 14047 13277 14059 13311
rect 14001 13271 14059 13277
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 14752 13308 14780 13348
rect 14424 13280 14780 13308
rect 14921 13311 14979 13317
rect 14424 13268 14430 13280
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 15010 13308 15016 13320
rect 14967 13280 15016 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 15120 13308 15148 13348
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16942 13376 16948 13388
rect 15896 13348 16948 13376
rect 15896 13336 15902 13348
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17696 13385 17724 13416
rect 17954 13385 17960 13388
rect 17129 13379 17187 13385
rect 17129 13345 17141 13379
rect 17175 13345 17187 13379
rect 17129 13339 17187 13345
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 17948 13339 17960 13385
rect 18012 13376 18018 13388
rect 18984 13376 19012 13416
rect 19398 13413 19410 13416
rect 19444 13413 19456 13447
rect 19398 13407 19456 13413
rect 19153 13379 19211 13385
rect 19153 13376 19165 13379
rect 18012 13348 18048 13376
rect 18984 13348 19165 13376
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 15120 13280 15761 13308
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15856 13308 15884 13336
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15856 13280 15945 13308
rect 15749 13271 15807 13277
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 16574 13308 16580 13320
rect 16535 13280 16580 13308
rect 15933 13271 15991 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 16669 13311 16727 13317
rect 16669 13277 16681 13311
rect 16715 13277 16727 13311
rect 17144 13308 17172 13339
rect 17954 13336 17960 13339
rect 18012 13336 18018 13348
rect 19153 13345 19165 13348
rect 19199 13376 19211 13379
rect 19242 13376 19248 13388
rect 19199 13348 19248 13376
rect 19199 13345 19211 13348
rect 19153 13339 19211 13345
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 20898 13376 20904 13388
rect 20859 13348 20904 13376
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 16669 13271 16727 13277
rect 16868 13280 17172 13308
rect 10594 13240 10600 13252
rect 9600 13212 10600 13240
rect 10594 13200 10600 13212
rect 10652 13200 10658 13252
rect 10689 13243 10747 13249
rect 10689 13209 10701 13243
rect 10735 13240 10747 13243
rect 12621 13243 12679 13249
rect 10735 13212 12572 13240
rect 10735 13209 10747 13212
rect 10689 13203 10747 13209
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 3326 13172 3332 13184
rect 2179 13144 3332 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 5442 13172 5448 13184
rect 5132 13144 5448 13172
rect 5132 13132 5138 13144
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13172 7895 13175
rect 8754 13172 8760 13184
rect 7883 13144 8760 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 8754 13132 8760 13144
rect 8812 13132 8818 13184
rect 9493 13175 9551 13181
rect 9493 13141 9505 13175
rect 9539 13172 9551 13175
rect 10318 13172 10324 13184
rect 9539 13144 10324 13172
rect 9539 13141 9551 13144
rect 9493 13135 9551 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 12253 13175 12311 13181
rect 12253 13141 12265 13175
rect 12299 13172 12311 13175
rect 12434 13172 12440 13184
rect 12299 13144 12440 13172
rect 12299 13141 12311 13144
rect 12253 13135 12311 13141
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 12544 13172 12572 13212
rect 12621 13209 12633 13243
rect 12667 13240 12679 13243
rect 15105 13243 15163 13249
rect 15105 13240 15117 13243
rect 12667 13212 15117 13240
rect 12667 13209 12679 13212
rect 12621 13203 12679 13209
rect 15105 13209 15117 13212
rect 15151 13209 15163 13243
rect 15105 13203 15163 13209
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 16117 13243 16175 13249
rect 16117 13240 16129 13243
rect 15620 13212 16129 13240
rect 15620 13200 15626 13212
rect 16117 13209 16129 13212
rect 16163 13209 16175 13243
rect 16117 13203 16175 13209
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 16684 13240 16712 13271
rect 16448 13212 16712 13240
rect 16448 13200 16454 13212
rect 12802 13172 12808 13184
rect 12544 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 16868 13172 16896 13280
rect 14056 13144 16896 13172
rect 14056 13132 14062 13144
rect 17034 13132 17040 13184
rect 17092 13172 17098 13184
rect 18782 13172 18788 13184
rect 17092 13144 18788 13172
rect 17092 13132 17098 13144
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 20438 13132 20444 13184
rect 20496 13172 20502 13184
rect 20533 13175 20591 13181
rect 20533 13172 20545 13175
rect 20496 13144 20545 13172
rect 20496 13132 20502 13144
rect 20533 13141 20545 13144
rect 20579 13141 20591 13175
rect 20533 13135 20591 13141
rect 20622 13132 20628 13184
rect 20680 13172 20686 13184
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 20680 13144 21097 13172
rect 20680 13132 20686 13144
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 21085 13135 21143 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1762 12968 1768 12980
rect 1723 12940 1768 12968
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 3878 12968 3884 12980
rect 2648 12940 3884 12968
rect 2648 12928 2654 12940
rect 2314 12792 2320 12844
rect 2372 12832 2378 12844
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 2372 12804 2513 12832
rect 2372 12792 2378 12804
rect 2501 12801 2513 12804
rect 2547 12801 2559 12835
rect 2958 12832 2964 12844
rect 2919 12804 2964 12832
rect 2501 12795 2559 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3252 12841 3280 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 5261 12971 5319 12977
rect 5261 12937 5273 12971
rect 5307 12968 5319 12971
rect 5350 12968 5356 12980
rect 5307 12940 5356 12968
rect 5307 12937 5319 12940
rect 5261 12931 5319 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5534 12968 5540 12980
rect 5447 12940 5540 12968
rect 4617 12903 4675 12909
rect 4617 12869 4629 12903
rect 4663 12900 4675 12903
rect 5460 12900 5488 12940
rect 5534 12928 5540 12940
rect 5592 12968 5598 12980
rect 6822 12968 6828 12980
rect 5592 12940 5948 12968
rect 6783 12940 6828 12968
rect 5592 12928 5598 12940
rect 4663 12872 5488 12900
rect 4663 12869 4675 12872
rect 4617 12863 4675 12869
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12801 3295 12835
rect 5718 12832 5724 12844
rect 5679 12804 5724 12832
rect 3237 12795 3295 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 5920 12841 5948 12940
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7650 12968 7656 12980
rect 7611 12940 7656 12968
rect 7650 12928 7656 12940
rect 7708 12928 7714 12980
rect 8202 12928 8208 12980
rect 8260 12968 8266 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 8260 12940 9505 12968
rect 8260 12928 8266 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 10410 12968 10416 12980
rect 10371 12940 10416 12968
rect 9493 12931 9551 12937
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 11112 12940 11253 12968
rect 11112 12928 11118 12940
rect 11241 12937 11253 12940
rect 11287 12937 11299 12971
rect 11241 12931 11299 12937
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13173 12971 13231 12977
rect 12492 12940 12572 12968
rect 12492 12928 12498 12940
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 6914 12900 6920 12912
rect 6788 12872 6920 12900
rect 6788 12860 6794 12872
rect 6914 12860 6920 12872
rect 6972 12900 6978 12912
rect 7190 12900 7196 12912
rect 6972 12872 7196 12900
rect 6972 12860 6978 12872
rect 7190 12860 7196 12872
rect 7248 12900 7254 12912
rect 7248 12872 8064 12900
rect 7248 12860 7254 12872
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12832 5963 12835
rect 6546 12832 6552 12844
rect 5951 12804 6552 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 8036 12841 8064 12872
rect 11514 12860 11520 12912
rect 11572 12900 11578 12912
rect 12250 12900 12256 12912
rect 11572 12872 12256 12900
rect 11572 12860 11578 12872
rect 12250 12860 12256 12872
rect 12308 12860 12314 12912
rect 12544 12900 12572 12940
rect 13173 12937 13185 12971
rect 13219 12968 13231 12971
rect 14734 12968 14740 12980
rect 13219 12940 14740 12968
rect 13219 12937 13231 12940
rect 13173 12931 13231 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15746 12968 15752 12980
rect 15344 12940 15752 12968
rect 15344 12928 15350 12940
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 16172 12940 16405 12968
rect 16172 12928 16178 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 16393 12931 16451 12937
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18506 12968 18512 12980
rect 18095 12940 18512 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 18748 12940 18889 12968
rect 18748 12928 18754 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 18877 12931 18935 12937
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19705 12971 19763 12977
rect 19705 12968 19717 12971
rect 19392 12940 19717 12968
rect 19392 12928 19398 12940
rect 19705 12937 19717 12940
rect 19751 12937 19763 12971
rect 19705 12931 19763 12937
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 20533 12971 20591 12977
rect 20533 12968 20545 12971
rect 20036 12940 20545 12968
rect 20036 12928 20042 12940
rect 20533 12937 20545 12940
rect 20579 12937 20591 12971
rect 20533 12931 20591 12937
rect 14366 12900 14372 12912
rect 12544 12872 14372 12900
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 14645 12903 14703 12909
rect 14645 12869 14657 12903
rect 14691 12900 14703 12903
rect 15102 12900 15108 12912
rect 14691 12872 15108 12900
rect 14691 12869 14703 12872
rect 14645 12863 14703 12869
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 19886 12900 19892 12912
rect 15988 12872 19892 12900
rect 15988 12860 15994 12872
rect 19886 12860 19892 12872
rect 19944 12860 19950 12912
rect 20088 12872 20300 12900
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 9214 12792 9220 12844
rect 9272 12832 9278 12844
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 9272 12804 10057 12832
rect 9272 12792 9278 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10836 12804 10977 12832
rect 10836 12792 10842 12804
rect 10965 12801 10977 12804
rect 11011 12832 11023 12835
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11011 12804 11805 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 11793 12795 11851 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15562 12832 15568 12844
rect 15335 12804 15568 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 16022 12832 16028 12844
rect 15983 12804 16028 12832
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16666 12792 16672 12844
rect 16724 12792 16730 12844
rect 16942 12832 16948 12844
rect 16903 12804 16948 12832
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18012 12804 18613 12832
rect 18012 12792 18018 12804
rect 18601 12801 18613 12804
rect 18647 12832 18659 12835
rect 18690 12832 18696 12844
rect 18647 12804 18696 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 18690 12792 18696 12804
rect 18748 12832 18754 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 18748 12804 19441 12832
rect 18748 12792 18754 12804
rect 19429 12801 19441 12804
rect 19475 12832 19487 12835
rect 20088 12832 20116 12872
rect 20272 12841 20300 12872
rect 19475 12804 20116 12832
rect 20257 12835 20315 12841
rect 19475 12801 19487 12804
rect 19429 12795 19487 12801
rect 20257 12801 20269 12835
rect 20303 12832 20315 12835
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 20303 12804 21097 12832
rect 20303 12801 20315 12804
rect 20257 12795 20315 12801
rect 21085 12801 21097 12804
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 1578 12764 1584 12776
rect 1539 12736 1584 12764
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 7190 12724 7196 12776
rect 7248 12764 7254 12776
rect 7248 12736 7293 12764
rect 7248 12724 7254 12736
rect 7558 12724 7564 12776
rect 7616 12764 7622 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7616 12736 7849 12764
rect 7616 12724 7622 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 8110 12724 8116 12776
rect 8168 12764 8174 12776
rect 8277 12767 8335 12773
rect 8277 12764 8289 12767
rect 8168 12736 8289 12764
rect 8168 12724 8174 12736
rect 8277 12733 8289 12736
rect 8323 12733 8335 12767
rect 8277 12727 8335 12733
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 9916 12736 9965 12764
rect 9916 12724 9922 12736
rect 9953 12733 9965 12736
rect 9999 12764 10011 12767
rect 10594 12764 10600 12776
rect 9999 12736 10600 12764
rect 9999 12733 10011 12736
rect 9953 12727 10011 12733
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 15930 12764 15936 12776
rect 13679 12736 15936 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 15930 12724 15936 12736
rect 15988 12764 15994 12776
rect 16684 12764 16712 12792
rect 15988 12736 16712 12764
rect 15988 12724 15994 12736
rect 17678 12724 17684 12776
rect 17736 12764 17742 12776
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 17736 12736 19349 12764
rect 17736 12724 17742 12736
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 20070 12764 20076 12776
rect 20031 12736 20076 12764
rect 19337 12727 19395 12733
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 20346 12724 20352 12776
rect 20404 12764 20410 12776
rect 20993 12767 21051 12773
rect 20993 12764 21005 12767
rect 20404 12736 21005 12764
rect 20404 12724 20410 12736
rect 20993 12733 21005 12736
rect 21039 12733 21051 12767
rect 20993 12727 21051 12733
rect 2038 12656 2044 12708
rect 2096 12696 2102 12708
rect 3510 12705 3516 12708
rect 2409 12699 2467 12705
rect 2409 12696 2421 12699
rect 2096 12668 2421 12696
rect 2096 12656 2102 12668
rect 2409 12665 2421 12668
rect 2455 12665 2467 12699
rect 2409 12659 2467 12665
rect 3504 12659 3516 12705
rect 3568 12696 3574 12708
rect 5629 12699 5687 12705
rect 3568 12668 3604 12696
rect 3510 12656 3516 12659
rect 3568 12656 3574 12668
rect 5629 12665 5641 12699
rect 5675 12696 5687 12699
rect 5718 12696 5724 12708
rect 5675 12668 5724 12696
rect 5675 12665 5687 12668
rect 5629 12659 5687 12665
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 7098 12656 7104 12708
rect 7156 12696 7162 12708
rect 7285 12699 7343 12705
rect 7285 12696 7297 12699
rect 7156 12668 7297 12696
rect 7156 12656 7162 12668
rect 7285 12665 7297 12668
rect 7331 12665 7343 12699
rect 7285 12659 7343 12665
rect 10226 12656 10232 12708
rect 10284 12696 10290 12708
rect 10781 12699 10839 12705
rect 10781 12696 10793 12699
rect 10284 12668 10793 12696
rect 10284 12656 10290 12668
rect 10781 12665 10793 12668
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 10873 12699 10931 12705
rect 10873 12665 10885 12699
rect 10919 12696 10931 12699
rect 10962 12696 10968 12708
rect 10919 12668 10968 12696
rect 10919 12665 10931 12668
rect 10873 12659 10931 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 11609 12699 11667 12705
rect 11609 12665 11621 12699
rect 11655 12696 11667 12699
rect 12069 12699 12127 12705
rect 12069 12696 12081 12699
rect 11655 12668 12081 12696
rect 11655 12665 11667 12668
rect 11609 12659 11667 12665
rect 12069 12665 12081 12668
rect 12115 12665 12127 12699
rect 12069 12659 12127 12665
rect 13541 12699 13599 12705
rect 13541 12665 13553 12699
rect 13587 12696 13599 12699
rect 14001 12699 14059 12705
rect 14001 12696 14013 12699
rect 13587 12668 14013 12696
rect 13587 12665 13599 12668
rect 13541 12659 13599 12665
rect 14001 12665 14013 12668
rect 14047 12665 14059 12699
rect 14001 12659 14059 12665
rect 15013 12699 15071 12705
rect 15013 12665 15025 12699
rect 15059 12696 15071 12699
rect 15841 12699 15899 12705
rect 15059 12668 15516 12696
rect 15059 12665 15071 12668
rect 15013 12659 15071 12665
rect 1762 12588 1768 12640
rect 1820 12628 1826 12640
rect 2317 12631 2375 12637
rect 2317 12628 2329 12631
rect 1820 12600 2329 12628
rect 1820 12588 1826 12600
rect 2317 12597 2329 12600
rect 2363 12597 2375 12631
rect 2317 12591 2375 12597
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 8478 12628 8484 12640
rect 8260 12600 8484 12628
rect 8260 12588 8266 12600
rect 8478 12588 8484 12600
rect 8536 12628 8542 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8536 12600 9413 12628
rect 8536 12588 8542 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 9861 12631 9919 12637
rect 9861 12597 9873 12631
rect 9907 12628 9919 12631
rect 11054 12628 11060 12640
rect 9907 12600 11060 12628
rect 9907 12597 9919 12600
rect 9861 12591 9919 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11204 12600 11713 12628
rect 11204 12588 11210 12600
rect 11701 12597 11713 12600
rect 11747 12628 11759 12631
rect 12618 12628 12624 12640
rect 11747 12600 12624 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 15102 12628 15108 12640
rect 15063 12600 15108 12628
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 15488 12637 15516 12668
rect 15841 12665 15853 12699
rect 15887 12696 15899 12699
rect 16666 12696 16672 12708
rect 15887 12668 16672 12696
rect 15887 12665 15899 12668
rect 15841 12659 15899 12665
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 16850 12696 16856 12708
rect 16763 12668 16856 12696
rect 16850 12656 16856 12668
rect 16908 12696 16914 12708
rect 17770 12696 17776 12708
rect 16908 12668 17776 12696
rect 16908 12656 16914 12668
rect 17770 12656 17776 12668
rect 17828 12656 17834 12708
rect 18782 12656 18788 12708
rect 18840 12696 18846 12708
rect 19150 12696 19156 12708
rect 18840 12668 19156 12696
rect 18840 12656 18846 12668
rect 19150 12656 19156 12668
rect 19208 12656 19214 12708
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 20901 12699 20959 12705
rect 20901 12696 20913 12699
rect 19484 12668 20913 12696
rect 19484 12656 19490 12668
rect 20901 12665 20913 12668
rect 20947 12665 20959 12699
rect 20901 12659 20959 12665
rect 15473 12631 15531 12637
rect 15473 12597 15485 12631
rect 15519 12597 15531 12631
rect 15473 12591 15531 12597
rect 15933 12631 15991 12637
rect 15933 12597 15945 12631
rect 15979 12628 15991 12631
rect 16114 12628 16120 12640
rect 15979 12600 16120 12628
rect 15979 12597 15991 12600
rect 15933 12591 15991 12597
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 16761 12631 16819 12637
rect 16761 12597 16773 12631
rect 16807 12628 16819 12631
rect 17310 12628 17316 12640
rect 16807 12600 17316 12628
rect 16807 12597 16819 12600
rect 16761 12591 16819 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18417 12631 18475 12637
rect 18417 12628 18429 12631
rect 18012 12600 18429 12628
rect 18012 12588 18018 12600
rect 18417 12597 18429 12600
rect 18463 12597 18475 12631
rect 18417 12591 18475 12597
rect 18509 12631 18567 12637
rect 18509 12597 18521 12631
rect 18555 12628 18567 12631
rect 18598 12628 18604 12640
rect 18555 12600 18604 12628
rect 18555 12597 18567 12600
rect 18509 12591 18567 12597
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 18932 12600 19257 12628
rect 18932 12588 18938 12600
rect 19245 12597 19257 12600
rect 19291 12597 19303 12631
rect 19245 12591 19303 12597
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20165 12631 20223 12637
rect 20165 12628 20177 12631
rect 19392 12600 20177 12628
rect 19392 12588 19398 12600
rect 20165 12597 20177 12600
rect 20211 12597 20223 12631
rect 20165 12591 20223 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3237 12427 3295 12433
rect 3237 12424 3249 12427
rect 2832 12396 3249 12424
rect 2832 12384 2838 12396
rect 3237 12393 3249 12396
rect 3283 12424 3295 12427
rect 3510 12424 3516 12436
rect 3283 12396 3516 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 7374 12424 7380 12436
rect 5592 12396 7380 12424
rect 5592 12384 5598 12396
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 8205 12427 8263 12433
rect 8205 12393 8217 12427
rect 8251 12424 8263 12427
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8251 12396 8585 12424
rect 8251 12393 8263 12396
rect 8205 12387 8263 12393
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 9033 12427 9091 12433
rect 9033 12393 9045 12427
rect 9079 12424 9091 12427
rect 11517 12427 11575 12433
rect 9079 12396 11468 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 3605 12359 3663 12365
rect 3605 12356 3617 12359
rect 1504 12328 3617 12356
rect 1504 12297 1532 12328
rect 3605 12325 3617 12328
rect 3651 12325 3663 12359
rect 3605 12319 3663 12325
rect 4709 12359 4767 12365
rect 4709 12325 4721 12359
rect 4755 12356 4767 12359
rect 4798 12356 4804 12368
rect 4755 12328 4804 12356
rect 4755 12325 4767 12328
rect 4709 12319 4767 12325
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 6730 12356 6736 12368
rect 5040 12328 6736 12356
rect 5040 12316 5046 12328
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 11440 12356 11468 12396
rect 11517 12393 11529 12427
rect 11563 12424 11575 12427
rect 11606 12424 11612 12436
rect 11563 12396 11612 12424
rect 11563 12393 11575 12396
rect 11517 12387 11575 12393
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 13354 12424 13360 12436
rect 11756 12396 13360 12424
rect 11756 12384 11762 12396
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 13998 12424 14004 12436
rect 13771 12396 14004 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 15102 12424 15108 12436
rect 14415 12396 15108 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16390 12424 16396 12436
rect 16264 12396 16396 12424
rect 16264 12384 16270 12396
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 16632 12396 16773 12424
rect 16632 12384 16638 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 16761 12387 16819 12393
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17267 12396 18644 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 11624 12356 11652 12384
rect 11854 12359 11912 12365
rect 11854 12356 11866 12359
rect 6972 12328 9444 12356
rect 11440 12328 11560 12356
rect 11624 12328 11866 12356
rect 6972 12316 6978 12328
rect 2130 12297 2136 12300
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12257 1547 12291
rect 2124 12288 2136 12297
rect 2091 12260 2136 12288
rect 1489 12251 1547 12257
rect 2124 12251 2136 12260
rect 2130 12248 2136 12251
rect 2188 12248 2194 12300
rect 3326 12288 3332 12300
rect 3287 12260 3332 12288
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 5000 12288 5028 12316
rect 4816 12260 5028 12288
rect 4816 12229 4844 12260
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 6356 12291 6414 12297
rect 6356 12288 6368 12291
rect 6236 12260 6368 12288
rect 6236 12248 6242 12260
rect 6356 12257 6368 12260
rect 6402 12288 6414 12291
rect 6402 12260 7328 12288
rect 6402 12257 6414 12260
rect 6356 12251 6414 12257
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12189 6147 12223
rect 7300 12220 7328 12260
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 7432 12260 8125 12288
rect 7432 12248 7438 12260
rect 8113 12257 8125 12260
rect 8159 12288 8171 12291
rect 8478 12288 8484 12300
rect 8159 12260 8484 12288
rect 8159 12257 8171 12260
rect 8113 12251 8171 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8938 12248 8944 12300
rect 8996 12288 9002 12300
rect 8996 12260 9041 12288
rect 8996 12248 9002 12260
rect 8202 12220 8208 12232
rect 7300 12192 8208 12220
rect 6089 12183 6147 12189
rect 1670 12084 1676 12096
rect 1631 12056 1676 12084
rect 1670 12044 1676 12056
rect 1728 12044 1734 12096
rect 1872 12084 1900 12183
rect 3970 12112 3976 12164
rect 4028 12152 4034 12164
rect 4908 12152 4936 12183
rect 4028 12124 4936 12152
rect 4028 12112 4034 12124
rect 2130 12084 2136 12096
rect 1872 12056 2136 12084
rect 2130 12044 2136 12056
rect 2188 12084 2194 12096
rect 2590 12084 2596 12096
rect 2188 12056 2596 12084
rect 2188 12044 2194 12056
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4706 12084 4712 12096
rect 4387 12056 4712 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 6104 12084 6132 12183
rect 8202 12180 8208 12192
rect 8260 12220 8266 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8260 12192 8309 12220
rect 8260 12180 8266 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 9214 12220 9220 12232
rect 9175 12192 9220 12220
rect 8297 12183 8355 12189
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 7466 12152 7472 12164
rect 7379 12124 7472 12152
rect 7466 12112 7472 12124
rect 7524 12152 7530 12164
rect 7834 12152 7840 12164
rect 7524 12124 7840 12152
rect 7524 12112 7530 12124
rect 7834 12112 7840 12124
rect 7892 12112 7898 12164
rect 6270 12084 6276 12096
rect 6104 12056 6276 12084
rect 6270 12044 6276 12056
rect 6328 12084 6334 12096
rect 6822 12084 6828 12096
rect 6328 12056 6828 12084
rect 6328 12044 6334 12056
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12084 7803 12087
rect 8662 12084 8668 12096
rect 7791 12056 8668 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9416 12084 9444 12328
rect 10404 12291 10462 12297
rect 10404 12257 10416 12291
rect 10450 12288 10462 12291
rect 10778 12288 10784 12300
rect 10450 12260 10784 12288
rect 10450 12257 10462 12260
rect 10404 12251 10462 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11532 12288 11560 12328
rect 11854 12325 11866 12328
rect 11900 12325 11912 12359
rect 11854 12319 11912 12325
rect 12158 12316 12164 12368
rect 12216 12356 12222 12368
rect 17862 12365 17868 12368
rect 17129 12359 17187 12365
rect 17129 12356 17141 12359
rect 12216 12328 17141 12356
rect 12216 12316 12222 12328
rect 17129 12325 17141 12328
rect 17175 12325 17187 12359
rect 17856 12356 17868 12365
rect 17823 12328 17868 12356
rect 17129 12319 17187 12325
rect 17856 12319 17868 12328
rect 17862 12316 17868 12319
rect 17920 12316 17926 12368
rect 18616 12356 18644 12396
rect 18690 12384 18696 12436
rect 18748 12424 18754 12436
rect 18969 12427 19027 12433
rect 18969 12424 18981 12427
rect 18748 12396 18981 12424
rect 18748 12384 18754 12396
rect 18969 12393 18981 12396
rect 19015 12393 19027 12427
rect 18969 12387 19027 12393
rect 19061 12427 19119 12433
rect 19061 12393 19073 12427
rect 19107 12424 19119 12427
rect 19426 12424 19432 12436
rect 19107 12396 19432 12424
rect 19107 12393 19119 12396
rect 19061 12387 19119 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 19794 12424 19800 12436
rect 19536 12396 19800 12424
rect 19536 12356 19564 12396
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 18616 12328 19564 12356
rect 19604 12359 19662 12365
rect 19604 12325 19616 12359
rect 19650 12356 19662 12359
rect 20438 12356 20444 12368
rect 19650 12328 20444 12356
rect 19650 12325 19662 12328
rect 19604 12319 19662 12325
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 11698 12288 11704 12300
rect 11532 12260 11704 12288
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 13906 12288 13912 12300
rect 13867 12260 13912 12288
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 14424 12260 14749 12288
rect 14424 12248 14430 12260
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 15378 12288 15384 12300
rect 14737 12251 14795 12257
rect 15028 12260 15384 12288
rect 9858 12220 9864 12232
rect 9692 12192 9864 12220
rect 9692 12084 9720 12192
rect 9858 12180 9864 12192
rect 9916 12220 9922 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9916 12192 10149 12220
rect 9916 12180 9922 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 15028 12229 15056 12260
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15562 12297 15568 12300
rect 15556 12288 15568 12297
rect 15475 12260 15568 12288
rect 15556 12251 15568 12260
rect 15620 12288 15626 12300
rect 16390 12288 16396 12300
rect 15620 12260 16396 12288
rect 15562 12248 15568 12251
rect 15620 12248 15626 12260
rect 16390 12248 16396 12260
rect 16448 12248 16454 12300
rect 17586 12288 17592 12300
rect 17547 12260 17592 12288
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19337 12291 19395 12297
rect 19337 12288 19349 12291
rect 19300 12260 19349 12288
rect 19300 12248 19306 12260
rect 19337 12257 19349 12260
rect 19383 12257 19395 12291
rect 20990 12288 20996 12300
rect 20951 12260 20996 12288
rect 19337 12251 19395 12257
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11572 12192 11621 12220
rect 11572 12180 11578 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 9416 12056 9720 12084
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 10502 12084 10508 12096
rect 10100 12056 10508 12084
rect 10100 12044 10106 12056
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10870 12044 10876 12096
rect 10928 12084 10934 12096
rect 11146 12084 11152 12096
rect 10928 12056 11152 12084
rect 10928 12044 10934 12056
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11624 12084 11652 12183
rect 14844 12152 14872 12183
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 15160 12192 15301 12220
rect 15160 12180 15166 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 16298 12180 16304 12232
rect 16356 12220 16362 12232
rect 16758 12220 16764 12232
rect 16356 12192 16764 12220
rect 16356 12180 16362 12192
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17313 12223 17371 12229
rect 17313 12189 17325 12223
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 15194 12152 15200 12164
rect 14844 12124 15200 12152
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 16669 12155 16727 12161
rect 16669 12121 16681 12155
rect 16715 12152 16727 12155
rect 16942 12152 16948 12164
rect 16715 12124 16948 12152
rect 16715 12121 16727 12124
rect 16669 12115 16727 12121
rect 16942 12112 16948 12124
rect 17000 12152 17006 12164
rect 17328 12152 17356 12183
rect 17000 12124 17356 12152
rect 17000 12112 17006 12124
rect 12342 12084 12348 12096
rect 11624 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12986 12084 12992 12096
rect 12947 12056 12992 12084
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14550 12084 14556 12096
rect 14148 12056 14556 12084
rect 14148 12044 14154 12056
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 18598 12084 18604 12096
rect 17368 12056 18604 12084
rect 17368 12044 17374 12056
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 20530 12044 20536 12096
rect 20588 12084 20594 12096
rect 20717 12087 20775 12093
rect 20717 12084 20729 12087
rect 20588 12056 20729 12084
rect 20588 12044 20594 12056
rect 20717 12053 20729 12056
rect 20763 12053 20775 12087
rect 21174 12084 21180 12096
rect 21135 12056 21180 12084
rect 20717 12047 20775 12053
rect 21174 12044 21180 12056
rect 21232 12044 21238 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 2130 11880 2136 11892
rect 1780 11852 2136 11880
rect 1780 11753 1808 11852
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 5074 11880 5080 11892
rect 4212 11852 5080 11880
rect 4212 11840 4218 11852
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 7098 11880 7104 11892
rect 5951 11852 7104 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7742 11840 7748 11892
rect 7800 11840 7806 11892
rect 8294 11880 8300 11892
rect 8255 11852 8300 11880
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 8938 11880 8944 11892
rect 8536 11852 8944 11880
rect 8536 11840 8542 11852
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 11790 11880 11796 11892
rect 9600 11852 11796 11880
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 7760 11812 7788 11840
rect 8205 11815 8263 11821
rect 8205 11812 8217 11815
rect 6236 11784 6500 11812
rect 7760 11784 8217 11812
rect 6236 11772 6242 11784
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 3936 11716 4261 11744
rect 3936 11704 3942 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4249 11707 4307 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 6472 11753 6500 11784
rect 8205 11781 8217 11784
rect 8251 11781 8263 11815
rect 8205 11775 8263 11781
rect 8303 11784 8892 11812
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11713 5135 11747
rect 6457 11747 6515 11753
rect 5077 11707 5135 11713
rect 5368 11716 6316 11744
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 5092 11676 5120 11707
rect 4028 11648 5120 11676
rect 4028 11636 4034 11648
rect 2032 11611 2090 11617
rect 2032 11577 2044 11611
rect 2078 11608 2090 11611
rect 2130 11608 2136 11620
rect 2078 11580 2136 11608
rect 2078 11577 2090 11580
rect 2032 11571 2090 11577
rect 2130 11568 2136 11580
rect 2188 11568 2194 11620
rect 3786 11568 3792 11620
rect 3844 11608 3850 11620
rect 5368 11608 5396 11716
rect 6288 11685 6316 11716
rect 6457 11713 6469 11747
rect 6503 11713 6515 11747
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 6457 11707 6515 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 8303 11744 8331 11784
rect 8754 11744 8760 11756
rect 7892 11716 8331 11744
rect 8715 11716 8760 11744
rect 7892 11704 7898 11716
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 8864 11753 8892 11784
rect 9600 11753 9628 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 15657 11883 15715 11889
rect 15657 11880 15669 11883
rect 15436 11852 15669 11880
rect 15436 11840 15442 11852
rect 15657 11849 15669 11852
rect 15703 11880 15715 11883
rect 16022 11880 16028 11892
rect 15703 11852 16028 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 16390 11840 16396 11892
rect 16448 11880 16454 11892
rect 17129 11883 17187 11889
rect 17129 11880 17141 11883
rect 16448 11852 17141 11880
rect 16448 11840 16454 11852
rect 17129 11849 17141 11852
rect 17175 11849 17187 11883
rect 17129 11843 17187 11849
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18049 11883 18107 11889
rect 18049 11880 18061 11883
rect 18012 11852 18061 11880
rect 18012 11840 18018 11852
rect 18049 11849 18061 11852
rect 18095 11849 18107 11883
rect 19702 11880 19708 11892
rect 18049 11843 18107 11849
rect 18340 11852 19708 11880
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 10042 11812 10048 11824
rect 9824 11784 10048 11812
rect 9824 11772 9830 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10229 11815 10287 11821
rect 10229 11781 10241 11815
rect 10275 11812 10287 11815
rect 10275 11784 11560 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 9677 11707 9735 11713
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11645 6331 11679
rect 6273 11639 6331 11645
rect 7092 11679 7150 11685
rect 7092 11645 7104 11679
rect 7138 11676 7150 11679
rect 7852 11676 7880 11704
rect 8662 11676 8668 11688
rect 7138 11648 7880 11676
rect 8623 11648 8668 11676
rect 7138 11645 7150 11648
rect 7092 11639 7150 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 9692 11676 9720 11707
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11532 11753 11560 11784
rect 16758 11772 16764 11824
rect 16816 11812 16822 11824
rect 18340 11812 18368 11852
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 16816 11784 18368 11812
rect 16816 11772 16822 11784
rect 18414 11772 18420 11824
rect 18472 11812 18478 11824
rect 19150 11812 19156 11824
rect 18472 11784 19156 11812
rect 18472 11772 18478 11784
rect 19150 11772 19156 11784
rect 19208 11772 19214 11824
rect 11517 11747 11575 11753
rect 10888 11716 11468 11744
rect 8772 11648 9720 11676
rect 10597 11679 10655 11685
rect 6454 11608 6460 11620
rect 3844 11580 5396 11608
rect 5460 11580 6460 11608
rect 3844 11568 3850 11580
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 2372 11512 3157 11540
rect 2372 11500 2378 11512
rect 3145 11509 3157 11512
rect 3191 11509 3203 11543
rect 3694 11540 3700 11552
rect 3655 11512 3700 11540
rect 3145 11503 3203 11509
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 4062 11540 4068 11552
rect 4023 11512 4068 11540
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4212 11512 4257 11540
rect 4212 11500 4218 11512
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4525 11543 4583 11549
rect 4525 11540 4537 11543
rect 4396 11512 4537 11540
rect 4396 11500 4402 11512
rect 4525 11509 4537 11512
rect 4571 11509 4583 11543
rect 4525 11503 4583 11509
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 4672 11512 4905 11540
rect 4672 11500 4678 11512
rect 4893 11509 4905 11512
rect 4939 11540 4951 11543
rect 5460 11540 5488 11580
rect 6454 11568 6460 11580
rect 6512 11568 6518 11620
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 8772 11608 8800 11648
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 10686 11676 10692 11688
rect 10643 11648 10692 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 6788 11580 8800 11608
rect 6788 11568 6794 11580
rect 9030 11568 9036 11620
rect 9088 11608 9094 11620
rect 10888 11608 10916 11716
rect 11440 11685 11468 11716
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11664 11716 11709 11744
rect 11664 11704 11670 11716
rect 17862 11704 17868 11756
rect 17920 11744 17926 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17920 11716 18613 11744
rect 17920 11704 17926 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 18690 11704 18696 11756
rect 18748 11744 18754 11756
rect 19429 11747 19487 11753
rect 19429 11744 19441 11747
rect 18748 11716 19441 11744
rect 18748 11704 18754 11716
rect 19429 11713 19441 11716
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 19702 11704 19708 11756
rect 19760 11744 19766 11756
rect 20165 11747 20223 11753
rect 20165 11744 20177 11747
rect 19760 11716 20177 11744
rect 19760 11704 19766 11716
rect 20165 11713 20177 11716
rect 20211 11713 20223 11747
rect 20346 11744 20352 11756
rect 20307 11716 20352 11744
rect 20165 11707 20223 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11744 20867 11747
rect 20898 11744 20904 11756
rect 20855 11716 20904 11744
rect 20855 11713 20867 11716
rect 20809 11707 20867 11713
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 12400 11648 12449 11676
rect 12400 11636 12406 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12704 11679 12762 11685
rect 12704 11645 12716 11679
rect 12750 11676 12762 11679
rect 12986 11676 12992 11688
rect 12750 11648 12992 11676
rect 12750 11645 12762 11648
rect 12704 11639 12762 11645
rect 12986 11636 12992 11648
rect 13044 11676 13050 11688
rect 13262 11676 13268 11688
rect 13044 11648 13268 11676
rect 13044 11636 13050 11648
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11676 14335 11679
rect 15102 11676 15108 11688
rect 14323 11648 15108 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 15102 11636 15108 11648
rect 15160 11676 15166 11688
rect 16022 11685 16028 11688
rect 15749 11679 15807 11685
rect 15749 11676 15761 11679
rect 15160 11648 15761 11676
rect 15160 11636 15166 11648
rect 15749 11645 15761 11648
rect 15795 11645 15807 11679
rect 16016 11676 16028 11685
rect 15983 11648 16028 11676
rect 15749 11639 15807 11645
rect 16016 11639 16028 11648
rect 16022 11636 16028 11639
rect 16080 11636 16086 11688
rect 18966 11636 18972 11688
rect 19024 11676 19030 11688
rect 19337 11679 19395 11685
rect 19337 11676 19349 11679
rect 19024 11648 19349 11676
rect 19024 11636 19030 11648
rect 19337 11645 19349 11648
rect 19383 11645 19395 11679
rect 20533 11679 20591 11685
rect 20533 11676 20545 11679
rect 19337 11639 19395 11645
rect 20180 11648 20545 11676
rect 9088 11580 10916 11608
rect 14544 11611 14602 11617
rect 9088 11568 9094 11580
rect 14544 11577 14556 11611
rect 14590 11608 14602 11611
rect 15286 11608 15292 11620
rect 14590 11580 15292 11608
rect 14590 11577 14602 11580
rect 14544 11571 14602 11577
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 18414 11608 18420 11620
rect 18375 11580 18420 11608
rect 18414 11568 18420 11580
rect 18472 11568 18478 11620
rect 20073 11611 20131 11617
rect 20073 11608 20085 11611
rect 18892 11580 20085 11608
rect 5626 11540 5632 11552
rect 4939 11512 5488 11540
rect 5587 11512 5632 11540
rect 4939 11509 4951 11512
rect 4893 11503 4951 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 6365 11543 6423 11549
rect 6365 11509 6377 11543
rect 6411 11540 6423 11543
rect 8938 11540 8944 11552
rect 6411 11512 8944 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 9272 11512 9505 11540
rect 9272 11500 9278 11512
rect 9493 11509 9505 11512
rect 9539 11509 9551 11543
rect 9493 11503 9551 11509
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 11057 11543 11115 11549
rect 10744 11512 10789 11540
rect 10744 11500 10750 11512
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 12894 11540 12900 11552
rect 11103 11512 12900 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 17586 11540 17592 11552
rect 17460 11512 17592 11540
rect 17460 11500 17466 11512
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 18506 11540 18512 11552
rect 18467 11512 18512 11540
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 18892 11549 18920 11580
rect 20073 11577 20085 11580
rect 20119 11577 20131 11611
rect 20073 11571 20131 11577
rect 18877 11543 18935 11549
rect 18877 11509 18889 11543
rect 18923 11509 18935 11543
rect 19242 11540 19248 11552
rect 19203 11512 19248 11540
rect 18877 11503 18935 11509
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 19705 11543 19763 11549
rect 19705 11509 19717 11543
rect 19751 11540 19763 11543
rect 20180 11540 20208 11648
rect 20533 11645 20545 11648
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 19751 11512 20208 11540
rect 19751 11509 19763 11512
rect 19705 11503 19763 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1854 11336 1860 11348
rect 1719 11308 1860 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 3694 11336 3700 11348
rect 2179 11308 3700 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4801 11339 4859 11345
rect 4801 11336 4813 11339
rect 4212 11308 4813 11336
rect 4212 11296 4218 11308
rect 4801 11305 4813 11308
rect 4847 11305 4859 11339
rect 4801 11299 4859 11305
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 6457 11339 6515 11345
rect 6457 11336 6469 11339
rect 5684 11308 6469 11336
rect 5684 11296 5690 11308
rect 6457 11305 6469 11308
rect 6503 11305 6515 11339
rect 11606 11336 11612 11348
rect 6457 11299 6515 11305
rect 7484 11308 11612 11336
rect 2041 11271 2099 11277
rect 2041 11237 2053 11271
rect 2087 11268 2099 11271
rect 3234 11268 3240 11280
rect 2087 11240 3240 11268
rect 2087 11237 2099 11240
rect 2041 11231 2099 11237
rect 3234 11228 3240 11240
rect 3292 11228 3298 11280
rect 3602 11228 3608 11280
rect 3660 11268 3666 11280
rect 6549 11271 6607 11277
rect 6549 11268 6561 11271
rect 3660 11240 6561 11268
rect 3660 11228 3666 11240
rect 6549 11237 6561 11240
rect 6595 11237 6607 11271
rect 6549 11231 6607 11237
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2590 11200 2596 11212
rect 2547 11172 2596 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 2768 11203 2826 11209
rect 2768 11169 2780 11203
rect 2814 11200 2826 11203
rect 3142 11200 3148 11212
rect 2814 11172 3148 11200
rect 2814 11169 2826 11172
rect 2768 11163 2826 11169
rect 3142 11160 3148 11172
rect 3200 11200 3206 11212
rect 3970 11200 3976 11212
rect 3200 11172 3976 11200
rect 3200 11160 3206 11172
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 6822 11200 6828 11212
rect 5215 11172 6828 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7484 11209 7512 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 14366 11336 14372 11348
rect 13412 11308 13952 11336
rect 14327 11308 14372 11336
rect 13412 11296 13418 11308
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 9122 11268 9128 11280
rect 8904 11240 9128 11268
rect 8904 11228 8910 11240
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 9490 11228 9496 11280
rect 9548 11268 9554 11280
rect 12888 11271 12946 11277
rect 9548 11240 12839 11268
rect 9548 11228 9554 11240
rect 7834 11209 7840 11212
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7828 11163 7840 11209
rect 7892 11200 7898 11212
rect 10505 11203 10563 11209
rect 7892 11172 7928 11200
rect 7834 11160 7840 11163
rect 7892 11160 7898 11172
rect 10505 11169 10517 11203
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 5258 11132 5264 11144
rect 5219 11104 5264 11132
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 5368 11064 5396 11095
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 6236 11104 6653 11132
rect 6236 11092 6242 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 6972 11104 7573 11132
rect 6972 11092 6978 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 8938 11092 8944 11144
rect 8996 11132 9002 11144
rect 9766 11132 9772 11144
rect 8996 11104 9772 11132
rect 8996 11092 9002 11104
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 4028 11036 5396 11064
rect 6089 11067 6147 11073
rect 4028 11024 4034 11036
rect 6089 11033 6101 11067
rect 6135 11064 6147 11067
rect 7190 11064 7196 11076
rect 6135 11036 7196 11064
rect 6135 11033 6147 11036
rect 6089 11027 6147 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7285 11067 7343 11073
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 7466 11064 7472 11076
rect 7331 11036 7472 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 9490 11024 9496 11076
rect 9548 11064 9554 11076
rect 10134 11064 10140 11076
rect 9548 11036 10140 11064
rect 9548 11024 9554 11036
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10520 11064 10548 11163
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 11664 11172 12265 11200
rect 11664 11160 11670 11172
rect 12253 11169 12265 11172
rect 12299 11200 12311 11203
rect 12710 11200 12716 11212
rect 12299 11172 12716 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 12811 11200 12839 11240
rect 12888 11237 12900 11271
rect 12934 11268 12946 11271
rect 13814 11268 13820 11280
rect 12934 11240 13820 11268
rect 12934 11237 12946 11240
rect 12888 11231 12946 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 13924 11268 13952 11308
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 15289 11339 15347 11345
rect 15289 11336 15301 11339
rect 15252 11308 15301 11336
rect 15252 11296 15258 11308
rect 15289 11305 15301 11308
rect 15335 11305 15347 11339
rect 16114 11336 16120 11348
rect 16075 11308 16120 11336
rect 15289 11299 15347 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 16356 11308 16589 11336
rect 16356 11296 16362 11308
rect 16577 11305 16589 11308
rect 16623 11305 16635 11339
rect 16577 11299 16635 11305
rect 17589 11339 17647 11345
rect 17589 11305 17601 11339
rect 17635 11336 17647 11339
rect 17678 11336 17684 11348
rect 17635 11308 17684 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 17678 11296 17684 11308
rect 17736 11296 17742 11348
rect 18417 11339 18475 11345
rect 18417 11305 18429 11339
rect 18463 11336 18475 11339
rect 19242 11336 19248 11348
rect 18463 11308 19248 11336
rect 18463 11305 18475 11308
rect 18417 11299 18475 11305
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 21082 11336 21088 11348
rect 21043 11308 21088 11336
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 14737 11271 14795 11277
rect 14737 11268 14749 11271
rect 13924 11240 14749 11268
rect 14737 11237 14749 11240
rect 14783 11237 14795 11271
rect 14737 11231 14795 11237
rect 16485 11271 16543 11277
rect 16485 11237 16497 11271
rect 16531 11268 16543 11271
rect 17034 11268 17040 11280
rect 16531 11240 17040 11268
rect 16531 11237 16543 11240
rect 16485 11231 16543 11237
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 18785 11271 18843 11277
rect 18785 11237 18797 11271
rect 18831 11268 18843 11271
rect 19426 11268 19432 11280
rect 18831 11240 19432 11268
rect 18831 11237 18843 11240
rect 18785 11231 18843 11237
rect 19426 11228 19432 11240
rect 19484 11228 19490 11280
rect 19604 11271 19662 11277
rect 19604 11237 19616 11271
rect 19650 11268 19662 11271
rect 19886 11268 19892 11280
rect 19650 11240 19892 11268
rect 19650 11237 19662 11240
rect 19604 11231 19662 11237
rect 19886 11228 19892 11240
rect 19944 11268 19950 11280
rect 20346 11268 20352 11280
rect 19944 11240 20352 11268
rect 19944 11228 19950 11240
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 14550 11200 14556 11212
rect 12811 11172 14556 11200
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 15286 11200 15292 11212
rect 14936 11172 15292 11200
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 12492 11104 12633 11132
rect 12492 11092 12498 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 14936 11141 14964 11172
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15654 11200 15660 11212
rect 15615 11172 15660 11200
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 17420 11172 17969 11200
rect 14829 11135 14887 11141
rect 14829 11132 14841 11135
rect 14424 11104 14841 11132
rect 14424 11092 14430 11104
rect 14829 11101 14841 11104
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15068 11104 15761 11132
rect 15068 11092 15074 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 16390 11132 16396 11144
rect 15887 11104 16396 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 10520 11036 12664 11064
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 5442 10996 5448 11008
rect 5040 10968 5448 10996
rect 5040 10956 5046 10968
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 8938 10996 8944 11008
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 11974 10996 11980 11008
rect 9180 10968 11980 10996
rect 9180 10956 9186 10968
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12636 10996 12664 11036
rect 13556 11036 15240 11064
rect 13556 10996 13584 11036
rect 12636 10968 13584 10996
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 14001 10999 14059 11005
rect 14001 10996 14013 10999
rect 13688 10968 14013 10996
rect 13688 10956 13694 10968
rect 14001 10965 14013 10968
rect 14047 10965 14059 10999
rect 15212 10996 15240 11036
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 15856 11064 15884 11095
rect 16390 11092 16396 11104
rect 16448 11132 16454 11144
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16448 11104 16681 11132
rect 16448 11092 16454 11104
rect 16669 11101 16681 11104
rect 16715 11101 16727 11135
rect 16942 11132 16948 11144
rect 16903 11104 16948 11132
rect 16669 11095 16727 11101
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17420 11141 17448 11172
rect 17957 11169 17969 11172
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 19334 11200 19340 11212
rect 18095 11172 18552 11200
rect 19295 11172 19340 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18524 11144 18552 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 20898 11200 20904 11212
rect 20859 11172 20904 11200
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 17368 11104 17417 11132
rect 17368 11092 17374 11104
rect 17405 11101 17417 11104
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 15344 11036 15884 11064
rect 17328 11036 17816 11064
rect 15344 11024 15350 11036
rect 17328 10996 17356 11036
rect 15212 10968 17356 10996
rect 17788 10996 17816 11036
rect 17862 11024 17868 11076
rect 17920 11064 17926 11076
rect 18156 11064 18184 11095
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 18874 11132 18880 11144
rect 18835 11104 18880 11132
rect 18874 11092 18880 11104
rect 18932 11092 18938 11144
rect 19061 11135 19119 11141
rect 19061 11101 19073 11135
rect 19107 11132 19119 11135
rect 19150 11132 19156 11144
rect 19107 11104 19156 11132
rect 19107 11101 19119 11104
rect 19061 11095 19119 11101
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 17920 11036 18184 11064
rect 17920 11024 17926 11036
rect 19610 10996 19616 11008
rect 17788 10968 19616 10996
rect 14001 10959 14059 10965
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 20714 10996 20720 11008
rect 20675 10968 20720 10996
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 1762 10792 1768 10804
rect 1627 10764 1768 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 3234 10792 3240 10804
rect 3195 10764 3240 10792
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 3786 10752 3792 10804
rect 3844 10792 3850 10804
rect 4893 10795 4951 10801
rect 3844 10764 4844 10792
rect 3844 10752 3850 10764
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4816 10724 4844 10764
rect 4893 10761 4905 10795
rect 4939 10792 4951 10795
rect 5258 10792 5264 10804
rect 4939 10764 5264 10792
rect 4939 10761 4951 10764
rect 4893 10755 4951 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7374 10792 7380 10804
rect 7248 10764 7380 10792
rect 7248 10752 7254 10764
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 9030 10792 9036 10804
rect 8991 10764 9036 10792
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 10778 10792 10784 10804
rect 9692 10764 10784 10792
rect 9122 10724 9128 10736
rect 4028 10696 4660 10724
rect 4816 10696 9128 10724
rect 4028 10684 4034 10696
rect 2130 10656 2136 10668
rect 2043 10628 2136 10656
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3142 10656 3148 10668
rect 3099 10628 3148 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3878 10656 3884 10668
rect 3252 10628 3884 10656
rect 2148 10588 2176 10616
rect 3252 10588 3280 10628
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4632 10665 4660 10696
rect 9122 10684 9128 10696
rect 9180 10684 9186 10736
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5500 10628 5545 10656
rect 5500 10616 5506 10628
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 6052 10628 6285 10656
rect 6052 10616 6058 10628
rect 6273 10625 6285 10628
rect 6319 10656 6331 10659
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 6319 10628 7573 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 8938 10656 8944 10668
rect 8895 10628 8944 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9692 10665 9720 10764
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 11204 10764 11345 10792
rect 11204 10752 11210 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 13354 10792 13360 10804
rect 12483 10764 13360 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 14645 10795 14703 10801
rect 14645 10761 14657 10795
rect 14691 10792 14703 10795
rect 15010 10792 15016 10804
rect 14691 10764 15016 10792
rect 14691 10761 14703 10764
rect 14645 10755 14703 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 16117 10795 16175 10801
rect 16117 10792 16129 10795
rect 15712 10764 16129 10792
rect 15712 10752 15718 10764
rect 16117 10761 16129 10764
rect 16163 10761 16175 10795
rect 16117 10755 16175 10761
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 16945 10795 17003 10801
rect 16945 10792 16957 10795
rect 16724 10764 16957 10792
rect 16724 10752 16730 10764
rect 16945 10761 16957 10764
rect 16991 10761 17003 10795
rect 19886 10792 19892 10804
rect 16945 10755 17003 10761
rect 17144 10764 19472 10792
rect 19847 10764 19892 10792
rect 10796 10724 10824 10752
rect 11241 10727 11299 10733
rect 11241 10724 11253 10727
rect 10796 10696 11253 10724
rect 11241 10693 11253 10696
rect 11287 10693 11299 10727
rect 11241 10687 11299 10693
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 12768 10696 13952 10724
rect 12768 10684 12774 10696
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9858 10656 9864 10668
rect 9819 10628 9864 10656
rect 9677 10619 9735 10625
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11072 10628 11897 10656
rect 2148 10560 3280 10588
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 4246 10588 4252 10600
rect 3743 10560 4252 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 4430 10588 4436 10600
rect 4391 10560 4436 10588
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 5258 10588 5264 10600
rect 5219 10560 5264 10588
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 8662 10588 8668 10600
rect 8623 10560 8668 10588
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 10870 10588 10876 10600
rect 8772 10560 10876 10588
rect 1949 10523 2007 10529
rect 1949 10489 1961 10523
rect 1995 10520 2007 10523
rect 2869 10523 2927 10529
rect 1995 10492 2452 10520
rect 1995 10489 2007 10492
rect 1949 10483 2007 10489
rect 2041 10455 2099 10461
rect 2041 10421 2053 10455
rect 2087 10452 2099 10455
rect 2222 10452 2228 10464
rect 2087 10424 2228 10452
rect 2087 10421 2099 10424
rect 2041 10415 2099 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2424 10461 2452 10492
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 3234 10520 3240 10532
rect 2915 10492 3240 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3234 10480 3240 10492
rect 3292 10480 3298 10532
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 4706 10520 4712 10532
rect 3651 10492 4712 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 4706 10480 4712 10492
rect 4764 10480 4770 10532
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 5353 10523 5411 10529
rect 5353 10520 5365 10523
rect 5040 10492 5365 10520
rect 5040 10480 5046 10492
rect 5353 10489 5365 10492
rect 5399 10489 5411 10523
rect 5353 10483 5411 10489
rect 6638 10480 6644 10532
rect 6696 10520 6702 10532
rect 8772 10520 8800 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 11072 10532 11100 10628
rect 11885 10625 11897 10628
rect 11931 10625 11943 10659
rect 12894 10656 12900 10668
rect 12855 10628 12900 10656
rect 11885 10619 11943 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10656 13047 10659
rect 13262 10656 13268 10668
rect 13035 10628 13268 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 13817 10659 13875 10665
rect 13817 10656 13829 10659
rect 13688 10628 13829 10656
rect 13688 10616 13694 10628
rect 13817 10625 13829 10628
rect 13863 10625 13875 10659
rect 13924 10656 13952 10696
rect 15289 10659 15347 10665
rect 13924 10628 14596 10656
rect 13817 10619 13875 10625
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11204 10560 11713 10588
rect 11204 10548 11210 10560
rect 11701 10557 11713 10560
rect 11747 10588 11759 10591
rect 12434 10588 12440 10600
rect 11747 10560 12440 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12802 10588 12808 10600
rect 12763 10560 12808 10588
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 13078 10548 13084 10600
rect 13136 10588 13142 10600
rect 14274 10588 14280 10600
rect 13136 10560 14280 10588
rect 13136 10548 13142 10560
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 14568 10597 14596 10628
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 15562 10656 15568 10668
rect 15335 10628 15568 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 15562 10616 15568 10628
rect 15620 10656 15626 10668
rect 16761 10659 16819 10665
rect 16761 10656 16773 10659
rect 15620 10628 16773 10656
rect 15620 10616 15626 10628
rect 16761 10625 16773 10628
rect 16807 10656 16819 10659
rect 17144 10656 17172 10764
rect 17310 10684 17316 10736
rect 17368 10724 17374 10736
rect 18230 10724 18236 10736
rect 17368 10696 18236 10724
rect 17368 10684 17374 10696
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 19444 10724 19472 10764
rect 19886 10752 19892 10764
rect 19944 10752 19950 10804
rect 20714 10724 20720 10736
rect 19444 10696 20720 10724
rect 20714 10684 20720 10696
rect 20772 10684 20778 10736
rect 20806 10684 20812 10736
rect 20864 10724 20870 10736
rect 22554 10724 22560 10736
rect 20864 10696 22560 10724
rect 20864 10684 20870 10696
rect 22554 10684 22560 10696
rect 22612 10684 22618 10736
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 16807 10628 17172 10656
rect 17420 10628 17509 10656
rect 16807 10625 16819 10628
rect 16761 10619 16819 10625
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16850 10588 16856 10600
rect 16531 10560 16856 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 17000 10560 17325 10588
rect 17000 10548 17006 10560
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 6696 10492 8800 10520
rect 10128 10523 10186 10529
rect 6696 10480 6702 10492
rect 10128 10489 10140 10523
rect 10174 10520 10186 10523
rect 11054 10520 11060 10532
rect 10174 10492 11060 10520
rect 10174 10489 10186 10492
rect 10128 10483 10186 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11790 10520 11796 10532
rect 11751 10492 11796 10520
rect 11790 10480 11796 10492
rect 11848 10480 11854 10532
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 13633 10523 13691 10529
rect 11940 10492 13308 10520
rect 11940 10480 11946 10492
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10421 2467 10455
rect 2409 10415 2467 10421
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2832 10424 2877 10452
rect 2832 10412 2838 10424
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 3844 10424 4077 10452
rect 3844 10412 3850 10424
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 5258 10452 5264 10464
rect 4571 10424 5264 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5902 10412 5908 10464
rect 5960 10452 5966 10464
rect 6089 10455 6147 10461
rect 6089 10452 6101 10455
rect 5960 10424 6101 10452
rect 5960 10412 5966 10424
rect 6089 10421 6101 10424
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 7006 10452 7012 10464
rect 6236 10424 6281 10452
rect 6967 10424 7012 10452
rect 6236 10412 6242 10424
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7374 10452 7380 10464
rect 7335 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 8202 10452 8208 10464
rect 7524 10424 7569 10452
rect 8163 10424 8208 10452
rect 7524 10412 7530 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8570 10452 8576 10464
rect 8531 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9030 10412 9036 10464
rect 9088 10452 9094 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9088 10424 9413 10452
rect 9088 10412 9094 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 11146 10452 11152 10464
rect 9539 10424 11152 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 13280 10461 13308 10492
rect 13633 10489 13645 10523
rect 13679 10520 13691 10523
rect 14093 10523 14151 10529
rect 14093 10520 14105 10523
rect 13679 10492 14105 10520
rect 13679 10489 13691 10492
rect 13633 10483 13691 10489
rect 14093 10489 14105 10492
rect 14139 10489 14151 10523
rect 15102 10520 15108 10532
rect 15063 10492 15108 10520
rect 14093 10483 14151 10489
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 16390 10480 16396 10532
rect 16448 10520 16454 10532
rect 17420 10520 17448 10628
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 20533 10659 20591 10665
rect 20533 10625 20545 10659
rect 20579 10625 20591 10659
rect 20990 10656 20996 10668
rect 20951 10628 20996 10656
rect 20533 10619 20591 10625
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 16448 10492 17448 10520
rect 16448 10480 16454 10492
rect 17494 10480 17500 10532
rect 17552 10520 17558 10532
rect 18524 10520 18552 10551
rect 19886 10548 19892 10600
rect 19944 10588 19950 10600
rect 20162 10588 20168 10600
rect 19944 10560 20168 10588
rect 19944 10548 19950 10560
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 20346 10588 20352 10600
rect 20307 10560 20352 10588
rect 20346 10548 20352 10560
rect 20404 10548 20410 10600
rect 17552 10492 18552 10520
rect 17552 10480 17558 10492
rect 18690 10480 18696 10532
rect 18748 10529 18754 10532
rect 18748 10523 18812 10529
rect 18748 10489 18766 10523
rect 18800 10520 18812 10523
rect 20548 10520 20576 10619
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 20806 10588 20812 10600
rect 20767 10560 20812 10588
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 18800 10492 20576 10520
rect 18800 10489 18812 10492
rect 18748 10483 18812 10489
rect 18748 10480 18754 10483
rect 13265 10455 13323 10461
rect 13265 10421 13277 10455
rect 13311 10421 13323 10455
rect 13722 10452 13728 10464
rect 13683 10424 13728 10452
rect 13265 10415 13323 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 13964 10424 14381 10452
rect 13964 10412 13970 10424
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 15010 10452 15016 10464
rect 14971 10424 15016 10452
rect 14369 10415 14427 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 16577 10455 16635 10461
rect 16577 10452 16589 10455
rect 15436 10424 16589 10452
rect 15436 10412 15442 10424
rect 16577 10421 16589 10424
rect 16623 10421 16635 10455
rect 16577 10415 16635 10421
rect 16758 10412 16764 10464
rect 16816 10452 16822 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 16816 10424 17417 10452
rect 16816 10412 16822 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 19702 10412 19708 10464
rect 19760 10452 19766 10464
rect 19981 10455 20039 10461
rect 19981 10452 19993 10455
rect 19760 10424 19993 10452
rect 19760 10412 19766 10424
rect 19981 10421 19993 10424
rect 20027 10421 20039 10455
rect 20438 10452 20444 10464
rect 20399 10424 20444 10452
rect 19981 10415 20039 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 1946 10248 1952 10260
rect 1627 10220 1952 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2087 10220 2421 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 2409 10217 2421 10220
rect 2455 10217 2467 10251
rect 2409 10211 2467 10217
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3237 10251 3295 10257
rect 3237 10248 3249 10251
rect 2832 10220 3249 10248
rect 2832 10208 2838 10220
rect 3237 10217 3249 10220
rect 3283 10217 3295 10251
rect 3237 10211 3295 10217
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3786 10248 3792 10260
rect 3568 10220 3792 10248
rect 3568 10208 3574 10220
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 6638 10248 6644 10260
rect 4120 10220 6644 10248
rect 4120 10208 4126 10220
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7466 10248 7472 10260
rect 6963 10220 7472 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 7576 10220 9137 10248
rect 2869 10183 2927 10189
rect 2869 10149 2881 10183
rect 2915 10180 2927 10183
rect 3694 10180 3700 10192
rect 2915 10152 3700 10180
rect 2915 10149 2927 10152
rect 2869 10143 2927 10149
rect 3694 10140 3700 10152
rect 3752 10140 3758 10192
rect 4338 10189 4344 10192
rect 4332 10143 4344 10189
rect 4396 10180 4402 10192
rect 5442 10180 5448 10192
rect 4396 10152 5448 10180
rect 4338 10140 4344 10143
rect 4396 10140 4402 10152
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 6730 10180 6736 10192
rect 6564 10152 6736 10180
rect 1946 10112 1952 10124
rect 1907 10084 1952 10112
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 2823 10084 3372 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3142 10044 3148 10056
rect 3099 10016 3148 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3344 10044 3372 10084
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 6270 10112 6276 10124
rect 3476 10084 5120 10112
rect 6231 10084 6276 10112
rect 3476 10072 3482 10084
rect 3510 10044 3516 10056
rect 3344 10016 3516 10044
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3936 10016 4077 10044
rect 3936 10004 3942 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 5092 10044 5120 10084
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6564 10053 6592 10152
rect 6730 10140 6736 10152
rect 6788 10180 6794 10192
rect 7576 10180 7604 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 10413 10251 10471 10257
rect 10413 10217 10425 10251
rect 10459 10248 10471 10251
rect 10686 10248 10692 10260
rect 10459 10220 10692 10248
rect 10459 10217 10471 10220
rect 10413 10211 10471 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 11241 10251 11299 10257
rect 11241 10248 11253 10251
rect 11204 10220 11253 10248
rect 11204 10208 11210 10220
rect 11241 10217 11253 10220
rect 11287 10217 11299 10251
rect 11241 10211 11299 10217
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 13722 10248 13728 10260
rect 12032 10220 13728 10248
rect 12032 10208 12038 10220
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13832 10220 13921 10248
rect 6788 10152 7604 10180
rect 6788 10140 6794 10152
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 5092 10016 6377 10044
rect 4065 10007 4123 10013
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 2774 9976 2780 9988
rect 2464 9948 2780 9976
rect 2464 9936 2470 9948
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 5902 9976 5908 9988
rect 5863 9948 5908 9976
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 3970 9868 3976 9920
rect 4028 9908 4034 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 4028 9880 5457 9908
rect 4028 9868 4034 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 7300 9908 7328 10075
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 7466 10044 7472 10056
rect 7423 10016 7472 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7576 10053 7604 10152
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 9214 10180 9220 10192
rect 8536 10152 9220 10180
rect 8536 10140 8542 10152
rect 9214 10140 9220 10152
rect 9272 10140 9278 10192
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 10781 10183 10839 10189
rect 10781 10180 10793 10183
rect 10652 10152 10793 10180
rect 10652 10140 10658 10152
rect 10781 10149 10793 10152
rect 10827 10149 10839 10183
rect 11698 10180 11704 10192
rect 11611 10152 11704 10180
rect 10781 10143 10839 10149
rect 11698 10140 11704 10152
rect 11756 10180 11762 10192
rect 13449 10183 13507 10189
rect 13449 10180 13461 10183
rect 11756 10152 13461 10180
rect 11756 10140 11762 10152
rect 13449 10149 13461 10152
rect 13495 10149 13507 10183
rect 13832 10180 13860 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 14001 10251 14059 10257
rect 14001 10217 14013 10251
rect 14047 10248 14059 10251
rect 14090 10248 14096 10260
rect 14047 10220 14096 10248
rect 14047 10217 14059 10220
rect 14001 10211 14059 10217
rect 14090 10208 14096 10220
rect 14148 10248 14154 10260
rect 14148 10220 15424 10248
rect 14148 10208 14154 10220
rect 13449 10143 13507 10149
rect 13740 10152 13860 10180
rect 15396 10180 15424 10220
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 16298 10248 16304 10260
rect 15804 10220 16304 10248
rect 15804 10208 15810 10220
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 16448 10220 16681 10248
rect 16448 10208 16454 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18748 10220 18889 10248
rect 18748 10208 18754 10220
rect 18877 10217 18889 10220
rect 18923 10217 18935 10251
rect 18877 10211 18935 10217
rect 19613 10251 19671 10257
rect 19613 10217 19625 10251
rect 19659 10248 19671 10251
rect 20346 10248 20352 10260
rect 19659 10220 20352 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 16022 10180 16028 10192
rect 15396 10152 16028 10180
rect 13740 10124 13768 10152
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 17764 10183 17822 10189
rect 17764 10149 17776 10183
rect 17810 10180 17822 10183
rect 17954 10180 17960 10192
rect 17810 10152 17960 10180
rect 17810 10149 17822 10152
rect 17764 10143 17822 10149
rect 17954 10140 17960 10152
rect 18012 10180 18018 10192
rect 19150 10180 19156 10192
rect 18012 10152 19156 10180
rect 18012 10140 18018 10152
rect 19150 10140 19156 10152
rect 19208 10180 19214 10192
rect 19208 10152 20208 10180
rect 19208 10140 19214 10152
rect 8012 10115 8070 10121
rect 8012 10081 8024 10115
rect 8058 10112 8070 10115
rect 8938 10112 8944 10124
rect 8058 10084 8944 10112
rect 8058 10081 8070 10084
rect 8012 10075 8070 10081
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 10318 10072 10324 10124
rect 10376 10112 10382 10124
rect 10873 10115 10931 10121
rect 10873 10112 10885 10115
rect 10376 10084 10885 10112
rect 10376 10072 10382 10084
rect 10873 10081 10885 10084
rect 10919 10081 10931 10115
rect 10873 10075 10931 10081
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 11146 10112 11152 10124
rect 11020 10084 11152 10112
rect 11020 10072 11026 10084
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12860 10084 13001 10112
rect 12860 10072 12866 10084
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13722 10072 13728 10124
rect 13780 10072 13786 10124
rect 14366 10072 14372 10124
rect 14424 10072 14430 10124
rect 14734 10112 14740 10124
rect 14695 10084 14740 10112
rect 14734 10072 14740 10084
rect 14792 10072 14798 10124
rect 15562 10121 15568 10124
rect 15556 10112 15568 10121
rect 15028 10084 15568 10112
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7561 10007 7619 10013
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10778 10044 10784 10056
rect 9824 10016 10784 10044
rect 9824 10004 9830 10016
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 11054 10044 11060 10056
rect 11015 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 11072 9976 11100 10004
rect 11808 9976 11836 10007
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 13078 10044 13084 10056
rect 12676 10016 13084 10044
rect 12676 10004 12682 10016
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 13262 10044 13268 10056
rect 13175 10016 13268 10044
rect 13262 10004 13268 10016
rect 13320 10044 13326 10056
rect 13630 10044 13636 10056
rect 13320 10016 13636 10044
rect 13320 10004 13326 10016
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 13998 10044 14004 10056
rect 13872 10016 14004 10044
rect 13872 10004 13878 10016
rect 13998 10004 14004 10016
rect 14056 10044 14062 10056
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 14056 10016 14197 10044
rect 14056 10004 14062 10016
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 12526 9976 12532 9988
rect 11072 9948 11836 9976
rect 11900 9948 12532 9976
rect 8478 9908 8484 9920
rect 7300 9880 8484 9908
rect 5445 9871 5503 9877
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 11900 9908 11928 9948
rect 12526 9936 12532 9948
rect 12584 9936 12590 9988
rect 13449 9979 13507 9985
rect 13449 9945 13461 9979
rect 13495 9976 13507 9979
rect 14090 9976 14096 9988
rect 13495 9948 14096 9976
rect 13495 9945 13507 9948
rect 13449 9939 13507 9945
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 14384 9985 14412 10072
rect 15028 10053 15056 10084
rect 15556 10075 15568 10084
rect 15562 10072 15568 10075
rect 15620 10072 15626 10124
rect 19978 10112 19984 10124
rect 19939 10084 19984 10112
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 15013 10047 15071 10053
rect 15013 10013 15025 10047
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 17494 10044 17500 10056
rect 15289 10007 15347 10013
rect 17328 10016 17500 10044
rect 14369 9979 14427 9985
rect 14369 9945 14381 9979
rect 14415 9945 14427 9979
rect 14844 9976 14872 10007
rect 15194 9976 15200 9988
rect 14844 9948 15200 9976
rect 14369 9939 14427 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 11848 9880 11928 9908
rect 11848 9868 11854 9880
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12032 9880 12633 9908
rect 12032 9868 12038 9880
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 12621 9871 12679 9877
rect 13541 9911 13599 9917
rect 13541 9877 13553 9911
rect 13587 9908 13599 9911
rect 15102 9908 15108 9920
rect 13587 9880 15108 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15304 9908 15332 10007
rect 15654 9908 15660 9920
rect 15304 9880 15660 9908
rect 15654 9868 15660 9880
rect 15712 9908 15718 9920
rect 17328 9908 17356 10016
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 20070 10044 20076 10056
rect 20031 10016 20076 10044
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20180 10053 20208 10152
rect 20165 10047 20223 10053
rect 20165 10013 20177 10047
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 15712 9880 17356 9908
rect 15712 9868 15718 9880
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 2133 9707 2191 9713
rect 2133 9704 2145 9707
rect 2004 9676 2145 9704
rect 2004 9664 2010 9676
rect 2133 9673 2145 9676
rect 2179 9673 2191 9707
rect 3142 9704 3148 9716
rect 2133 9667 2191 9673
rect 2792 9676 3148 9704
rect 2792 9577 2820 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4341 9707 4399 9713
rect 4341 9704 4353 9707
rect 4304 9676 4353 9704
rect 4304 9664 4310 9676
rect 4341 9673 4353 9676
rect 4387 9673 4399 9707
rect 4341 9667 4399 9673
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 6052 9676 8217 9704
rect 6052 9664 6058 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8205 9667 8263 9673
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 12802 9704 12808 9716
rect 8352 9676 12808 9704
rect 8352 9664 8358 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 14292 9676 14688 9704
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8536 9608 8585 9636
rect 8536 9596 8542 9608
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 10318 9636 10324 9648
rect 8573 9599 8631 9605
rect 8680 9608 10324 9636
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 6270 9568 6276 9580
rect 6231 9540 6276 9568
rect 2777 9531 2835 9537
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2038 9500 2044 9512
rect 1811 9472 2044 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2038 9460 2044 9472
rect 2096 9460 2102 9512
rect 2498 9500 2504 9512
rect 2459 9472 2504 9500
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 4801 9503 4859 9509
rect 3007 9472 3924 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 3896 9444 3924 9472
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 5068 9503 5126 9509
rect 5068 9469 5080 9503
rect 5114 9500 5126 9503
rect 5994 9500 6000 9512
rect 5114 9472 6000 9500
rect 5114 9469 5126 9472
rect 5068 9463 5126 9469
rect 1964 9404 3004 9432
rect 1964 9373 1992 9404
rect 2976 9376 3004 9404
rect 3050 9392 3056 9444
rect 3108 9432 3114 9444
rect 3206 9435 3264 9441
rect 3206 9432 3218 9435
rect 3108 9404 3218 9432
rect 3108 9392 3114 9404
rect 3206 9401 3218 9404
rect 3252 9401 3264 9435
rect 3206 9395 3264 9401
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4062 9432 4068 9444
rect 3936 9404 4068 9432
rect 3936 9392 3942 9404
rect 4062 9392 4068 9404
rect 4120 9432 4126 9444
rect 4816 9432 4844 9463
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6104 9472 6837 9500
rect 6104 9432 6132 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 7616 9472 8493 9500
rect 7616 9460 7622 9472
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 4120 9404 6132 9432
rect 4120 9392 4126 9404
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 7070 9435 7128 9441
rect 7070 9432 7082 9435
rect 6788 9404 7082 9432
rect 6788 9392 6794 9404
rect 7070 9401 7082 9404
rect 7116 9401 7128 9435
rect 8680 9432 8708 9608
rect 10318 9596 10324 9608
rect 10376 9636 10382 9648
rect 10962 9636 10968 9648
rect 10376 9608 10968 9636
rect 10376 9596 10382 9608
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 11517 9639 11575 9645
rect 11517 9605 11529 9639
rect 11563 9605 11575 9639
rect 11517 9599 11575 9605
rect 13909 9639 13967 9645
rect 13909 9605 13921 9639
rect 13955 9636 13967 9639
rect 14292 9636 14320 9676
rect 14660 9636 14688 9676
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 17494 9704 17500 9716
rect 15252 9676 17500 9704
rect 15252 9664 15258 9676
rect 17494 9664 17500 9676
rect 17552 9704 17558 9716
rect 17552 9676 19564 9704
rect 17552 9664 17558 9676
rect 15565 9639 15623 9645
rect 13955 9608 14320 9636
rect 14384 9608 14596 9636
rect 14660 9608 15424 9636
rect 13955 9605 13967 9608
rect 13909 9599 13967 9605
rect 8938 9528 8944 9580
rect 8996 9568 9002 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8996 9540 9137 9568
rect 8996 9528 9002 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 9916 9540 10057 9568
rect 9916 9528 9922 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 11330 9568 11336 9580
rect 11291 9540 11336 9568
rect 10045 9531 10103 9537
rect 11330 9528 11336 9540
rect 11388 9528 11394 9580
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11532 9568 11560 9599
rect 11974 9568 11980 9580
rect 11480 9540 11560 9568
rect 11935 9540 11980 9568
rect 11480 9528 11486 9540
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12158 9568 12164 9580
rect 12119 9540 12164 9568
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14384 9568 14412 9608
rect 14568 9577 14596 9608
rect 14056 9540 14412 9568
rect 14553 9571 14611 9577
rect 14056 9528 14062 9540
rect 14553 9537 14565 9571
rect 14599 9537 14611 9571
rect 14553 9531 14611 9537
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 14976 9540 15301 9568
rect 14976 9528 14982 9540
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9490 9500 9496 9512
rect 9079 9472 9496 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9490 9460 9496 9472
rect 9548 9500 9554 9512
rect 11149 9503 11207 9509
rect 9548 9472 11008 9500
rect 9548 9460 9554 9472
rect 8938 9432 8944 9444
rect 7070 9395 7128 9401
rect 7208 9404 8708 9432
rect 8899 9404 8944 9432
rect 1949 9367 2007 9373
rect 1949 9333 1961 9367
rect 1995 9333 2007 9367
rect 1949 9327 2007 9333
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 2682 9364 2688 9376
rect 2639 9336 2688 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 6052 9336 6193 9364
rect 6052 9324 6058 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 7208 9364 7236 9404
rect 8938 9392 8944 9404
rect 8996 9392 9002 9444
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9432 9919 9435
rect 10502 9432 10508 9444
rect 9907 9404 10508 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 6880 9336 7236 9364
rect 6880 9324 6886 9336
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 8260 9336 8309 9364
rect 8260 9324 8266 9336
rect 8297 9333 8309 9336
rect 8343 9333 8355 9367
rect 9490 9364 9496 9376
rect 9451 9336 9496 9364
rect 8297 9327 8355 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10689 9367 10747 9373
rect 10008 9336 10053 9364
rect 10008 9324 10014 9336
rect 10689 9333 10701 9367
rect 10735 9364 10747 9367
rect 10870 9364 10876 9376
rect 10735 9336 10876 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 10980 9364 11008 9472
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11882 9500 11888 9512
rect 11195 9472 11744 9500
rect 11843 9472 11888 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11057 9435 11115 9441
rect 11057 9401 11069 9435
rect 11103 9432 11115 9435
rect 11422 9432 11428 9444
rect 11103 9404 11428 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 11716 9432 11744 9472
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 12434 9500 12440 9512
rect 12395 9472 12440 9500
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 15102 9500 15108 9512
rect 15063 9472 15108 9500
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15396 9500 15424 9608
rect 15565 9605 15577 9639
rect 15611 9636 15623 9639
rect 17678 9636 17684 9648
rect 15611 9608 17684 9636
rect 15611 9605 15623 9608
rect 15565 9599 15623 9605
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 18049 9639 18107 9645
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 18874 9636 18880 9648
rect 18095 9608 18880 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 18874 9596 18880 9608
rect 18932 9596 18938 9648
rect 19426 9636 19432 9648
rect 19387 9608 19432 9636
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 19536 9636 19564 9676
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 20257 9707 20315 9713
rect 20257 9704 20269 9707
rect 20036 9676 20269 9704
rect 20036 9664 20042 9676
rect 20257 9673 20269 9676
rect 20303 9673 20315 9707
rect 20257 9667 20315 9673
rect 19536 9608 20944 9636
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15528 9540 16037 9568
rect 15528 9528 15534 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 16758 9568 16764 9580
rect 16255 9540 16764 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 16758 9528 16764 9540
rect 16816 9568 16822 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16816 9540 17049 9568
rect 16816 9528 16822 9540
rect 17037 9537 17049 9540
rect 17083 9568 17095 9571
rect 18693 9571 18751 9577
rect 18693 9568 18705 9571
rect 17083 9540 18705 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 18693 9537 18705 9540
rect 18739 9568 18751 9571
rect 19334 9568 19340 9580
rect 18739 9540 19340 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 19334 9528 19340 9540
rect 19392 9568 19398 9580
rect 19981 9571 20039 9577
rect 19981 9568 19993 9571
rect 19392 9540 19993 9568
rect 19392 9528 19398 9540
rect 19981 9537 19993 9540
rect 20027 9568 20039 9571
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 20027 9540 20821 9568
rect 20027 9537 20039 9540
rect 19981 9531 20039 9537
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 17310 9500 17316 9512
rect 15243 9472 15424 9500
rect 15856 9472 17316 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 11974 9432 11980 9444
rect 11716 9404 11980 9432
rect 11974 9392 11980 9404
rect 12032 9392 12038 9444
rect 12704 9435 12762 9441
rect 12704 9401 12716 9435
rect 12750 9432 12762 9435
rect 13262 9432 13268 9444
rect 12750 9404 13268 9432
rect 12750 9401 12762 9404
rect 12704 9395 12762 9401
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 14369 9435 14427 9441
rect 13363 9404 13952 9432
rect 13363 9364 13391 9404
rect 13814 9364 13820 9376
rect 10980 9336 13391 9364
rect 13775 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 13924 9364 13952 9404
rect 14369 9401 14381 9435
rect 14415 9432 14427 9435
rect 14458 9432 14464 9444
rect 14415 9404 14464 9432
rect 14415 9401 14427 9404
rect 14369 9395 14427 9401
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 15856 9432 15884 9472
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 18417 9503 18475 9509
rect 18417 9469 18429 9503
rect 18463 9500 18475 9503
rect 18782 9500 18788 9512
rect 18463 9472 18788 9500
rect 18463 9469 18475 9472
rect 18417 9463 18475 9469
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 19794 9460 19800 9512
rect 19852 9500 19858 9512
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 19852 9472 20637 9500
rect 19852 9460 19858 9472
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 20717 9503 20775 9509
rect 20717 9469 20729 9503
rect 20763 9500 20775 9503
rect 20916 9500 20944 9608
rect 21358 9596 21364 9648
rect 21416 9596 21422 9648
rect 21376 9568 21404 9596
rect 21542 9568 21548 9580
rect 21376 9540 21548 9568
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 20763 9472 20944 9500
rect 20763 9469 20775 9472
rect 20717 9463 20775 9469
rect 14559 9404 15884 9432
rect 15933 9435 15991 9441
rect 14277 9367 14335 9373
rect 14277 9364 14289 9367
rect 13924 9336 14289 9364
rect 14277 9333 14289 9336
rect 14323 9364 14335 9367
rect 14559 9364 14587 9404
rect 15933 9401 15945 9435
rect 15979 9432 15991 9435
rect 16114 9432 16120 9444
rect 15979 9404 16120 9432
rect 15979 9401 15991 9404
rect 15933 9395 15991 9401
rect 16114 9392 16120 9404
rect 16172 9392 16178 9444
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 16684 9404 16865 9432
rect 14323 9336 14587 9364
rect 14737 9367 14795 9373
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 14737 9333 14749 9367
rect 14783 9364 14795 9367
rect 15194 9364 15200 9376
rect 14783 9336 15200 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 16390 9364 16396 9376
rect 16351 9336 16396 9364
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 16684 9364 16712 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 16853 9395 16911 9401
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 19978 9432 19984 9444
rect 19300 9404 19984 9432
rect 19300 9392 19306 9404
rect 19978 9392 19984 9404
rect 20036 9392 20042 9444
rect 16632 9336 16712 9364
rect 16761 9367 16819 9373
rect 16632 9324 16638 9336
rect 16761 9333 16773 9367
rect 16807 9364 16819 9367
rect 16942 9364 16948 9376
rect 16807 9336 16948 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 17276 9336 18521 9364
rect 17276 9324 17282 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 19794 9364 19800 9376
rect 19755 9336 19800 9364
rect 18509 9327 18567 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 19886 9324 19892 9376
rect 19944 9364 19950 9376
rect 19944 9336 19989 9364
rect 19944 9324 19950 9336
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 20530 9364 20536 9376
rect 20220 9336 20536 9364
rect 20220 9324 20226 9336
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2409 9163 2467 9169
rect 2409 9160 2421 9163
rect 2280 9132 2421 9160
rect 2280 9120 2286 9132
rect 2409 9129 2421 9132
rect 2455 9129 2467 9163
rect 2409 9123 2467 9129
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 3384 9132 5365 9160
rect 3384 9120 3390 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 5718 9160 5724 9172
rect 5679 9132 5724 9160
rect 5353 9123 5411 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 6236 9132 6285 9160
rect 6236 9120 6242 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 6273 9123 6331 9129
rect 6733 9163 6791 9169
rect 6733 9129 6745 9163
rect 6779 9160 6791 9163
rect 6822 9160 6828 9172
rect 6779 9132 6828 9160
rect 6779 9129 6791 9132
rect 6733 9123 6791 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7374 9160 7380 9172
rect 7331 9132 7380 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7745 9163 7803 9169
rect 7745 9129 7757 9163
rect 7791 9160 7803 9163
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7791 9132 8125 9160
rect 7791 9129 7803 9132
rect 7745 9123 7803 9129
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 9582 9160 9588 9172
rect 8113 9123 8171 9129
rect 8496 9132 9588 9160
rect 2777 9095 2835 9101
rect 2777 9061 2789 9095
rect 2823 9092 2835 9095
rect 2958 9092 2964 9104
rect 2823 9064 2964 9092
rect 2823 9061 2835 9064
rect 2777 9055 2835 9061
rect 2958 9052 2964 9064
rect 3016 9092 3022 9104
rect 3418 9092 3424 9104
rect 3016 9064 3424 9092
rect 3016 9052 3022 9064
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 5813 9095 5871 9101
rect 5813 9061 5825 9095
rect 5859 9092 5871 9095
rect 7006 9092 7012 9104
rect 5859 9064 7012 9092
rect 5859 9061 5871 9064
rect 5813 9055 5871 9061
rect 7006 9052 7012 9064
rect 7064 9052 7070 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 8496 9101 8524 9132
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 11756 9132 13645 9160
rect 11756 9120 11762 9132
rect 13633 9129 13645 9132
rect 13679 9160 13691 9163
rect 13679 9132 14504 9160
rect 13679 9129 13691 9132
rect 13633 9123 13691 9129
rect 8481 9095 8539 9101
rect 8481 9092 8493 9095
rect 7616 9064 8493 9092
rect 7616 9052 7622 9064
rect 8481 9061 8493 9064
rect 8527 9061 8539 9095
rect 8481 9055 8539 9061
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 10962 9092 10968 9104
rect 8628 9064 8673 9092
rect 9784 9064 10968 9092
rect 8628 9052 8634 9064
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 9024 2927 9027
rect 2915 8996 3464 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3142 8956 3148 8968
rect 3099 8928 3148 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3436 8956 3464 8996
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 6641 9027 6699 9033
rect 6641 9024 6653 9027
rect 3568 8996 6653 9024
rect 3568 8984 3574 8996
rect 6641 8993 6653 8996
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 7156 8996 7665 9024
rect 7156 8984 7162 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 9784 9024 9812 9064
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 11968 9095 12026 9101
rect 11968 9061 11980 9095
rect 12014 9092 12026 9095
rect 12158 9092 12164 9104
rect 12014 9064 12164 9092
rect 12014 9061 12026 9064
rect 11968 9055 12026 9061
rect 12158 9052 12164 9064
rect 12216 9092 12222 9104
rect 13814 9092 13820 9104
rect 12216 9064 13820 9092
rect 12216 9052 12222 9064
rect 13814 9052 13820 9064
rect 13872 9092 13878 9104
rect 14366 9092 14372 9104
rect 13872 9064 14136 9092
rect 14327 9064 14372 9092
rect 13872 9052 13878 9064
rect 8352 8996 9812 9024
rect 9944 9027 10002 9033
rect 8352 8984 8358 8996
rect 9944 8993 9956 9027
rect 9990 9024 10002 9027
rect 9990 8996 10723 9024
rect 9990 8993 10002 8996
rect 9944 8987 10002 8993
rect 3602 8956 3608 8968
rect 3436 8928 3608 8956
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6788 8928 6837 8956
rect 6788 8916 6794 8928
rect 6825 8925 6837 8928
rect 6871 8956 6883 8959
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 6871 8928 7849 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 7837 8925 7849 8928
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 8846 8956 8852 8968
rect 8803 8928 8852 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 9674 8956 9680 8968
rect 9635 8928 9680 8956
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 10695 8956 10723 8996
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 13446 9024 13452 9036
rect 10928 8996 13452 9024
rect 10928 8984 10934 8996
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 11054 8956 11060 8968
rect 10695 8928 11060 8956
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11698 8956 11704 8968
rect 11659 8928 11704 8956
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 12802 8916 12808 8968
rect 12860 8916 12866 8968
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13556 8956 13584 8987
rect 12952 8928 13584 8956
rect 13817 8959 13875 8965
rect 12952 8916 12958 8928
rect 13817 8925 13829 8959
rect 13863 8956 13875 8959
rect 13998 8956 14004 8968
rect 13863 8928 14004 8956
rect 13863 8925 13875 8928
rect 13817 8919 13875 8925
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 14108 8956 14136 9064
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 14476 9092 14504 9132
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 15194 9160 15200 9172
rect 15068 9132 15200 9160
rect 15068 9120 15074 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15381 9163 15439 9169
rect 15381 9129 15393 9163
rect 15427 9160 15439 9163
rect 15470 9160 15476 9172
rect 15427 9132 15476 9160
rect 15427 9129 15439 9132
rect 15381 9123 15439 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15746 9160 15752 9172
rect 15707 9132 15752 9160
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 18012 9132 18061 9160
rect 18012 9120 18018 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 18509 9163 18567 9169
rect 18509 9129 18521 9163
rect 18555 9160 18567 9163
rect 18598 9160 18604 9172
rect 18555 9132 18604 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 18598 9120 18604 9132
rect 18656 9160 18662 9172
rect 18874 9160 18880 9172
rect 18656 9132 18880 9160
rect 18656 9120 18662 9132
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 19981 9163 20039 9169
rect 19981 9129 19993 9163
rect 20027 9160 20039 9163
rect 20070 9160 20076 9172
rect 20027 9132 20076 9160
rect 20027 9129 20039 9132
rect 19981 9123 20039 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 16666 9092 16672 9104
rect 14476 9064 16672 9092
rect 16666 9052 16672 9064
rect 16724 9052 16730 9104
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 16914 9095 16972 9101
rect 16914 9092 16926 9095
rect 16816 9064 16926 9092
rect 16816 9052 16822 9064
rect 16914 9061 16926 9064
rect 16960 9061 16972 9095
rect 19426 9092 19432 9104
rect 16914 9055 16972 9061
rect 17032 9064 19432 9092
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 9024 14519 9027
rect 15010 9024 15016 9036
rect 14507 8996 15016 9024
rect 14507 8993 14519 8996
rect 14461 8987 14519 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 15841 9027 15899 9033
rect 15841 9024 15853 9027
rect 15252 8996 15853 9024
rect 15252 8984 15258 8996
rect 15841 8993 15853 8996
rect 15887 8993 15899 9027
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 15841 8987 15899 8993
rect 15948 8996 16405 9024
rect 14553 8959 14611 8965
rect 14553 8956 14565 8959
rect 14108 8928 14565 8956
rect 14553 8925 14565 8928
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 14826 8916 14832 8968
rect 14884 8956 14890 8968
rect 15948 8956 15976 8996
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 17032 9024 17060 9064
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 19521 9095 19579 9101
rect 19521 9061 19533 9095
rect 19567 9092 19579 9095
rect 20530 9092 20536 9104
rect 19567 9064 20536 9092
rect 19567 9061 19579 9064
rect 19521 9055 19579 9061
rect 20530 9052 20536 9064
rect 20588 9052 20594 9104
rect 16393 8987 16451 8993
rect 16500 8996 17060 9024
rect 14884 8928 15976 8956
rect 16025 8959 16083 8965
rect 14884 8916 14890 8928
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 16500 8956 16528 8996
rect 18506 8984 18512 9036
rect 18564 9024 18570 9036
rect 19242 9024 19248 9036
rect 18564 8996 19248 9024
rect 18564 8984 18570 8996
rect 19242 8984 19248 8996
rect 19300 9024 19306 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19300 8996 19625 9024
rect 19300 8984 19306 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 9024 20407 9027
rect 20622 9024 20628 9036
rect 20395 8996 20628 9024
rect 20395 8993 20407 8996
rect 20349 8987 20407 8993
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 16071 8928 16528 8956
rect 16669 8959 16727 8965
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 16669 8925 16681 8959
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 6638 8888 6644 8900
rect 4764 8860 6644 8888
rect 4764 8848 4770 8860
rect 6638 8848 6644 8860
rect 6696 8888 6702 8900
rect 7926 8888 7932 8900
rect 6696 8860 7932 8888
rect 6696 8848 6702 8860
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 12820 8888 12848 8916
rect 15470 8888 15476 8900
rect 12820 8860 15476 8888
rect 15470 8848 15476 8860
rect 15528 8848 15534 8900
rect 15654 8848 15660 8900
rect 15712 8888 15718 8900
rect 16209 8891 16267 8897
rect 16209 8888 16221 8891
rect 15712 8860 16221 8888
rect 15712 8848 15718 8860
rect 16209 8857 16221 8860
rect 16255 8888 16267 8891
rect 16684 8888 16712 8919
rect 17770 8916 17776 8968
rect 17828 8956 17834 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 17828 8928 18613 8956
rect 17828 8916 17834 8928
rect 18601 8925 18613 8928
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8956 18751 8959
rect 19334 8956 19340 8968
rect 18739 8928 19340 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 19334 8916 19340 8928
rect 19392 8956 19398 8968
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19392 8928 19717 8956
rect 19392 8916 19398 8928
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19720 8888 19748 8919
rect 19978 8916 19984 8968
rect 20036 8956 20042 8968
rect 20441 8959 20499 8965
rect 20441 8956 20453 8959
rect 20036 8928 20453 8956
rect 20036 8916 20042 8928
rect 20441 8925 20453 8928
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8925 20591 8959
rect 20533 8919 20591 8925
rect 20254 8888 20260 8900
rect 16255 8860 16712 8888
rect 17604 8860 18644 8888
rect 19720 8860 20260 8888
rect 16255 8857 16267 8860
rect 16209 8851 16267 8857
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 6822 8820 6828 8832
rect 3476 8792 6828 8820
rect 3476 8780 3482 8792
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 8110 8820 8116 8832
rect 7064 8792 8116 8820
rect 7064 8780 7070 8792
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 10870 8820 10876 8832
rect 8720 8792 10876 8820
rect 8720 8780 8726 8792
rect 10870 8780 10876 8792
rect 10928 8820 10934 8832
rect 12802 8820 12808 8832
rect 10928 8792 12808 8820
rect 10928 8780 10934 8792
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 12986 8780 12992 8832
rect 13044 8820 13050 8832
rect 13081 8823 13139 8829
rect 13081 8820 13093 8823
rect 13044 8792 13093 8820
rect 13044 8780 13050 8792
rect 13081 8789 13093 8792
rect 13127 8789 13139 8823
rect 13081 8783 13139 8789
rect 13173 8823 13231 8829
rect 13173 8789 13185 8823
rect 13219 8820 13231 8823
rect 13722 8820 13728 8832
rect 13219 8792 13728 8820
rect 13219 8789 13231 8792
rect 13173 8783 13231 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14001 8823 14059 8829
rect 14001 8820 14013 8823
rect 13872 8792 14013 8820
rect 13872 8780 13878 8792
rect 14001 8789 14013 8792
rect 14047 8789 14059 8823
rect 14001 8783 14059 8789
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 17604 8820 17632 8860
rect 18616 8832 18644 8860
rect 20254 8848 20260 8860
rect 20312 8888 20318 8900
rect 20548 8888 20576 8919
rect 20312 8860 20576 8888
rect 20312 8848 20318 8860
rect 14516 8792 17632 8820
rect 18141 8823 18199 8829
rect 14516 8780 14522 8792
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18506 8820 18512 8832
rect 18187 8792 18512 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 18598 8780 18604 8832
rect 18656 8780 18662 8832
rect 19150 8820 19156 8832
rect 19111 8792 19156 8820
rect 19150 8780 19156 8792
rect 19208 8780 19214 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 2866 8616 2872 8628
rect 1719 8588 2872 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7653 8619 7711 8625
rect 7653 8616 7665 8619
rect 7340 8588 7665 8616
rect 7340 8576 7346 8588
rect 7653 8585 7665 8588
rect 7699 8585 7711 8619
rect 7653 8579 7711 8585
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 10502 8616 10508 8628
rect 7984 8588 10508 8616
rect 7984 8576 7990 8588
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11112 8588 11529 8616
rect 11112 8576 11118 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 12434 8616 12440 8628
rect 11756 8588 12440 8616
rect 11756 8576 11762 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 14366 8616 14372 8628
rect 12667 8588 14372 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14553 8619 14611 8625
rect 14553 8585 14565 8619
rect 14599 8616 14611 8619
rect 16850 8616 16856 8628
rect 14599 8588 16856 8616
rect 14599 8585 14611 8588
rect 14553 8579 14611 8585
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 16945 8619 17003 8625
rect 16945 8585 16957 8619
rect 16991 8616 17003 8619
rect 17126 8616 17132 8628
rect 16991 8588 17132 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18598 8616 18604 8628
rect 18095 8588 18604 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 20806 8616 20812 8628
rect 18923 8588 20812 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8517 2467 8551
rect 5445 8551 5503 8557
rect 5445 8548 5457 8551
rect 2409 8511 2467 8517
rect 2884 8520 5457 8548
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 1486 8412 1492 8424
rect 1447 8384 1492 8412
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 2424 8412 2452 8511
rect 2884 8489 2912 8520
rect 5445 8517 5457 8520
rect 5491 8517 5503 8551
rect 5445 8511 5503 8517
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 6972 8520 7696 8548
rect 6972 8508 6978 8520
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 2869 8443 2927 8449
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3878 8480 3884 8492
rect 3839 8452 3884 8480
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5592 8452 6009 8480
rect 5592 8440 5598 8452
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6880 8452 7389 8480
rect 6880 8440 6886 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 1903 8384 2452 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 3326 8372 3332 8424
rect 3384 8412 3390 8424
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3384 8384 3709 8412
rect 3384 8372 3390 8384
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 6696 8384 7297 8412
rect 6696 8372 6702 8384
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 3605 8347 3663 8353
rect 3605 8313 3617 8347
rect 3651 8344 3663 8347
rect 3970 8344 3976 8356
rect 3651 8316 3976 8344
rect 3651 8313 3663 8316
rect 3605 8307 3663 8313
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 5813 8347 5871 8353
rect 5813 8313 5825 8347
rect 5859 8344 5871 8347
rect 7193 8347 7251 8353
rect 5859 8316 6868 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 2832 8248 2877 8276
rect 2832 8236 2838 8248
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 3237 8279 3295 8285
rect 3237 8276 3249 8279
rect 3200 8248 3249 8276
rect 3200 8236 3206 8248
rect 3237 8245 3249 8248
rect 3283 8245 3295 8279
rect 3237 8239 3295 8245
rect 3786 8236 3792 8288
rect 3844 8276 3850 8288
rect 5074 8276 5080 8288
rect 3844 8248 5080 8276
rect 3844 8236 3850 8248
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5902 8276 5908 8288
rect 5863 8248 5908 8276
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6840 8285 6868 8316
rect 7193 8313 7205 8347
rect 7239 8344 7251 8347
rect 7466 8344 7472 8356
rect 7239 8316 7472 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 7668 8344 7696 8520
rect 9858 8508 9864 8560
rect 9916 8548 9922 8560
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 9916 8520 10057 8548
rect 9916 8508 9922 8520
rect 10045 8517 10057 8520
rect 10091 8548 10103 8551
rect 10091 8520 10171 8548
rect 10091 8517 10103 8520
rect 10045 8511 10103 8517
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 8168 8452 8217 8480
rect 8168 8440 8174 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 10143 8480 10171 8520
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 12216 8520 13391 8548
rect 12216 8508 12222 8520
rect 10143 8452 10272 8480
rect 8205 8443 8263 8449
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 7800 8384 8677 8412
rect 7800 8372 7806 8384
rect 8665 8381 8677 8384
rect 8711 8412 8723 8415
rect 9674 8412 9680 8424
rect 8711 8384 9680 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10144 8415 10202 8421
rect 10144 8412 10156 8415
rect 10060 8384 10156 8412
rect 8021 8347 8079 8353
rect 8021 8344 8033 8347
rect 7668 8316 8033 8344
rect 8021 8313 8033 8316
rect 8067 8313 8079 8347
rect 8021 8307 8079 8313
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8344 8171 8347
rect 8570 8344 8576 8356
rect 8159 8316 8576 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 8932 8347 8990 8353
rect 8932 8313 8944 8347
rect 8978 8344 8990 8347
rect 9582 8344 9588 8356
rect 8978 8316 9588 8344
rect 8978 8313 8990 8316
rect 8932 8307 8990 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 9692 8344 9720 8372
rect 10060 8344 10088 8384
rect 10144 8381 10156 8384
rect 10190 8381 10202 8415
rect 10244 8412 10272 8452
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 12986 8480 12992 8492
rect 11204 8452 12992 8480
rect 11204 8440 11210 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13262 8480 13268 8492
rect 13223 8452 13268 8480
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13363 8480 13391 8520
rect 13446 8508 13452 8560
rect 13504 8548 13510 8560
rect 13725 8551 13783 8557
rect 13725 8548 13737 8551
rect 13504 8520 13737 8548
rect 13504 8508 13510 8520
rect 13725 8517 13737 8520
rect 13771 8548 13783 8551
rect 14734 8548 14740 8560
rect 13771 8520 14740 8548
rect 13771 8517 13783 8520
rect 13725 8511 13783 8517
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 15838 8548 15844 8560
rect 14844 8520 15844 8548
rect 14844 8480 14872 8520
rect 15838 8508 15844 8520
rect 15896 8508 15902 8560
rect 16117 8551 16175 8557
rect 16117 8517 16129 8551
rect 16163 8548 16175 8551
rect 16163 8520 17356 8548
rect 16163 8517 16175 8520
rect 16117 8511 16175 8517
rect 15102 8480 15108 8492
rect 13363 8452 14872 8480
rect 15063 8452 15108 8480
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 16390 8440 16396 8492
rect 16448 8480 16454 8492
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16448 8452 16681 8480
rect 16448 8440 16454 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 10393 8415 10451 8421
rect 10393 8412 10405 8415
rect 10244 8384 10405 8412
rect 10144 8375 10202 8381
rect 10393 8381 10405 8384
rect 10439 8381 10451 8415
rect 10393 8375 10451 8381
rect 13081 8415 13139 8421
rect 13081 8381 13093 8415
rect 13127 8412 13139 8415
rect 13722 8412 13728 8424
rect 13127 8384 13728 8412
rect 13127 8381 13139 8384
rect 13081 8375 13139 8381
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 13906 8412 13912 8424
rect 13867 8384 13912 8412
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 14366 8372 14372 8424
rect 14424 8412 14430 8424
rect 17328 8421 17356 8520
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 20257 8551 20315 8557
rect 20257 8548 20269 8551
rect 17736 8520 18736 8548
rect 17736 8508 17742 8520
rect 17402 8440 17408 8492
rect 17460 8480 17466 8492
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 17460 8452 17509 8480
rect 17460 8440 17466 8452
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18598 8480 18604 8492
rect 18012 8452 18604 8480
rect 18012 8440 18018 8452
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 18708 8480 18736 8520
rect 18892 8520 20269 8548
rect 18892 8480 18920 8520
rect 20257 8517 20269 8520
rect 20303 8517 20315 8551
rect 20257 8511 20315 8517
rect 18708 8452 18920 8480
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 19702 8480 19708 8492
rect 19567 8452 19708 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19852 8452 19901 8480
rect 19852 8440 19858 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 19889 8443 19947 8449
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20220 8452 20821 8480
rect 20220 8440 20226 8452
rect 20809 8449 20821 8452
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 14424 8384 16589 8412
rect 14424 8372 14430 8384
rect 16577 8381 16589 8384
rect 16623 8381 16635 8415
rect 16577 8375 16635 8381
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 18417 8415 18475 8421
rect 17828 8384 18368 8412
rect 17828 8372 17834 8384
rect 9692 8316 10088 8344
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 14458 8344 14464 8356
rect 10560 8316 14464 8344
rect 10560 8304 10566 8316
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 14550 8304 14556 8356
rect 14608 8344 14614 8356
rect 14921 8347 14979 8353
rect 14921 8344 14933 8347
rect 14608 8316 14933 8344
rect 14608 8304 14614 8316
rect 14921 8313 14933 8316
rect 14967 8313 14979 8347
rect 14921 8307 14979 8313
rect 16485 8347 16543 8353
rect 16485 8313 16497 8347
rect 16531 8344 16543 8347
rect 17034 8344 17040 8356
rect 16531 8316 17040 8344
rect 16531 8313 16543 8316
rect 16485 8307 16543 8313
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 6825 8279 6883 8285
rect 6825 8245 6837 8279
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 7558 8236 7564 8288
rect 7616 8276 7622 8288
rect 8386 8276 8392 8288
rect 7616 8248 8392 8276
rect 7616 8236 7622 8248
rect 8386 8236 8392 8248
rect 8444 8276 8450 8288
rect 9674 8276 9680 8288
rect 8444 8248 9680 8276
rect 8444 8236 8450 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 11606 8236 11612 8288
rect 11664 8276 11670 8288
rect 11664 8248 11709 8276
rect 11664 8236 11670 8248
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 12989 8279 13047 8285
rect 12989 8276 13001 8279
rect 12860 8248 13001 8276
rect 12860 8236 12866 8248
rect 12989 8245 13001 8248
rect 13035 8245 13047 8279
rect 12989 8239 13047 8245
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14274 8276 14280 8288
rect 13872 8248 14280 8276
rect 13872 8236 13878 8248
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 15068 8248 15113 8276
rect 15068 8236 15074 8248
rect 15378 8236 15384 8288
rect 15436 8276 15442 8288
rect 15746 8276 15752 8288
rect 15436 8248 15752 8276
rect 15436 8236 15442 8248
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 18340 8276 18368 8384
rect 18417 8381 18429 8415
rect 18463 8412 18475 8415
rect 18506 8412 18512 8424
rect 18463 8384 18512 8412
rect 18463 8381 18475 8384
rect 18417 8375 18475 8381
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 19334 8412 19340 8424
rect 19295 8384 19340 8412
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 20717 8415 20775 8421
rect 20717 8412 20729 8415
rect 20680 8384 20729 8412
rect 20680 8372 20686 8384
rect 20717 8381 20729 8384
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 19245 8347 19303 8353
rect 19245 8313 19257 8347
rect 19291 8344 19303 8347
rect 19886 8344 19892 8356
rect 19291 8316 19892 8344
rect 19291 8313 19303 8316
rect 19245 8307 19303 8313
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 20588 8316 20668 8344
rect 20588 8304 20594 8316
rect 20640 8285 20668 8316
rect 18509 8279 18567 8285
rect 18509 8276 18521 8279
rect 18340 8248 18521 8276
rect 18509 8245 18521 8248
rect 18555 8245 18567 8279
rect 18509 8239 18567 8245
rect 20625 8279 20683 8285
rect 20625 8245 20637 8279
rect 20671 8245 20683 8279
rect 20625 8239 20683 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 3050 8072 3056 8084
rect 3007 8044 3056 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3602 8072 3608 8084
rect 3559 8044 3608 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 3602 8032 3608 8044
rect 3660 8072 3666 8084
rect 3786 8072 3792 8084
rect 3660 8044 3792 8072
rect 3660 8032 3666 8044
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 5960 8044 6285 8072
rect 5960 8032 5966 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 6687 8044 7113 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 7101 8035 7159 8041
rect 7469 8075 7527 8081
rect 7469 8041 7481 8075
rect 7515 8072 7527 8075
rect 7558 8072 7564 8084
rect 7515 8044 7564 8072
rect 7515 8041 7527 8044
rect 7469 8035 7527 8041
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8435 8044 8769 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8757 8041 8769 8044
rect 8803 8041 8815 8075
rect 8757 8035 8815 8041
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 9677 8075 9735 8081
rect 8996 8044 9628 8072
rect 8996 8032 9002 8044
rect 3878 8004 3884 8016
rect 3791 7976 3884 8004
rect 1848 7939 1906 7945
rect 1848 7905 1860 7939
rect 1894 7936 1906 7939
rect 3418 7936 3424 7948
rect 1894 7908 3424 7936
rect 1894 7905 1906 7908
rect 1848 7899 1906 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 3804 7877 3832 7976
rect 3878 7964 3884 7976
rect 3936 8004 3942 8016
rect 4424 8007 4482 8013
rect 4424 8004 4436 8007
rect 3936 7976 4436 8004
rect 3936 7964 3942 7976
rect 4424 7973 4436 7976
rect 4470 8004 4482 8007
rect 6822 8004 6828 8016
rect 4470 7976 6828 8004
rect 4470 7973 4482 7976
rect 4424 7967 4482 7973
rect 6822 7964 6828 7976
rect 6880 8004 6886 8016
rect 8297 8007 8355 8013
rect 6880 7976 6960 8004
rect 6880 7964 6886 7976
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4157 7939 4215 7945
rect 4157 7936 4169 7939
rect 4120 7908 4169 7936
rect 4120 7896 4126 7908
rect 4157 7905 4169 7908
rect 4203 7936 4215 7939
rect 4246 7936 4252 7948
rect 4203 7908 4252 7936
rect 4203 7905 4215 7908
rect 4157 7899 4215 7905
rect 4246 7896 4252 7908
rect 4304 7936 4310 7948
rect 5905 7939 5963 7945
rect 4304 7908 5212 7936
rect 4304 7896 4310 7908
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 5184 7800 5212 7908
rect 5905 7905 5917 7939
rect 5951 7936 5963 7939
rect 6270 7936 6276 7948
rect 5951 7908 6276 7936
rect 5951 7905 5963 7908
rect 5905 7899 5963 7905
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6932 7877 6960 7976
rect 8297 7973 8309 8007
rect 8343 8004 8355 8007
rect 9490 8004 9496 8016
rect 8343 7976 9496 8004
rect 8343 7973 8355 7976
rect 8297 7967 8355 7973
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 9600 8004 9628 8044
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 9950 8072 9956 8084
rect 9723 8044 9956 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11606 8072 11612 8084
rect 10919 8044 11612 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 14090 8072 14096 8084
rect 11716 8044 14096 8072
rect 9766 8004 9772 8016
rect 9600 7976 9772 8004
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10502 7964 10508 8016
rect 10560 8004 10566 8016
rect 11716 8004 11744 8044
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14366 8072 14372 8084
rect 14327 8044 14372 8072
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 15378 8072 15384 8084
rect 14516 8044 15384 8072
rect 14516 8032 14522 8044
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 17402 8072 17408 8084
rect 16807 8044 17408 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 18509 8075 18567 8081
rect 18509 8041 18521 8075
rect 18555 8072 18567 8075
rect 19150 8072 19156 8084
rect 18555 8044 19156 8072
rect 18555 8041 18567 8044
rect 18509 8035 18567 8041
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 20312 8044 20545 8072
rect 20312 8032 20318 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 20533 8035 20591 8041
rect 10560 7976 11744 8004
rect 12796 8007 12854 8013
rect 10560 7964 10566 7976
rect 12796 7973 12808 8007
rect 12842 8004 12854 8007
rect 12986 8004 12992 8016
rect 12842 7976 12992 8004
rect 12842 7973 12854 7976
rect 12796 7967 12854 7973
rect 12986 7964 12992 7976
rect 13044 7964 13050 8016
rect 13078 7964 13084 8016
rect 13136 8004 13142 8016
rect 13722 8004 13728 8016
rect 13136 7976 13728 8004
rect 13136 7964 13142 7976
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 17129 8007 17187 8013
rect 17129 7973 17141 8007
rect 17175 8004 17187 8007
rect 17678 8004 17684 8016
rect 17175 7976 17684 8004
rect 17175 7973 17187 7976
rect 17129 7967 17187 7973
rect 17678 7964 17684 7976
rect 17736 7964 17742 8016
rect 18417 8007 18475 8013
rect 18417 7973 18429 8007
rect 18463 8004 18475 8007
rect 18690 8004 18696 8016
rect 18463 7976 18696 8004
rect 18463 7973 18475 7976
rect 18417 7967 18475 7973
rect 18690 7964 18696 7976
rect 18748 7964 18754 8016
rect 19426 8013 19432 8016
rect 19420 8004 19432 8013
rect 19387 7976 19432 8004
rect 19420 7967 19432 7976
rect 19426 7964 19432 7967
rect 19484 7964 19490 8016
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 7616 7908 7661 7936
rect 7616 7896 7622 7908
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 9125 7939 9183 7945
rect 9125 7936 9137 7939
rect 8444 7908 9137 7936
rect 8444 7896 8450 7908
rect 9125 7905 9137 7908
rect 9171 7905 9183 7939
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9125 7899 9183 7905
rect 9324 7908 10057 7936
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7868 7803 7871
rect 7834 7868 7840 7880
rect 7791 7840 7840 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 5721 7803 5779 7809
rect 5721 7800 5733 7803
rect 5184 7772 5733 7800
rect 5721 7769 5733 7772
rect 5767 7769 5779 7803
rect 5721 7763 5779 7769
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 6178 7800 6184 7812
rect 5960 7772 6184 7800
rect 5960 7760 5966 7772
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6748 7800 6776 7831
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 7190 7800 7196 7812
rect 6748 7772 7196 7800
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 8588 7800 8616 7831
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 8812 7840 9229 7868
rect 8812 7828 8818 7840
rect 9217 7837 9229 7840
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 8938 7800 8944 7812
rect 7852 7772 8524 7800
rect 8588 7772 8944 7800
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 3234 7732 3240 7744
rect 3191 7704 3240 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 7852 7732 7880 7772
rect 4120 7704 7880 7732
rect 7929 7735 7987 7741
rect 4120 7692 4126 7704
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8294 7732 8300 7744
rect 7975 7704 8300 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8496 7732 8524 7772
rect 8938 7760 8944 7772
rect 8996 7760 9002 7812
rect 9324 7732 9352 7908
rect 10045 7905 10057 7908
rect 10091 7936 10103 7939
rect 10686 7936 10692 7948
rect 10091 7908 10692 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10962 7936 10968 7948
rect 10875 7908 10968 7936
rect 10962 7896 10968 7908
rect 11020 7936 11026 7948
rect 12250 7936 12256 7948
rect 11020 7908 12256 7936
rect 11020 7896 11026 7908
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 14056 7908 14749 7936
rect 14056 7896 14062 7908
rect 14737 7905 14749 7908
rect 14783 7905 14795 7939
rect 15102 7936 15108 7948
rect 15015 7908 15108 7936
rect 14737 7899 14795 7905
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9858 7868 9864 7880
rect 9447 7840 9864 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10134 7868 10140 7880
rect 10047 7840 10140 7868
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 11057 7871 11115 7877
rect 11057 7868 11069 7871
rect 10321 7831 10379 7837
rect 10888 7840 11069 7868
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 10152 7800 10180 7828
rect 9824 7772 10180 7800
rect 10336 7800 10364 7831
rect 10888 7800 10916 7840
rect 11057 7837 11069 7840
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12492 7840 12541 7868
rect 12492 7828 12498 7840
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 13630 7868 13636 7880
rect 13543 7840 13636 7868
rect 12529 7831 12587 7837
rect 10336 7772 10916 7800
rect 9824 7760 9830 7772
rect 8496 7704 9352 7732
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 10336 7732 10364 7772
rect 11238 7760 11244 7812
rect 11296 7800 11302 7812
rect 11296 7772 12572 7800
rect 11296 7760 11302 7772
rect 9640 7704 10364 7732
rect 10505 7735 10563 7741
rect 9640 7692 9646 7704
rect 10505 7701 10517 7735
rect 10551 7732 10563 7735
rect 10686 7732 10692 7744
rect 10551 7704 10692 7732
rect 10551 7701 10563 7704
rect 10505 7695 10563 7701
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 12342 7732 12348 7744
rect 11112 7704 12348 7732
rect 11112 7692 11118 7704
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 12544 7732 12572 7772
rect 13556 7732 13584 7840
rect 13630 7828 13636 7840
rect 13688 7868 13694 7880
rect 15028 7877 15056 7908
rect 15102 7896 15108 7908
rect 15160 7936 15166 7948
rect 15556 7939 15614 7945
rect 15556 7936 15568 7939
rect 15160 7908 15568 7936
rect 15160 7896 15166 7908
rect 15556 7905 15568 7908
rect 15602 7936 15614 7939
rect 16666 7936 16672 7948
rect 15602 7908 16672 7936
rect 15602 7905 15614 7908
rect 15556 7899 15614 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 16850 7896 16856 7948
rect 16908 7936 16914 7948
rect 17221 7939 17279 7945
rect 17221 7936 17233 7939
rect 16908 7908 17233 7936
rect 16908 7896 16914 7908
rect 17221 7905 17233 7908
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 19153 7939 19211 7945
rect 19153 7936 19165 7939
rect 18564 7908 19165 7936
rect 18564 7896 18570 7908
rect 19153 7905 19165 7908
rect 19199 7905 19211 7939
rect 19153 7899 19211 7905
rect 14829 7871 14887 7877
rect 14829 7868 14841 7871
rect 13688 7840 14841 7868
rect 13688 7828 13694 7840
rect 14829 7837 14841 7840
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 17313 7871 17371 7877
rect 17313 7868 17325 7871
rect 15289 7831 15347 7837
rect 16684 7840 17325 7868
rect 12544 7704 13584 7732
rect 13630 7692 13636 7744
rect 13688 7732 13694 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 13688 7704 13921 7732
rect 13688 7692 13694 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 15304 7732 15332 7831
rect 15654 7732 15660 7744
rect 15304 7704 15660 7732
rect 13909 7695 13967 7701
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 16390 7692 16396 7744
rect 16448 7732 16454 7744
rect 16684 7741 16712 7840
rect 17313 7837 17325 7840
rect 17359 7837 17371 7871
rect 18598 7868 18604 7880
rect 18559 7840 18604 7868
rect 17313 7831 17371 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 18049 7803 18107 7809
rect 18049 7769 18061 7803
rect 18095 7800 18107 7803
rect 18966 7800 18972 7812
rect 18095 7772 18972 7800
rect 18095 7769 18107 7772
rect 18049 7763 18107 7769
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 16669 7735 16727 7741
rect 16669 7732 16681 7735
rect 16448 7704 16681 7732
rect 16448 7692 16454 7704
rect 16669 7701 16681 7704
rect 16715 7701 16727 7735
rect 16669 7695 16727 7701
rect 16758 7692 16764 7744
rect 16816 7732 16822 7744
rect 17678 7732 17684 7744
rect 16816 7704 17684 7732
rect 16816 7692 16822 7704
rect 17678 7692 17684 7704
rect 17736 7732 17742 7744
rect 20162 7732 20168 7744
rect 17736 7704 20168 7732
rect 17736 7692 17742 7704
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 2832 7500 2877 7528
rect 2832 7488 2838 7500
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 3697 7531 3755 7537
rect 3697 7528 3709 7531
rect 3660 7500 3709 7528
rect 3660 7488 3666 7500
rect 3697 7497 3709 7500
rect 3743 7497 3755 7531
rect 3697 7491 3755 7497
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 12342 7528 12348 7540
rect 4120 7500 12348 7528
rect 4120 7488 4126 7500
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 14274 7528 14280 7540
rect 12492 7500 14280 7528
rect 12492 7488 12498 7500
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15470 7528 15476 7540
rect 14783 7500 15476 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 18598 7528 18604 7540
rect 15580 7500 18604 7528
rect 3786 7460 3792 7472
rect 3344 7432 3792 7460
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1544 7364 1593 7392
rect 1544 7352 1550 7364
rect 1581 7361 1593 7364
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2774 7392 2780 7404
rect 2639 7364 2780 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 3234 7392 3240 7404
rect 3195 7364 3240 7392
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7293 1455 7327
rect 3142 7324 3148 7336
rect 3103 7296 3148 7324
rect 1397 7287 1455 7293
rect 1412 7188 1440 7287
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 1949 7191 2007 7197
rect 1949 7188 1961 7191
rect 1412 7160 1961 7188
rect 1949 7157 1961 7160
rect 1995 7157 2007 7191
rect 2314 7188 2320 7200
rect 2275 7160 2320 7188
rect 1949 7151 2007 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 2409 7191 2467 7197
rect 2409 7157 2421 7191
rect 2455 7188 2467 7191
rect 2958 7188 2964 7200
rect 2455 7160 2964 7188
rect 2455 7157 2467 7160
rect 2409 7151 2467 7157
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3344 7188 3372 7432
rect 3786 7420 3792 7432
rect 3844 7420 3850 7472
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 4430 7460 4436 7472
rect 3936 7432 4436 7460
rect 3936 7420 3942 7432
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 4264 7401 4292 7432
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7460 5963 7463
rect 6822 7460 6828 7472
rect 5951 7432 6828 7460
rect 5951 7429 5963 7432
rect 5905 7423 5963 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 7101 7463 7159 7469
rect 7101 7429 7113 7463
rect 7147 7460 7159 7463
rect 7190 7460 7196 7472
rect 7147 7432 7196 7460
rect 7147 7429 7159 7432
rect 7101 7423 7159 7429
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 7742 7420 7748 7472
rect 7800 7460 7806 7472
rect 7929 7463 7987 7469
rect 7929 7460 7941 7463
rect 7800 7432 7941 7460
rect 7800 7420 7806 7432
rect 7929 7429 7941 7432
rect 7975 7429 7987 7463
rect 7929 7423 7987 7429
rect 8110 7420 8116 7472
rect 8168 7420 8174 7472
rect 8386 7460 8392 7472
rect 8347 7432 8392 7460
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10410 7460 10416 7472
rect 10008 7432 10416 7460
rect 10008 7420 10014 7432
rect 10410 7420 10416 7432
rect 10468 7420 10474 7472
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 15580 7460 15608 7500
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 19886 7528 19892 7540
rect 19847 7500 19892 7528
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 17034 7460 17040 7472
rect 12124 7432 15608 7460
rect 16995 7432 17040 7460
rect 12124 7420 12130 7432
rect 17034 7420 17040 7432
rect 17092 7420 17098 7472
rect 19426 7420 19432 7472
rect 19484 7460 19490 7472
rect 19797 7463 19855 7469
rect 19797 7460 19809 7463
rect 19484 7432 19809 7460
rect 19484 7420 19490 7432
rect 19797 7429 19809 7432
rect 19843 7429 19855 7463
rect 19797 7423 19855 7429
rect 4249 7395 4307 7401
rect 3476 7364 3521 7392
rect 3476 7352 3482 7364
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 4396 7364 4537 7392
rect 4396 7352 4402 7364
rect 4525 7361 4537 7364
rect 4571 7361 4583 7395
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 4525 7355 4583 7361
rect 7208 7364 7665 7392
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 3752 7296 4108 7324
rect 3752 7284 3758 7296
rect 4080 7256 4108 7296
rect 7208 7268 7236 7364
rect 7653 7361 7665 7364
rect 7699 7392 7711 7395
rect 7834 7392 7840 7404
rect 7699 7364 7840 7392
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 8128 7392 8156 7420
rect 7944 7364 8156 7392
rect 9033 7395 9091 7401
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7324 7527 7327
rect 7558 7324 7564 7336
rect 7515 7296 7564 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 4157 7259 4215 7265
rect 4157 7256 4169 7259
rect 4080 7228 4169 7256
rect 4157 7225 4169 7228
rect 4203 7225 4215 7259
rect 4157 7219 4215 7225
rect 4430 7216 4436 7268
rect 4488 7256 4494 7268
rect 4770 7259 4828 7265
rect 4770 7256 4782 7259
rect 4488 7228 4782 7256
rect 4488 7216 4494 7228
rect 4770 7225 4782 7228
rect 4816 7256 4828 7259
rect 7190 7256 7196 7268
rect 4816 7228 7196 7256
rect 4816 7225 4828 7228
rect 4770 7219 4828 7225
rect 7190 7216 7196 7228
rect 7248 7216 7254 7268
rect 3292 7160 3372 7188
rect 3292 7148 3298 7160
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 3844 7160 4077 7188
rect 3844 7148 3850 7160
rect 4065 7157 4077 7160
rect 4111 7157 4123 7191
rect 4065 7151 4123 7157
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7484 7188 7512 7287
rect 7558 7284 7564 7296
rect 7616 7324 7622 7336
rect 7944 7324 7972 7364
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9582 7392 9588 7404
rect 9079 7364 9588 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10226 7392 10232 7404
rect 9907 7364 10232 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10226 7352 10232 7364
rect 10284 7392 10290 7404
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10284 7364 10609 7392
rect 10284 7352 10290 7364
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 13630 7392 13636 7404
rect 13591 7364 13636 7392
rect 10597 7355 10655 7361
rect 13630 7352 13636 7364
rect 13688 7392 13694 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 13688 7364 14473 7392
rect 13688 7352 13694 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 15289 7395 15347 7401
rect 15289 7392 15301 7395
rect 14608 7364 15301 7392
rect 14608 7352 14614 7364
rect 15289 7361 15301 7364
rect 15335 7361 15347 7395
rect 17678 7392 17684 7404
rect 15289 7355 15347 7361
rect 15396 7364 15700 7392
rect 17639 7364 17684 7392
rect 7616 7296 7972 7324
rect 8113 7327 8171 7333
rect 7616 7284 7622 7296
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8202 7324 8208 7336
rect 8159 7296 8208 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 10502 7324 10508 7336
rect 10463 7296 10508 7324
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 12434 7324 12440 7336
rect 10919 7296 12440 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11348 7268 11376 7296
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7324 12679 7327
rect 13446 7324 13452 7336
rect 12667 7296 13452 7324
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7324 13599 7327
rect 13814 7324 13820 7336
rect 13587 7296 13820 7324
rect 13587 7293 13599 7296
rect 13541 7287 13599 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 13964 7296 14381 7324
rect 13964 7284 13970 7296
rect 14369 7293 14381 7296
rect 14415 7324 14427 7327
rect 15396 7324 15424 7364
rect 14415 7296 15424 7324
rect 15565 7327 15623 7333
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 15565 7293 15577 7327
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 7926 7256 7932 7268
rect 7576 7228 7932 7256
rect 7576 7197 7604 7228
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 8938 7256 8944 7268
rect 8027 7228 8944 7256
rect 7055 7160 7512 7188
rect 7561 7191 7619 7197
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7561 7157 7573 7191
rect 7607 7157 7619 7191
rect 7561 7151 7619 7157
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 8027 7188 8055 7228
rect 8938 7216 8944 7228
rect 8996 7216 9002 7268
rect 10413 7259 10471 7265
rect 9692 7228 10364 7256
rect 7708 7160 8055 7188
rect 7708 7148 7714 7160
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 8757 7191 8815 7197
rect 8757 7188 8769 7191
rect 8720 7160 8769 7188
rect 8720 7148 8726 7160
rect 8757 7157 8769 7160
rect 8803 7157 8815 7191
rect 8757 7151 8815 7157
rect 8849 7191 8907 7197
rect 8849 7157 8861 7191
rect 8895 7188 8907 7191
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8895 7160 9229 7188
rect 8895 7157 8907 7160
rect 8849 7151 8907 7157
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 9217 7151 9275 7157
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 9692 7197 9720 7228
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 9548 7160 9597 7188
rect 9548 7148 9554 7160
rect 9585 7157 9597 7160
rect 9631 7157 9643 7191
rect 9585 7151 9643 7157
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7157 9735 7191
rect 9677 7151 9735 7157
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 9824 7160 10057 7188
rect 9824 7148 9830 7160
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 10336 7188 10364 7228
rect 10413 7225 10425 7259
rect 10459 7256 10471 7259
rect 10594 7256 10600 7268
rect 10459 7228 10600 7256
rect 10459 7225 10471 7228
rect 10413 7219 10471 7225
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 11146 7265 11152 7268
rect 11140 7256 11152 7265
rect 11107 7228 11152 7256
rect 11140 7219 11152 7228
rect 11146 7216 11152 7219
rect 11204 7216 11210 7268
rect 11330 7216 11336 7268
rect 11388 7216 11394 7268
rect 11514 7216 11520 7268
rect 11572 7256 11578 7268
rect 12713 7259 12771 7265
rect 11572 7228 12296 7256
rect 11572 7216 11578 7228
rect 12158 7188 12164 7200
rect 10336 7160 12164 7188
rect 10045 7151 10103 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12268 7197 12296 7228
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 14277 7259 14335 7265
rect 14277 7256 14289 7259
rect 12759 7228 14289 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 14277 7225 14289 7228
rect 14323 7225 14335 7259
rect 14277 7219 14335 7225
rect 15010 7216 15016 7268
rect 15068 7256 15074 7268
rect 15105 7259 15163 7265
rect 15105 7256 15117 7259
rect 15068 7228 15117 7256
rect 15068 7216 15074 7228
rect 15105 7225 15117 7228
rect 15151 7225 15163 7259
rect 15105 7219 15163 7225
rect 15197 7259 15255 7265
rect 15197 7225 15209 7259
rect 15243 7256 15255 7259
rect 15378 7256 15384 7268
rect 15243 7228 15384 7256
rect 15243 7225 15255 7228
rect 15197 7219 15255 7225
rect 15378 7216 15384 7228
rect 15436 7216 15442 7268
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12342 7188 12348 7200
rect 12299 7160 12348 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13081 7191 13139 7197
rect 13081 7188 13093 7191
rect 12952 7160 13093 7188
rect 12952 7148 12958 7160
rect 13081 7157 13093 7160
rect 13127 7157 13139 7191
rect 13446 7188 13452 7200
rect 13407 7160 13452 7188
rect 13081 7151 13139 7157
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13906 7188 13912 7200
rect 13867 7160 13912 7188
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 15580 7188 15608 7287
rect 15672 7256 15700 7364
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 20438 7392 20444 7404
rect 20399 7364 20444 7392
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 15832 7327 15890 7333
rect 15832 7293 15844 7327
rect 15878 7324 15890 7327
rect 16390 7324 16396 7336
rect 15878 7296 16396 7324
rect 15878 7293 15890 7296
rect 15832 7287 15890 7293
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 17497 7327 17555 7333
rect 17497 7324 17509 7327
rect 16500 7296 17509 7324
rect 15930 7256 15936 7268
rect 15672 7228 15936 7256
rect 15930 7216 15936 7228
rect 15988 7256 15994 7268
rect 16500 7256 16528 7296
rect 17497 7293 17509 7296
rect 17543 7293 17555 7327
rect 17497 7287 17555 7293
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18506 7324 18512 7336
rect 18463 7296 18512 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 18684 7327 18742 7333
rect 18684 7293 18696 7327
rect 18730 7324 18742 7327
rect 19702 7324 19708 7336
rect 18730 7296 19708 7324
rect 18730 7293 18742 7296
rect 18684 7287 18742 7293
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 17405 7259 17463 7265
rect 15988 7228 16528 7256
rect 16684 7228 17356 7256
rect 15988 7216 15994 7228
rect 14516 7160 15608 7188
rect 14516 7148 14522 7160
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16684 7188 16712 7228
rect 15804 7160 16712 7188
rect 16945 7191 17003 7197
rect 15804 7148 15810 7160
rect 16945 7157 16957 7191
rect 16991 7188 17003 7191
rect 17218 7188 17224 7200
rect 16991 7160 17224 7188
rect 16991 7157 17003 7160
rect 16945 7151 17003 7157
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 17328 7188 17356 7228
rect 17405 7225 17417 7259
rect 17451 7256 17463 7259
rect 18049 7259 18107 7265
rect 18049 7256 18061 7259
rect 17451 7228 18061 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 18049 7225 18061 7228
rect 18095 7225 18107 7259
rect 18049 7219 18107 7225
rect 18874 7216 18880 7268
rect 18932 7256 18938 7268
rect 20349 7259 20407 7265
rect 20349 7256 20361 7259
rect 18932 7228 20361 7256
rect 18932 7216 18938 7228
rect 20349 7225 20361 7228
rect 20395 7225 20407 7259
rect 20349 7219 20407 7225
rect 18138 7188 18144 7200
rect 17328 7160 18144 7188
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 19242 7188 19248 7200
rect 18656 7160 19248 7188
rect 18656 7148 18662 7160
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 19518 7148 19524 7200
rect 19576 7188 19582 7200
rect 19794 7188 19800 7200
rect 19576 7160 19800 7188
rect 19576 7148 19582 7160
rect 19794 7148 19800 7160
rect 19852 7148 19858 7200
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 2314 6984 2320 6996
rect 1719 6956 2320 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 3878 6984 3884 6996
rect 3839 6956 3884 6984
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 7006 6984 7012 6996
rect 4948 6956 7012 6984
rect 4948 6944 4954 6956
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 8478 6984 8484 6996
rect 7147 6956 8484 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 8754 6984 8760 6996
rect 8715 6956 8760 6984
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 9125 6987 9183 6993
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9677 6987 9735 6993
rect 9677 6984 9689 6987
rect 9171 6956 9689 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9677 6953 9689 6956
rect 9723 6953 9735 6987
rect 9677 6947 9735 6953
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 11054 6984 11060 6996
rect 10091 6956 11060 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 11204 6956 12664 6984
rect 11204 6944 11210 6956
rect 2038 6916 2044 6928
rect 1999 6888 2044 6916
rect 2038 6876 2044 6888
rect 2096 6876 2102 6928
rect 3602 6916 3608 6928
rect 2516 6888 3608 6916
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 2516 6857 2544 6888
rect 3602 6876 3608 6888
rect 3660 6916 3666 6928
rect 3660 6888 4384 6916
rect 3660 6876 3666 6888
rect 4356 6860 4384 6888
rect 4982 6876 4988 6928
rect 5040 6916 5046 6928
rect 5166 6916 5172 6928
rect 5040 6888 5172 6916
rect 5040 6876 5046 6888
rect 5166 6876 5172 6888
rect 5224 6876 5230 6928
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 7248 6888 7972 6916
rect 7248 6876 7254 6888
rect 2774 6857 2780 6860
rect 2501 6851 2559 6857
rect 2501 6848 2513 6851
rect 1636 6820 2513 6848
rect 1636 6808 1642 6820
rect 2501 6817 2513 6820
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 2768 6811 2780 6857
rect 2832 6848 2838 6860
rect 2832 6820 2868 6848
rect 2774 6808 2780 6811
rect 2832 6808 2838 6820
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 4028 6820 4077 6848
rect 4028 6808 4034 6820
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 4396 6820 4813 6848
rect 4396 6808 4402 6820
rect 4801 6817 4813 6820
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 5068 6851 5126 6857
rect 5068 6817 5080 6851
rect 5114 6848 5126 6851
rect 5994 6848 6000 6860
rect 5114 6820 6000 6848
rect 5114 6817 5126 6820
rect 5068 6811 5126 6817
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6748 6820 7021 6848
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2363 6752 2544 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2516 6644 2544 6752
rect 6638 6712 6644 6724
rect 6599 6684 6644 6712
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 6748 6656 6776 6820
rect 7009 6817 7021 6820
rect 7055 6848 7067 6851
rect 7650 6848 7656 6860
rect 7055 6820 7656 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 7834 6848 7840 6860
rect 7795 6820 7840 6848
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 7944 6848 7972 6888
rect 8018 6876 8024 6928
rect 8076 6916 8082 6928
rect 8938 6916 8944 6928
rect 8076 6888 8944 6916
rect 8076 6876 8082 6888
rect 8938 6876 8944 6888
rect 8996 6916 9002 6928
rect 9306 6916 9312 6928
rect 8996 6888 9312 6916
rect 8996 6876 9002 6888
rect 9306 6876 9312 6888
rect 9364 6876 9370 6928
rect 10134 6916 10140 6928
rect 10047 6888 10140 6916
rect 10134 6876 10140 6888
rect 10192 6916 10198 6928
rect 10502 6916 10508 6928
rect 10192 6888 10508 6916
rect 10192 6876 10198 6888
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 10962 6876 10968 6928
rect 11020 6876 11026 6928
rect 11514 6876 11520 6928
rect 11572 6925 11578 6928
rect 11572 6919 11636 6925
rect 11572 6885 11590 6919
rect 11624 6885 11636 6919
rect 12636 6916 12664 6956
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12768 6956 12909 6984
rect 12768 6944 12774 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13044 6956 13737 6984
rect 13044 6944 13050 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 13725 6947 13783 6953
rect 14660 6956 15669 6984
rect 14660 6928 14688 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 15657 6947 15715 6953
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 19150 6984 19156 6996
rect 15896 6956 19156 6984
rect 15896 6944 15902 6956
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 19702 6984 19708 6996
rect 19663 6956 19708 6984
rect 19702 6944 19708 6956
rect 19760 6944 19766 6996
rect 19797 6987 19855 6993
rect 19797 6953 19809 6987
rect 19843 6984 19855 6987
rect 20254 6984 20260 6996
rect 19843 6956 20260 6984
rect 19843 6953 19855 6956
rect 19797 6947 19855 6953
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 13630 6916 13636 6928
rect 12636 6888 13636 6916
rect 11572 6879 11636 6885
rect 11572 6876 11578 6879
rect 9217 6851 9275 6857
rect 7944 6820 8064 6848
rect 7190 6780 7196 6792
rect 7151 6752 7196 6780
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7926 6780 7932 6792
rect 7300 6752 7932 6780
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 7300 6712 7328 6752
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 8036 6789 8064 6820
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9766 6848 9772 6860
rect 9263 6820 9772 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10980 6848 11008 6876
rect 10008 6820 11008 6848
rect 10008 6808 10014 6820
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 13262 6848 13268 6860
rect 11112 6820 12388 6848
rect 13223 6820 13268 6848
rect 11112 6808 11118 6820
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9582 6780 9588 6792
rect 9447 6752 9588 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10284 6752 10329 6780
rect 10284 6740 10290 6752
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11330 6780 11336 6792
rect 11020 6752 11336 6780
rect 11020 6740 11026 6752
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 7466 6712 7472 6724
rect 7064 6684 7328 6712
rect 7427 6684 7472 6712
rect 7064 6672 7070 6684
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 7558 6672 7564 6724
rect 7616 6712 7622 6724
rect 12360 6712 12388 6820
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 13464 6789 13492 6888
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 14090 6916 14096 6928
rect 14051 6888 14096 6916
rect 14090 6876 14096 6888
rect 14148 6876 14154 6928
rect 14642 6876 14648 6928
rect 14700 6876 14706 6928
rect 15102 6876 15108 6928
rect 15160 6916 15166 6928
rect 16390 6916 16396 6928
rect 15160 6888 16396 6916
rect 15160 6876 15166 6888
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 17405 6919 17463 6925
rect 17405 6885 17417 6919
rect 17451 6916 17463 6919
rect 17954 6916 17960 6928
rect 17451 6888 17960 6916
rect 17451 6885 17463 6888
rect 17405 6879 17463 6885
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 18138 6876 18144 6928
rect 18196 6916 18202 6928
rect 18196 6888 19748 6916
rect 18196 6876 18202 6888
rect 15120 6848 15148 6876
rect 19720 6860 19748 6888
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 13648 6820 15148 6848
rect 15764 6820 16129 6848
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 13372 6712 13400 6743
rect 13648 6712 13676 6820
rect 15764 6792 15792 6820
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18325 6851 18383 6857
rect 18325 6848 18337 6851
rect 17920 6820 18337 6848
rect 17920 6808 17926 6820
rect 18325 6817 18337 6820
rect 18371 6848 18383 6851
rect 18414 6848 18420 6860
rect 18371 6820 18420 6848
rect 18371 6817 18383 6820
rect 18325 6811 18383 6817
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18592 6851 18650 6857
rect 18592 6817 18604 6851
rect 18638 6848 18650 6851
rect 19426 6848 19432 6860
rect 18638 6820 19432 6848
rect 18638 6817 18650 6820
rect 18592 6811 18650 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 19702 6808 19708 6860
rect 19760 6808 19766 6860
rect 20162 6848 20168 6860
rect 20123 6820 20168 6848
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 14182 6780 14188 6792
rect 14143 6752 14188 6780
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6780 14427 6783
rect 14918 6780 14924 6792
rect 14415 6752 14924 6780
rect 14415 6749 14427 6752
rect 14369 6743 14427 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15746 6780 15752 6792
rect 15707 6752 15752 6780
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 17727 6752 18276 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 7616 6684 11183 6712
rect 12360 6684 13676 6712
rect 7616 6672 7622 6684
rect 2866 6644 2872 6656
rect 2516 6616 2872 6644
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 6178 6644 6184 6656
rect 6139 6616 6184 6644
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 6730 6644 6736 6656
rect 6595 6616 6736 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 9950 6644 9956 6656
rect 8536 6616 9956 6644
rect 8536 6604 8542 6616
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10502 6644 10508 6656
rect 10463 6616 10508 6644
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 11155 6644 11183 6684
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 15010 6712 15016 6724
rect 13872 6684 15016 6712
rect 13872 6672 13878 6684
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 15289 6715 15347 6721
rect 15289 6681 15301 6715
rect 15335 6712 15347 6715
rect 17512 6712 17540 6743
rect 15335 6684 17540 6712
rect 15335 6681 15347 6684
rect 15289 6675 15347 6681
rect 12434 6644 12440 6656
rect 11155 6616 12440 6644
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 12526 6604 12532 6656
rect 12584 6644 12590 6656
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12584 6616 12725 6644
rect 12584 6604 12590 6616
rect 12713 6613 12725 6616
rect 12759 6644 12771 6647
rect 14550 6644 14556 6656
rect 12759 6616 14556 6644
rect 12759 6613 12771 6616
rect 12713 6607 12771 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 17034 6644 17040 6656
rect 16995 6616 17040 6644
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 18248 6644 18276 6752
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 19576 6752 20269 6780
rect 19576 6740 19582 6752
rect 20257 6749 20269 6752
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 19242 6644 19248 6656
rect 18248 6616 19248 6644
rect 19242 6604 19248 6616
rect 19300 6644 19306 6656
rect 20364 6644 20392 6743
rect 19300 6616 20392 6644
rect 19300 6604 19306 6616
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2958 6440 2964 6452
rect 2919 6412 2964 6440
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 6270 6440 6276 6452
rect 4028 6412 6276 6440
rect 4028 6400 4034 6412
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 7466 6440 7472 6452
rect 6840 6412 7472 6440
rect 2774 6332 2780 6384
rect 2832 6372 2838 6384
rect 2869 6375 2927 6381
rect 2869 6372 2881 6375
rect 2832 6344 2881 6372
rect 2832 6332 2838 6344
rect 2869 6341 2881 6344
rect 2915 6341 2927 6375
rect 2869 6335 2927 6341
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 6730 6372 6736 6384
rect 4120 6344 6736 6372
rect 4120 6332 4126 6344
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3513 6307 3571 6313
rect 3513 6304 3525 6307
rect 3016 6276 3525 6304
rect 3016 6264 3022 6276
rect 3513 6273 3525 6276
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 4304 6276 4353 6304
rect 4304 6264 4310 6276
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 5166 6304 5172 6316
rect 5127 6276 5172 6304
rect 4341 6267 4399 6273
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6304 6147 6307
rect 6178 6304 6184 6316
rect 6135 6276 6184 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6840 6313 6868 6412
rect 7466 6400 7472 6412
rect 7524 6440 7530 6452
rect 7742 6440 7748 6452
rect 7524 6412 7748 6440
rect 7524 6400 7530 6412
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 12434 6440 12440 6452
rect 8588 6412 12440 6440
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6236 1547 6239
rect 1578 6236 1584 6248
rect 1535 6208 1584 6236
rect 1535 6205 1547 6208
rect 1489 6199 1547 6205
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 1756 6239 1814 6245
rect 1756 6205 1768 6239
rect 1802 6236 1814 6239
rect 2976 6236 3004 6264
rect 1802 6208 3004 6236
rect 3421 6239 3479 6245
rect 1802 6205 1814 6208
rect 1756 6199 1814 6205
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 4154 6236 4160 6248
rect 3467 6208 4160 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4672 6208 4997 6236
rect 4672 6196 4678 6208
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 4985 6199 5043 6205
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5810 6236 5816 6248
rect 5123 6208 5816 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 7092 6239 7150 6245
rect 7092 6205 7104 6239
rect 7138 6236 7150 6239
rect 8588 6236 8616 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 12529 6443 12587 6449
rect 12529 6409 12541 6443
rect 12575 6440 12587 6443
rect 15378 6440 15384 6452
rect 12575 6412 15384 6440
rect 12575 6409 12587 6412
rect 12529 6403 12587 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 17034 6400 17040 6452
rect 17092 6440 17098 6452
rect 19150 6440 19156 6452
rect 17092 6412 19156 6440
rect 17092 6400 17098 6412
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19426 6440 19432 6452
rect 19339 6412 19432 6440
rect 19426 6400 19432 6412
rect 19484 6440 19490 6452
rect 20438 6440 20444 6452
rect 19484 6412 20444 6440
rect 19484 6400 19490 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 10505 6375 10563 6381
rect 10505 6341 10517 6375
rect 10551 6372 10563 6375
rect 13906 6372 13912 6384
rect 10551 6344 12020 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 11146 6304 11152 6316
rect 11107 6276 11152 6304
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11992 6313 12020 6344
rect 12084 6344 13912 6372
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 7138 6208 8616 6236
rect 8665 6239 8723 6245
rect 7138 6205 7150 6208
rect 7092 6199 7150 6205
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 3329 6171 3387 6177
rect 3329 6137 3341 6171
rect 3375 6168 3387 6171
rect 7742 6168 7748 6180
rect 3375 6140 3832 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 3804 6109 3832 6140
rect 4172 6140 7748 6168
rect 4172 6109 4200 6140
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 7834 6128 7840 6180
rect 7892 6168 7898 6180
rect 8680 6168 8708 6199
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 11885 6239 11943 6245
rect 10560 6208 11652 6236
rect 10560 6196 10566 6208
rect 7892 6140 8708 6168
rect 7892 6128 7898 6140
rect 8846 6128 8852 6180
rect 8904 6177 8910 6180
rect 8904 6171 8968 6177
rect 8904 6137 8922 6171
rect 8956 6168 8968 6171
rect 10226 6168 10232 6180
rect 8956 6140 10232 6168
rect 8956 6137 8968 6140
rect 8904 6131 8968 6137
rect 8904 6128 8910 6131
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 10652 6140 10977 6168
rect 10652 6128 10658 6140
rect 10965 6137 10977 6140
rect 11011 6137 11023 6171
rect 10965 6131 11023 6137
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6069 3847 6103
rect 3789 6063 3847 6069
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6069 4215 6103
rect 4157 6063 4215 6069
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4295 6072 4629 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 5442 6100 5448 6112
rect 5403 6072 5448 6100
rect 4617 6063 4675 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 5813 6103 5871 6109
rect 5813 6100 5825 6103
rect 5776 6072 5825 6100
rect 5776 6060 5782 6072
rect 5813 6069 5825 6072
rect 5859 6069 5871 6103
rect 5813 6063 5871 6069
rect 5905 6103 5963 6109
rect 5905 6069 5917 6103
rect 5951 6100 5963 6103
rect 6546 6100 6552 6112
rect 5951 6072 6552 6100
rect 5951 6069 5963 6072
rect 5905 6063 5963 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8662 6100 8668 6112
rect 8251 6072 8668 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9640 6072 10057 6100
rect 9640 6060 9646 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10192 6072 10885 6100
rect 10192 6060 10198 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 11514 6100 11520 6112
rect 11475 6072 11520 6100
rect 10873 6063 10931 6069
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 11624 6100 11652 6208
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 12084 6236 12112 6344
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 13998 6332 14004 6384
rect 14056 6332 14062 6384
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6304 12219 6307
rect 12250 6304 12256 6316
rect 12207 6276 12256 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 12250 6264 12256 6276
rect 12308 6304 12314 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 12308 6276 13093 6304
rect 12308 6264 12314 6276
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 14016 6304 14044 6332
rect 13081 6267 13139 6273
rect 13188 6276 14044 6304
rect 11931 6208 12112 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 12768 6208 13001 6236
rect 12768 6196 12774 6208
rect 12989 6205 13001 6208
rect 13035 6205 13047 6239
rect 13188 6236 13216 6276
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15712 6276 15853 6304
rect 15712 6264 15718 6276
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 19981 6307 20039 6313
rect 19981 6273 19993 6307
rect 20027 6304 20039 6307
rect 20162 6304 20168 6316
rect 20027 6276 20168 6304
rect 20027 6273 20039 6276
rect 19981 6267 20039 6273
rect 20162 6264 20168 6276
rect 20220 6264 20226 6316
rect 20806 6304 20812 6316
rect 20767 6276 20812 6304
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 12989 6199 13047 6205
rect 13096 6208 13216 6236
rect 13909 6239 13967 6245
rect 11698 6128 11704 6180
rect 11756 6168 11762 6180
rect 12894 6168 12900 6180
rect 11756 6140 12388 6168
rect 12855 6140 12900 6168
rect 11756 6128 11762 6140
rect 11974 6100 11980 6112
rect 11624 6072 11980 6100
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12360 6100 12388 6140
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 13096 6100 13124 6208
rect 13909 6205 13921 6239
rect 13955 6236 13967 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13955 6208 14013 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 16108 6239 16166 6245
rect 16108 6205 16120 6239
rect 16154 6236 16166 6239
rect 17218 6236 17224 6248
rect 16154 6208 17224 6236
rect 16154 6205 16166 6208
rect 16108 6199 16166 6205
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17972 6208 18061 6236
rect 14268 6171 14326 6177
rect 14268 6137 14280 6171
rect 14314 6168 14326 6171
rect 14314 6140 15976 6168
rect 14314 6137 14326 6140
rect 14268 6131 14326 6137
rect 15948 6112 15976 6140
rect 16666 6128 16672 6180
rect 16724 6168 16730 6180
rect 17862 6168 17868 6180
rect 16724 6140 17868 6168
rect 16724 6128 16730 6140
rect 17862 6128 17868 6140
rect 17920 6168 17926 6180
rect 17972 6168 18000 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 19610 6196 19616 6248
rect 19668 6196 19674 6248
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 20717 6239 20775 6245
rect 20717 6236 20729 6239
rect 20680 6208 20729 6236
rect 20680 6196 20686 6208
rect 20717 6205 20729 6208
rect 20763 6205 20775 6239
rect 20717 6199 20775 6205
rect 17920 6140 18000 6168
rect 18316 6171 18374 6177
rect 17920 6128 17926 6140
rect 18316 6137 18328 6171
rect 18362 6168 18374 6171
rect 19242 6168 19248 6180
rect 18362 6140 19248 6168
rect 18362 6137 18374 6140
rect 18316 6131 18374 6137
rect 19242 6128 19248 6140
rect 19300 6128 19306 6180
rect 19628 6168 19656 6196
rect 20162 6168 20168 6180
rect 19628 6140 20168 6168
rect 20162 6128 20168 6140
rect 20220 6168 20226 6180
rect 20220 6140 20668 6168
rect 20220 6128 20226 6140
rect 13906 6100 13912 6112
rect 12360 6072 13124 6100
rect 13819 6072 13912 6100
rect 13906 6060 13912 6072
rect 13964 6100 13970 6112
rect 14366 6100 14372 6112
rect 13964 6072 14372 6100
rect 13964 6060 13970 6072
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 15381 6103 15439 6109
rect 15381 6100 15393 6103
rect 15068 6072 15393 6100
rect 15068 6060 15074 6072
rect 15381 6069 15393 6072
rect 15427 6069 15439 6103
rect 15381 6063 15439 6069
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 17221 6103 17279 6109
rect 17221 6100 17233 6103
rect 15988 6072 17233 6100
rect 15988 6060 15994 6072
rect 17221 6069 17233 6072
rect 17267 6069 17279 6103
rect 17221 6063 17279 6069
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 20640 6109 20668 6140
rect 20257 6103 20315 6109
rect 20257 6100 20269 6103
rect 19668 6072 20269 6100
rect 19668 6060 19674 6072
rect 20257 6069 20269 6072
rect 20303 6069 20315 6103
rect 20257 6063 20315 6069
rect 20625 6103 20683 6109
rect 20625 6069 20637 6103
rect 20671 6069 20683 6103
rect 20625 6063 20683 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 2958 5896 2964 5908
rect 2919 5868 2964 5896
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 3510 5856 3516 5908
rect 3568 5856 3574 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4120 5868 6316 5896
rect 4120 5856 4126 5868
rect 1762 5788 1768 5840
rect 1820 5828 1826 5840
rect 3421 5831 3479 5837
rect 3421 5828 3433 5831
rect 1820 5800 3433 5828
rect 1820 5788 1826 5800
rect 3421 5797 3433 5800
rect 3467 5828 3479 5831
rect 3528 5828 3556 5856
rect 3467 5800 3556 5828
rect 4341 5831 4399 5837
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 4341 5797 4353 5831
rect 4387 5828 4399 5831
rect 4893 5831 4951 5837
rect 4893 5828 4905 5831
rect 4387 5800 4905 5828
rect 4387 5797 4399 5800
rect 4341 5791 4399 5797
rect 4893 5797 4905 5800
rect 4939 5828 4951 5831
rect 5074 5828 5080 5840
rect 4939 5800 5080 5828
rect 4939 5797 4951 5800
rect 4893 5791 4951 5797
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5629 5831 5687 5837
rect 5629 5797 5641 5831
rect 5675 5828 5687 5831
rect 6178 5828 6184 5840
rect 5675 5800 6184 5828
rect 5675 5797 5687 5800
rect 5629 5791 5687 5797
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 6288 5828 6316 5868
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 6420 5868 6561 5896
rect 6420 5856 6426 5868
rect 6549 5865 6561 5868
rect 6595 5865 6607 5899
rect 6549 5859 6607 5865
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7558 5896 7564 5908
rect 6972 5868 7564 5896
rect 6972 5856 6978 5868
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 7800 5868 8125 5896
rect 7800 5856 7806 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 9490 5896 9496 5908
rect 8260 5868 9496 5896
rect 8260 5856 8266 5868
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 10226 5896 10232 5908
rect 10183 5868 10232 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10744 5868 10885 5896
rect 10744 5856 10750 5868
rect 10873 5865 10885 5868
rect 10919 5896 10931 5899
rect 11790 5896 11796 5908
rect 10919 5868 11796 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 11885 5899 11943 5905
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 12066 5896 12072 5908
rect 11931 5868 12072 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 14182 5896 14188 5908
rect 12943 5868 14188 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 15289 5899 15347 5905
rect 15289 5896 15301 5899
rect 14783 5868 15301 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15289 5865 15301 5868
rect 15335 5865 15347 5899
rect 15289 5859 15347 5865
rect 15378 5856 15384 5908
rect 15436 5896 15442 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15436 5868 15761 5896
rect 15436 5856 15442 5868
rect 15749 5865 15761 5868
rect 15795 5896 15807 5899
rect 17862 5896 17868 5908
rect 15795 5868 17868 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18233 5899 18291 5905
rect 18233 5896 18245 5899
rect 18012 5868 18245 5896
rect 18012 5856 18018 5868
rect 18233 5865 18245 5868
rect 18279 5865 18291 5899
rect 18233 5859 18291 5865
rect 18601 5899 18659 5905
rect 18601 5865 18613 5899
rect 18647 5896 18659 5899
rect 18782 5896 18788 5908
rect 18647 5868 18788 5896
rect 18647 5865 18659 5868
rect 18601 5859 18659 5865
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 19521 5899 19579 5905
rect 19521 5865 19533 5899
rect 19567 5896 19579 5899
rect 19981 5899 20039 5905
rect 19981 5896 19993 5899
rect 19567 5868 19993 5896
rect 19567 5865 19579 5868
rect 19521 5859 19579 5865
rect 19981 5865 19993 5868
rect 20027 5865 20039 5899
rect 19981 5859 20039 5865
rect 20070 5856 20076 5908
rect 20128 5896 20134 5908
rect 20349 5899 20407 5905
rect 20349 5896 20361 5899
rect 20128 5868 20361 5896
rect 20128 5856 20134 5868
rect 20349 5865 20361 5868
rect 20395 5865 20407 5899
rect 20349 5859 20407 5865
rect 6457 5831 6515 5837
rect 6457 5828 6469 5831
rect 6288 5800 6469 5828
rect 6457 5797 6469 5800
rect 6503 5828 6515 5831
rect 6730 5828 6736 5840
rect 6503 5800 6736 5828
rect 6503 5797 6515 5800
rect 6457 5791 6515 5797
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 7653 5831 7711 5837
rect 7653 5828 7665 5831
rect 6880 5800 7665 5828
rect 6880 5788 6886 5800
rect 7653 5797 7665 5800
rect 7699 5797 7711 5831
rect 7653 5791 7711 5797
rect 8481 5831 8539 5837
rect 8481 5797 8493 5831
rect 8527 5828 8539 5831
rect 10778 5828 10784 5840
rect 8527 5800 10784 5828
rect 8527 5797 8539 5800
rect 8481 5791 8539 5797
rect 10778 5788 10784 5800
rect 10836 5828 10842 5840
rect 11698 5828 11704 5840
rect 10836 5800 11704 5828
rect 10836 5788 10842 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 19061 5831 19119 5837
rect 12308 5800 15516 5828
rect 12308 5788 12314 5800
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 1848 5763 1906 5769
rect 1848 5729 1860 5763
rect 1894 5760 1906 5763
rect 2682 5760 2688 5772
rect 1894 5732 2688 5760
rect 1894 5729 1906 5732
rect 1848 5723 1906 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 4062 5760 4068 5772
rect 3559 5732 4068 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 4062 5720 4068 5732
rect 4120 5760 4126 5772
rect 4706 5760 4712 5772
rect 4120 5732 4712 5760
rect 4120 5720 4126 5732
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5760 4859 5763
rect 5350 5760 5356 5772
rect 4847 5732 5356 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 5350 5720 5356 5732
rect 5408 5760 5414 5772
rect 6546 5760 6552 5772
rect 5408 5732 6552 5760
rect 5408 5720 5414 5732
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 7190 5720 7196 5732
rect 7248 5760 7254 5772
rect 7742 5760 7748 5772
rect 7248 5732 7748 5760
rect 7248 5720 7254 5732
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 8570 5760 8576 5772
rect 8531 5732 8576 5760
rect 8570 5720 8576 5732
rect 8628 5760 8634 5772
rect 9214 5760 9220 5772
rect 8628 5732 9220 5760
rect 8628 5720 8634 5732
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 10796 5732 13277 5760
rect 3694 5692 3700 5704
rect 3607 5664 3700 5692
rect 3694 5652 3700 5664
rect 3752 5692 3758 5704
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 3752 5664 5089 5692
rect 3752 5652 3758 5664
rect 5077 5661 5089 5664
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5092 5624 5120 5655
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5592 5664 5733 5692
rect 5592 5652 5598 5664
rect 5721 5661 5733 5664
rect 5767 5692 5779 5695
rect 5810 5692 5816 5704
rect 5767 5664 5816 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 6730 5692 6736 5704
rect 6691 5664 6736 5692
rect 5905 5655 5963 5661
rect 5166 5624 5172 5636
rect 5079 5596 5172 5624
rect 5166 5584 5172 5596
rect 5224 5624 5230 5636
rect 5920 5624 5948 5655
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8386 5692 8392 5704
rect 7975 5664 8392 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8662 5692 8668 5704
rect 8623 5664 8668 5692
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9950 5692 9956 5704
rect 9416 5664 9956 5692
rect 8680 5624 8708 5652
rect 5224 5596 8708 5624
rect 5224 5584 5230 5596
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 4433 5559 4491 5565
rect 3108 5528 3153 5556
rect 3108 5516 3114 5528
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 5074 5556 5080 5568
rect 4479 5528 5080 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 5258 5556 5264 5568
rect 5219 5528 5264 5556
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6270 5556 6276 5568
rect 6135 5528 6276 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 9416 5556 9444 5664
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10284 5664 10329 5692
rect 10284 5652 10290 5664
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 10796 5624 10824 5732
rect 13265 5729 13277 5732
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 13722 5760 13728 5772
rect 13403 5732 13728 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14829 5763 14887 5769
rect 14829 5729 14841 5763
rect 14875 5760 14887 5763
rect 15194 5760 15200 5772
rect 14875 5732 15200 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10928 5664 10977 5692
rect 10928 5652 10934 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11112 5664 11157 5692
rect 11112 5652 11118 5664
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11974 5692 11980 5704
rect 11296 5664 11980 5692
rect 11296 5652 11302 5664
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 14182 5692 14188 5704
rect 13587 5664 14188 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 9548 5596 10824 5624
rect 11072 5624 11100 5652
rect 12084 5624 12112 5655
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 15010 5692 15016 5704
rect 14971 5664 15016 5692
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15102 5624 15108 5636
rect 11072 5596 12112 5624
rect 12176 5596 15108 5624
rect 9548 5584 9554 5596
rect 9674 5556 9680 5568
rect 7616 5528 9444 5556
rect 9635 5528 9680 5556
rect 7616 5516 7622 5528
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 10502 5556 10508 5568
rect 10463 5528 10508 5556
rect 10502 5516 10508 5528
rect 10560 5516 10566 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 10870 5556 10876 5568
rect 10744 5528 10876 5556
rect 10744 5516 10750 5528
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 11517 5559 11575 5565
rect 11517 5525 11529 5559
rect 11563 5556 11575 5559
rect 11698 5556 11704 5568
rect 11563 5528 11704 5556
rect 11563 5525 11575 5528
rect 11517 5519 11575 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12176 5556 12204 5596
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 14366 5556 14372 5568
rect 12032 5528 12204 5556
rect 14327 5528 14372 5556
rect 12032 5516 12038 5528
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 15488 5556 15516 5800
rect 18524 5800 18828 5828
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 15838 5760 15844 5772
rect 15703 5732 15844 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 17017 5763 17075 5769
rect 17017 5760 17029 5763
rect 16080 5732 17029 5760
rect 16080 5720 16086 5732
rect 17017 5729 17029 5732
rect 17063 5760 17075 5763
rect 18524 5760 18552 5800
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 17063 5732 18552 5760
rect 18616 5732 18705 5760
rect 17063 5729 17075 5732
rect 17017 5723 17075 5729
rect 15930 5692 15936 5704
rect 15891 5664 15936 5692
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 15654 5584 15660 5636
rect 15712 5624 15718 5636
rect 16666 5624 16672 5636
rect 15712 5596 16672 5624
rect 15712 5584 15718 5596
rect 16666 5584 16672 5596
rect 16724 5624 16730 5636
rect 16776 5624 16804 5655
rect 17954 5652 17960 5704
rect 18012 5692 18018 5704
rect 18616 5692 18644 5732
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 18800 5760 18828 5800
rect 19061 5797 19073 5831
rect 19107 5828 19119 5831
rect 19426 5828 19432 5840
rect 19107 5800 19432 5828
rect 19107 5797 19119 5800
rect 19061 5791 19119 5797
rect 19426 5788 19432 5800
rect 19484 5788 19490 5840
rect 19610 5828 19616 5840
rect 19571 5800 19616 5828
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 20530 5828 20536 5840
rect 20456 5800 20536 5828
rect 18800 5732 20208 5760
rect 18800 5701 18828 5732
rect 18012 5664 18644 5692
rect 18785 5695 18843 5701
rect 18012 5652 18018 5664
rect 18785 5661 18797 5695
rect 18831 5661 18843 5695
rect 18785 5655 18843 5661
rect 19242 5652 19248 5704
rect 19300 5692 19306 5704
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19300 5664 19717 5692
rect 19300 5652 19306 5664
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 16724 5596 16804 5624
rect 18141 5627 18199 5633
rect 16724 5584 16730 5596
rect 18141 5593 18153 5627
rect 18187 5624 18199 5627
rect 19260 5624 19288 5652
rect 18187 5596 19288 5624
rect 20180 5624 20208 5732
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20456 5701 20484 5800
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 20441 5695 20499 5701
rect 20441 5692 20453 5695
rect 20312 5664 20453 5692
rect 20312 5652 20318 5664
rect 20441 5661 20453 5664
rect 20487 5661 20499 5695
rect 20441 5655 20499 5661
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 20548 5624 20576 5655
rect 20714 5624 20720 5636
rect 20180 5596 20720 5624
rect 18187 5593 18199 5596
rect 18141 5587 18199 5593
rect 20714 5584 20720 5596
rect 20772 5584 20778 5636
rect 19061 5559 19119 5565
rect 19061 5556 19073 5559
rect 15488 5528 19073 5556
rect 19061 5525 19073 5528
rect 19107 5525 19119 5559
rect 19061 5519 19119 5525
rect 19153 5559 19211 5565
rect 19153 5525 19165 5559
rect 19199 5556 19211 5559
rect 20070 5556 20076 5568
rect 19199 5528 20076 5556
rect 19199 5525 19211 5528
rect 19153 5519 19211 5525
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2130 5352 2136 5364
rect 2091 5324 2136 5352
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 3568 5324 4108 5352
rect 3568 5312 3574 5324
rect 4080 5284 4108 5324
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4212 5324 4629 5352
rect 4212 5312 4218 5324
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 4617 5315 4675 5321
rect 4982 5312 4988 5364
rect 5040 5352 5046 5364
rect 8846 5352 8852 5364
rect 5040 5324 8432 5352
rect 8807 5324 8852 5352
rect 5040 5312 5046 5324
rect 6362 5284 6368 5296
rect 4080 5256 6368 5284
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 8404 5284 8432 5324
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9122 5312 9128 5364
rect 9180 5352 9186 5364
rect 9398 5352 9404 5364
rect 9180 5324 9404 5352
rect 9180 5312 9186 5324
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 10226 5312 10232 5364
rect 10284 5352 10290 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 10284 5324 11805 5352
rect 10284 5312 10290 5324
rect 11793 5321 11805 5324
rect 11839 5321 11851 5355
rect 11793 5315 11851 5321
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 13998 5352 14004 5364
rect 13044 5324 14004 5352
rect 13044 5312 13050 5324
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 14148 5324 14381 5352
rect 14148 5312 14154 5324
rect 14369 5321 14381 5324
rect 14415 5321 14427 5355
rect 15194 5352 15200 5364
rect 15155 5324 15200 5352
rect 14369 5315 14427 5321
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 18874 5352 18880 5364
rect 18835 5324 18880 5352
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19705 5355 19763 5361
rect 19705 5352 19717 5355
rect 19392 5324 19717 5352
rect 19392 5312 19398 5324
rect 19705 5321 19717 5324
rect 19751 5321 19763 5355
rect 19705 5315 19763 5321
rect 12802 5284 12808 5296
rect 8404 5256 10364 5284
rect 2682 5216 2688 5228
rect 2643 5188 2688 5216
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 5074 5216 5080 5228
rect 5035 5188 5080 5216
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 5224 5188 5269 5216
rect 5224 5176 5230 5188
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6178 5216 6184 5228
rect 5684 5188 6184 5216
rect 5684 5176 5690 5188
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6730 5216 6736 5228
rect 6595 5188 6736 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 7282 5216 7288 5228
rect 6880 5188 7288 5216
rect 6880 5176 6886 5188
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 10042 5216 10048 5228
rect 9355 5188 10048 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10192 5188 10237 5216
rect 10192 5176 10198 5188
rect 2498 5148 2504 5160
rect 2459 5120 2504 5148
rect 2498 5108 2504 5120
rect 2556 5108 2562 5160
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5148 2651 5151
rect 3050 5148 3056 5160
rect 2639 5120 3056 5148
rect 2639 5117 2651 5120
rect 2593 5111 2651 5117
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 3412 5151 3470 5157
rect 3412 5117 3424 5151
rect 3458 5148 3470 5151
rect 3694 5148 3700 5160
rect 3458 5120 3700 5148
rect 3458 5117 3470 5120
rect 3412 5111 3470 5117
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 3160 5080 3188 5111
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5258 5148 5264 5160
rect 5031 5120 5264 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 9950 5148 9956 5160
rect 6196 5120 7420 5148
rect 3602 5080 3608 5092
rect 2924 5052 3608 5080
rect 2924 5040 2930 5052
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 6196 5080 6224 5120
rect 4120 5052 6224 5080
rect 6273 5083 6331 5089
rect 4120 5040 4126 5052
rect 6273 5049 6285 5083
rect 6319 5080 6331 5083
rect 6825 5083 6883 5089
rect 6825 5080 6837 5083
rect 6319 5052 6837 5080
rect 6319 5049 6331 5052
rect 6273 5043 6331 5049
rect 6825 5049 6837 5052
rect 6871 5049 6883 5083
rect 7392 5080 7420 5120
rect 7668 5120 9956 5148
rect 7668 5080 7696 5120
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 7392 5052 7696 5080
rect 7736 5083 7794 5089
rect 6825 5043 6883 5049
rect 7736 5049 7748 5083
rect 7782 5049 7794 5083
rect 10336 5080 10364 5256
rect 11440 5256 12808 5284
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5148 10471 5151
rect 10962 5148 10968 5160
rect 10459 5120 10968 5148
rect 10459 5117 10471 5120
rect 10413 5111 10471 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 10680 5083 10738 5089
rect 10336 5052 10640 5080
rect 7736 5043 7794 5049
rect 1857 5015 1915 5021
rect 1857 4981 1869 5015
rect 1903 5012 1915 5015
rect 2222 5012 2228 5024
rect 1903 4984 2228 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 2740 4984 4537 5012
rect 2740 4972 2746 4984
rect 4525 4981 4537 4984
rect 4571 5012 4583 5015
rect 5166 5012 5172 5024
rect 4571 4984 5172 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 6178 5012 6184 5024
rect 5951 4984 6184 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 5012 6423 5015
rect 6546 5012 6552 5024
rect 6411 4984 6552 5012
rect 6411 4981 6423 4984
rect 6365 4975 6423 4981
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 7558 4972 7564 5024
rect 7616 5012 7622 5024
rect 7751 5012 7779 5043
rect 9582 5012 9588 5024
rect 7616 4984 7779 5012
rect 9543 4984 9588 5012
rect 7616 4972 7622 4984
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 10045 5015 10103 5021
rect 10045 4981 10057 5015
rect 10091 5012 10103 5015
rect 10318 5012 10324 5024
rect 10091 4984 10324 5012
rect 10091 4981 10103 4984
rect 10045 4975 10103 4981
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 10612 5012 10640 5052
rect 10680 5049 10692 5083
rect 10726 5080 10738 5083
rect 11054 5080 11060 5092
rect 10726 5052 11060 5080
rect 10726 5049 10738 5052
rect 10680 5043 10738 5049
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11440 5012 11468 5256
rect 12802 5244 12808 5256
rect 12860 5284 12866 5296
rect 12860 5256 14044 5284
rect 12860 5244 12866 5256
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 11940 5188 13124 5216
rect 11940 5176 11946 5188
rect 13096 5148 13124 5188
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 13906 5216 13912 5228
rect 13320 5188 13912 5216
rect 13320 5176 13326 5188
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 14016 5225 14044 5256
rect 16114 5244 16120 5296
rect 16172 5284 16178 5296
rect 17402 5284 17408 5296
rect 16172 5256 17408 5284
rect 16172 5244 16178 5256
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 18049 5287 18107 5293
rect 18049 5253 18061 5287
rect 18095 5284 18107 5287
rect 19518 5284 19524 5296
rect 18095 5256 19524 5284
rect 18095 5253 18107 5256
rect 18049 5247 18107 5253
rect 19518 5244 19524 5256
rect 19576 5244 19582 5296
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14182 5216 14188 5228
rect 14095 5188 14188 5216
rect 14001 5179 14059 5185
rect 14182 5176 14188 5188
rect 14240 5216 14246 5228
rect 15013 5219 15071 5225
rect 15013 5216 15025 5219
rect 14240 5188 15025 5216
rect 14240 5176 14246 5188
rect 15013 5185 15025 5188
rect 15059 5216 15071 5219
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15059 5188 15853 5216
rect 15059 5185 15071 5188
rect 15013 5179 15071 5185
rect 15841 5185 15853 5188
rect 15887 5216 15899 5219
rect 15930 5216 15936 5228
rect 15887 5188 15936 5216
rect 15887 5185 15899 5188
rect 15841 5179 15899 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 17129 5219 17187 5225
rect 17129 5216 17141 5219
rect 16632 5188 17141 5216
rect 16632 5176 16638 5188
rect 17129 5185 17141 5188
rect 17175 5216 17187 5219
rect 17586 5216 17592 5228
rect 17175 5188 17592 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 18564 5188 18613 5216
rect 18564 5176 18570 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 19242 5176 19248 5228
rect 19300 5216 19306 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19300 5188 19441 5216
rect 19300 5176 19306 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19429 5179 19487 5185
rect 19536 5188 20177 5216
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 13096 5120 14749 5148
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 15654 5148 15660 5160
rect 15615 5120 15660 5148
rect 14737 5111 14795 5117
rect 15654 5108 15660 5120
rect 15712 5148 15718 5160
rect 16114 5148 16120 5160
rect 15712 5120 16120 5148
rect 15712 5108 15718 5120
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 16942 5148 16948 5160
rect 16899 5120 16948 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 16942 5108 16948 5120
rect 17000 5148 17006 5160
rect 17678 5148 17684 5160
rect 17000 5120 17684 5148
rect 17000 5108 17006 5120
rect 17678 5108 17684 5120
rect 17736 5108 17742 5160
rect 19150 5108 19156 5160
rect 19208 5148 19214 5160
rect 19536 5148 19564 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 20349 5219 20407 5225
rect 20349 5185 20361 5219
rect 20395 5216 20407 5219
rect 20438 5216 20444 5228
rect 20395 5188 20444 5216
rect 20395 5185 20407 5188
rect 20349 5179 20407 5185
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 20898 5216 20904 5228
rect 20855 5188 20904 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 20898 5176 20904 5188
rect 20956 5176 20962 5228
rect 20070 5148 20076 5160
rect 19208 5120 19564 5148
rect 20031 5120 20076 5148
rect 19208 5108 19214 5120
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 11514 5040 11520 5092
rect 11572 5080 11578 5092
rect 17954 5080 17960 5092
rect 11572 5052 17960 5080
rect 11572 5040 11578 5052
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 18046 5040 18052 5092
rect 18104 5080 18110 5092
rect 19337 5083 19395 5089
rect 19337 5080 19349 5083
rect 18104 5052 19349 5080
rect 18104 5040 18110 5052
rect 19337 5049 19349 5052
rect 19383 5049 19395 5083
rect 19337 5043 19395 5049
rect 10612 4984 11468 5012
rect 13262 4972 13268 5024
rect 13320 5012 13326 5024
rect 13357 5015 13415 5021
rect 13357 5012 13369 5015
rect 13320 4984 13369 5012
rect 13320 4972 13326 4984
rect 13357 4981 13369 4984
rect 13403 4981 13415 5015
rect 13538 5012 13544 5024
rect 13499 4984 13544 5012
rect 13357 4975 13415 4981
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 13906 5012 13912 5024
rect 13867 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14829 5015 14887 5021
rect 14829 5012 14841 5015
rect 14056 4984 14841 5012
rect 14056 4972 14062 4984
rect 14829 4981 14841 4984
rect 14875 4981 14887 5015
rect 15562 5012 15568 5024
rect 15523 4984 15568 5012
rect 14829 4975 14887 4981
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 16485 5015 16543 5021
rect 16485 4981 16497 5015
rect 16531 5012 16543 5015
rect 16758 5012 16764 5024
rect 16531 4984 16764 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 16945 5015 17003 5021
rect 16945 5012 16957 5015
rect 16908 4984 16957 5012
rect 16908 4972 16914 4984
rect 16945 4981 16957 4984
rect 16991 4981 17003 5015
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 16945 4975 17003 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 18509 5015 18567 5021
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 18598 5012 18604 5024
rect 18555 4984 18604 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 18598 4972 18604 4984
rect 18656 4972 18662 5024
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19150 5012 19156 5024
rect 18840 4984 19156 5012
rect 18840 4972 18846 4984
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 19245 5015 19303 5021
rect 19245 4981 19257 5015
rect 19291 5012 19303 5015
rect 19426 5012 19432 5024
rect 19291 4984 19432 5012
rect 19291 4981 19303 4984
rect 19245 4975 19303 4981
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 2038 4808 2044 4820
rect 1903 4780 2044 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 5353 4811 5411 4817
rect 5353 4808 5365 4811
rect 4939 4780 5365 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5353 4777 5365 4780
rect 5399 4808 5411 4811
rect 5994 4808 6000 4820
rect 5399 4780 6000 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6178 4808 6184 4820
rect 6139 4780 6184 4808
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6880 4780 7021 4808
rect 6880 4768 6886 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7009 4771 7067 4777
rect 7101 4811 7159 4817
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 7147 4780 7481 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 7469 4777 7481 4780
rect 7515 4777 7527 4811
rect 7469 4771 7527 4777
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9582 4808 9588 4820
rect 9263 4780 9588 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 10318 4808 10324 4820
rect 10279 4780 10324 4808
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 10502 4768 10508 4820
rect 10560 4808 10566 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 10560 4780 11621 4808
rect 10560 4768 10566 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 12342 4808 12348 4820
rect 11609 4771 11667 4777
rect 12268 4780 12348 4808
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 5776 4712 6408 4740
rect 5776 4700 5782 4712
rect 2958 4672 2964 4684
rect 2332 4644 2964 4672
rect 2332 4616 2360 4644
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3418 4672 3424 4684
rect 3379 4644 3424 4672
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 6270 4672 6276 4684
rect 3712 4644 5672 4672
rect 6231 4644 6276 4672
rect 3712 4616 3740 4644
rect 5644 4616 5672 4644
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 6380 4672 6408 4712
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 7837 4743 7895 4749
rect 7837 4740 7849 4743
rect 7340 4712 7849 4740
rect 7340 4700 7346 4712
rect 7837 4709 7849 4712
rect 7883 4740 7895 4743
rect 8294 4740 8300 4752
rect 7883 4712 8300 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8662 4740 8668 4752
rect 8496 4712 8668 4740
rect 7466 4672 7472 4684
rect 6380 4644 7472 4672
rect 7466 4632 7472 4644
rect 7524 4672 7530 4684
rect 8496 4672 8524 4712
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 9125 4743 9183 4749
rect 9125 4709 9137 4743
rect 9171 4740 9183 4743
rect 9674 4740 9680 4752
rect 9171 4712 9680 4740
rect 9171 4709 9183 4712
rect 9125 4703 9183 4709
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 10229 4743 10287 4749
rect 10229 4709 10241 4743
rect 10275 4740 10287 4743
rect 12268 4740 12296 4780
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12618 4808 12624 4820
rect 12579 4780 12624 4808
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 14366 4808 14372 4820
rect 12759 4780 14372 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 18046 4808 18052 4820
rect 15335 4780 18052 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18414 4768 18420 4820
rect 18472 4808 18478 4820
rect 18509 4811 18567 4817
rect 18509 4808 18521 4811
rect 18472 4780 18521 4808
rect 18472 4768 18478 4780
rect 18509 4777 18521 4780
rect 18555 4777 18567 4811
rect 18509 4771 18567 4777
rect 18782 4768 18788 4820
rect 18840 4808 18846 4820
rect 19978 4808 19984 4820
rect 18840 4780 19984 4808
rect 18840 4768 18846 4780
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 15749 4743 15807 4749
rect 15749 4740 15761 4743
rect 10275 4712 12296 4740
rect 12360 4712 15761 4740
rect 10275 4709 10287 4712
rect 10229 4703 10287 4709
rect 10686 4672 10692 4684
rect 7524 4644 8524 4672
rect 8588 4644 10692 4672
rect 7524 4632 7530 4644
rect 2314 4604 2320 4616
rect 2275 4576 2320 4604
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 2682 4604 2688 4616
rect 2547 4576 2688 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 3513 4607 3571 4613
rect 3513 4604 3525 4607
rect 3384 4576 3525 4604
rect 3384 4564 3390 4576
rect 3513 4573 3525 4576
rect 3559 4573 3571 4607
rect 3694 4604 3700 4616
rect 3607 4576 3700 4604
rect 3513 4567 3571 4573
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 4764 4576 5457 4604
rect 4764 4564 4770 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5626 4604 5632 4616
rect 5587 4576 5632 4604
rect 5445 4567 5503 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 5776 4576 6377 4604
rect 5776 4564 5782 4576
rect 6365 4573 6377 4576
rect 6411 4604 6423 4607
rect 6822 4604 6828 4616
rect 6411 4576 6828 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 6822 4564 6828 4576
rect 6880 4604 6886 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6880 4576 7205 4604
rect 6880 4564 6886 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7800 4576 7941 4604
rect 7800 4564 7806 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8478 4604 8484 4616
rect 8159 4576 8484 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 8588 4536 8616 4644
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 11204 4644 11529 4672
rect 11204 4632 11210 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12360 4672 12388 4712
rect 15749 4709 15761 4712
rect 15795 4709 15807 4743
rect 15749 4703 15807 4709
rect 17034 4700 17040 4752
rect 17092 4740 17098 4752
rect 17304 4743 17362 4749
rect 17304 4740 17316 4743
rect 17092 4712 17316 4740
rect 17092 4700 17098 4712
rect 17304 4709 17316 4712
rect 17350 4740 17362 4743
rect 17350 4712 19104 4740
rect 17350 4709 17362 4712
rect 17304 4703 17362 4709
rect 13078 4672 13084 4684
rect 12032 4644 12388 4672
rect 13039 4644 13084 4672
rect 12032 4632 12038 4644
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13348 4675 13406 4681
rect 13348 4641 13360 4675
rect 13394 4672 13406 4675
rect 13906 4672 13912 4684
rect 13394 4644 13912 4672
rect 13394 4641 13406 4644
rect 13348 4635 13406 4641
rect 13906 4632 13912 4644
rect 13964 4632 13970 4684
rect 14090 4632 14096 4684
rect 14148 4632 14154 4684
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 16206 4672 16212 4684
rect 15764 4644 16212 4672
rect 9398 4604 9404 4616
rect 9359 4576 9404 4604
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10060 4576 10241 4604
rect 4120 4508 8616 4536
rect 4120 4496 4126 4508
rect 9214 4496 9220 4548
rect 9272 4536 9278 4548
rect 10060 4536 10088 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10594 4564 10600 4616
rect 10652 4604 10658 4616
rect 10781 4607 10839 4613
rect 10781 4604 10793 4607
rect 10652 4576 10793 4604
rect 10652 4564 10658 4576
rect 10781 4573 10793 4576
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11054 4604 11060 4616
rect 11011 4576 11060 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 11054 4564 11060 4576
rect 11112 4604 11118 4616
rect 11606 4604 11612 4616
rect 11112 4576 11612 4604
rect 11112 4564 11118 4576
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4573 12955 4607
rect 14108 4604 14136 4632
rect 15764 4604 15792 4644
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 16942 4672 16948 4684
rect 16448 4644 16948 4672
rect 16448 4632 16454 4644
rect 16942 4632 16948 4644
rect 17000 4632 17006 4684
rect 18874 4672 18880 4684
rect 18835 4644 18880 4672
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 14108 4576 15792 4604
rect 15933 4607 15991 4613
rect 12897 4567 12955 4573
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16022 4604 16028 4616
rect 15979 4576 16028 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 9272 4508 10088 4536
rect 9272 4496 9278 4508
rect 10134 4496 10140 4548
rect 10192 4536 10198 4548
rect 11716 4536 11744 4567
rect 11790 4536 11796 4548
rect 10192 4508 11796 4536
rect 10192 4496 10198 4508
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3053 4471 3111 4477
rect 3053 4468 3065 4471
rect 2832 4440 3065 4468
rect 2832 4428 2838 4440
rect 3053 4437 3065 4440
rect 3099 4437 3111 4471
rect 4982 4468 4988 4480
rect 4943 4440 4988 4468
rect 3053 4431 3111 4437
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5810 4468 5816 4480
rect 5771 4440 5816 4468
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 6641 4471 6699 4477
rect 6641 4437 6653 4471
rect 6687 4468 6699 4471
rect 8202 4468 8208 4480
rect 6687 4440 8208 4468
rect 6687 4437 6699 4440
rect 6641 4431 6699 4437
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 8757 4471 8815 4477
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 10042 4468 10048 4480
rect 8803 4440 10048 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11149 4471 11207 4477
rect 11149 4468 11161 4471
rect 11112 4440 11161 4468
rect 11112 4428 11118 4440
rect 11149 4437 11161 4440
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 12253 4471 12311 4477
rect 12253 4437 12265 4471
rect 12299 4468 12311 4471
rect 12710 4468 12716 4480
rect 12299 4440 12716 4468
rect 12299 4437 12311 4440
rect 12253 4431 12311 4437
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 12912 4468 12940 4567
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 16850 4604 16856 4616
rect 16724 4576 16856 4604
rect 16724 4564 16730 4576
rect 16850 4564 16856 4576
rect 16908 4604 16914 4616
rect 17037 4607 17095 4613
rect 17037 4604 17049 4607
rect 16908 4576 17049 4604
rect 16908 4564 16914 4576
rect 17037 4573 17049 4576
rect 17083 4573 17095 4607
rect 18506 4604 18512 4616
rect 17037 4567 17095 4573
rect 18432 4576 18512 4604
rect 13722 4468 13728 4480
rect 12912 4440 13728 4468
rect 13722 4428 13728 4440
rect 13780 4468 13786 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 13780 4440 14473 4468
rect 13780 4428 13786 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 17052 4468 17080 4567
rect 18432 4545 18460 4576
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18966 4604 18972 4616
rect 18927 4576 18972 4604
rect 18966 4564 18972 4576
rect 19024 4564 19030 4616
rect 19076 4613 19104 4712
rect 19610 4681 19616 4684
rect 19337 4675 19395 4681
rect 19337 4641 19349 4675
rect 19383 4672 19395 4675
rect 19383 4644 19463 4672
rect 19383 4641 19395 4644
rect 19337 4635 19395 4641
rect 19061 4607 19119 4613
rect 19061 4573 19073 4607
rect 19107 4573 19119 4607
rect 19435 4604 19463 4644
rect 19604 4635 19616 4681
rect 19668 4672 19674 4684
rect 19668 4644 19704 4672
rect 19610 4632 19616 4635
rect 19668 4632 19674 4644
rect 21266 4632 21272 4684
rect 21324 4672 21330 4684
rect 22186 4672 22192 4684
rect 21324 4644 22192 4672
rect 21324 4632 21330 4644
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 19061 4567 19119 4573
rect 19352 4576 19463 4604
rect 18417 4539 18475 4545
rect 18417 4505 18429 4539
rect 18463 4505 18475 4539
rect 18417 4499 18475 4505
rect 19352 4468 19380 4576
rect 17052 4440 19380 4468
rect 14461 4431 14519 4437
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 4249 4267 4307 4273
rect 4249 4264 4261 4267
rect 2608 4236 4261 4264
rect 2608 4140 2636 4236
rect 4249 4233 4261 4236
rect 4295 4264 4307 4267
rect 4890 4264 4896 4276
rect 4295 4236 4896 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 6788 4236 7604 4264
rect 6788 4224 6794 4236
rect 4724 4168 5028 4196
rect 2590 4128 2596 4140
rect 2551 4100 2596 4128
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 2774 4060 2780 4072
rect 2455 4032 2780 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 3136 4063 3194 4069
rect 3136 4029 3148 4063
rect 3182 4060 3194 4063
rect 3694 4060 3700 4072
rect 3182 4032 3700 4060
rect 3182 4029 3194 4032
rect 3136 4023 3194 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4724 4060 4752 4168
rect 4890 4128 4896 4140
rect 4851 4100 4896 4128
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5000 4128 5028 4168
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 7576 4196 7604 4236
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 7708 4236 8524 4264
rect 7708 4224 7714 4236
rect 6880 4168 7512 4196
rect 7576 4168 8340 4196
rect 6880 4156 6886 4168
rect 5718 4128 5724 4140
rect 5000 4100 5580 4128
rect 5679 4100 5724 4128
rect 4120 4032 4752 4060
rect 4801 4063 4859 4069
rect 4120 4020 4126 4032
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 4982 4060 4988 4072
rect 4847 4032 4988 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 5442 4060 5448 4072
rect 5092 4032 5448 4060
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 5092 3992 5120 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5552 4060 5580 4100
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 7484 4137 7512 4168
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 7469 4091 7527 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8312 4137 8340 4168
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8496 4128 8524 4236
rect 8662 4224 8668 4276
rect 8720 4264 8726 4276
rect 11882 4264 11888 4276
rect 8720 4236 11888 4264
rect 8720 4224 8726 4236
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 12158 4224 12164 4276
rect 12216 4264 12222 4276
rect 18966 4264 18972 4276
rect 12216 4236 18972 4264
rect 12216 4224 12222 4236
rect 18966 4224 18972 4236
rect 19024 4224 19030 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 19705 4267 19763 4273
rect 19705 4264 19717 4267
rect 19668 4236 19717 4264
rect 19668 4224 19674 4236
rect 19705 4233 19717 4236
rect 19751 4233 19763 4267
rect 19705 4227 19763 4233
rect 9950 4156 9956 4208
rect 10008 4196 10014 4208
rect 10226 4196 10232 4208
rect 10008 4168 10232 4196
rect 10008 4156 10014 4168
rect 10226 4156 10232 4168
rect 10284 4156 10290 4208
rect 10505 4199 10563 4205
rect 10505 4165 10517 4199
rect 10551 4196 10563 4199
rect 11146 4196 11152 4208
rect 10551 4168 11152 4196
rect 10551 4165 10563 4168
rect 10505 4159 10563 4165
rect 11146 4156 11152 4168
rect 11204 4156 11210 4208
rect 11790 4156 11796 4208
rect 11848 4196 11854 4208
rect 13722 4196 13728 4208
rect 11848 4168 11928 4196
rect 11848 4156 11854 4168
rect 8757 4131 8815 4137
rect 8757 4128 8769 4131
rect 8496 4100 8769 4128
rect 8297 4091 8355 4097
rect 8757 4097 8769 4100
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 6914 4060 6920 4072
rect 5552 4032 6920 4060
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 8772 4060 8800 4091
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10870 4128 10876 4140
rect 9824 4100 10876 4128
rect 9824 4088 9830 4100
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 11606 4128 11612 4140
rect 11103 4100 11612 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 11606 4088 11612 4100
rect 11664 4128 11670 4140
rect 11900 4137 11928 4168
rect 13188 4168 13728 4196
rect 13188 4137 13216 4168
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 13906 4156 13912 4208
rect 13964 4196 13970 4208
rect 13964 4168 15056 4196
rect 13964 4156 13970 4168
rect 11885 4131 11943 4137
rect 11664 4100 11836 4128
rect 11664 4088 11670 4100
rect 8846 4060 8852 4072
rect 7331 4032 8340 4060
rect 8772 4032 8852 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 8312 4004 8340 4032
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 9024 4063 9082 4069
rect 9024 4029 9036 4063
rect 9070 4060 9082 4063
rect 10134 4060 10140 4072
rect 9070 4032 10140 4060
rect 9070 4029 9082 4032
rect 9024 4023 9082 4029
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 11808 4060 11836 4100
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 14016 4137 14044 4168
rect 15028 4140 15056 4168
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13596 4100 13829 4128
rect 13596 4088 13602 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14826 4128 14832 4140
rect 14787 4100 14832 4128
rect 14001 4091 14059 4097
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15010 4128 15016 4140
rect 14971 4100 15016 4128
rect 15010 4088 15016 4100
rect 15068 4088 15074 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 17034 4128 17040 4140
rect 15988 4100 16896 4128
rect 16995 4100 17040 4128
rect 15988 4088 15994 4100
rect 16868 4072 16896 4100
rect 17034 4088 17040 4100
rect 17092 4128 17098 4140
rect 17310 4128 17316 4140
rect 17092 4100 17316 4128
rect 17092 4088 17098 4100
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 12158 4060 12164 4072
rect 11808 4032 12164 4060
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 13446 4060 13452 4072
rect 12268 4032 13452 4060
rect 4755 3964 5120 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 5629 3995 5687 4001
rect 5629 3992 5641 3995
rect 5408 3964 5641 3992
rect 5408 3952 5414 3964
rect 5629 3961 5641 3964
rect 5675 3961 5687 3995
rect 8113 3995 8171 4001
rect 8113 3992 8125 3995
rect 5629 3955 5687 3961
rect 6932 3964 8125 3992
rect 2038 3924 2044 3936
rect 1999 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 2866 3924 2872 3936
rect 2547 3896 2872 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 3752 3896 4353 3924
rect 3752 3884 3758 3896
rect 4341 3893 4353 3896
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 4672 3896 5181 3924
rect 4672 3884 4678 3896
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 5534 3924 5540 3936
rect 5495 3896 5540 3924
rect 5169 3887 5227 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6932 3933 6960 3964
rect 8113 3961 8125 3964
rect 8159 3961 8171 3995
rect 8113 3955 8171 3961
rect 8294 3952 8300 4004
rect 8352 3952 8358 4004
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 10965 3995 11023 4001
rect 10965 3992 10977 3995
rect 9548 3964 10977 3992
rect 9548 3952 9554 3964
rect 10965 3961 10977 3964
rect 11011 3992 11023 3995
rect 12268 3992 12296 4032
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4060 13783 4063
rect 13906 4060 13912 4072
rect 13771 4032 13912 4060
rect 13771 4029 13783 4032
rect 13725 4023 13783 4029
rect 13906 4020 13912 4032
rect 13964 4060 13970 4072
rect 16482 4060 16488 4072
rect 13964 4032 16488 4060
rect 13964 4020 13970 4032
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16724 4032 16773 4060
rect 16724 4020 16730 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 16850 4020 16856 4072
rect 16908 4060 16914 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 16908 4032 18337 4060
rect 16908 4020 16914 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18592 4063 18650 4069
rect 18592 4060 18604 4063
rect 18325 4023 18383 4029
rect 18524 4032 18604 4060
rect 18524 4004 18552 4032
rect 18592 4029 18604 4032
rect 18638 4060 18650 4063
rect 18966 4060 18972 4072
rect 18638 4032 18972 4060
rect 18638 4029 18650 4032
rect 18592 4023 18650 4029
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 11011 3964 12296 3992
rect 12897 3995 12955 4001
rect 11011 3961 11023 3964
rect 10965 3955 11023 3961
rect 12897 3961 12909 3995
rect 12943 3992 12955 3995
rect 14737 3995 14795 4001
rect 12943 3964 13492 3992
rect 12943 3961 12955 3964
rect 12897 3955 12955 3961
rect 6917 3927 6975 3933
rect 6917 3893 6929 3927
rect 6963 3893 6975 3927
rect 7374 3924 7380 3936
rect 7335 3896 7380 3924
rect 6917 3887 6975 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 8938 3924 8944 3936
rect 7791 3896 8944 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 10134 3924 10140 3936
rect 9456 3896 10140 3924
rect 9456 3884 9462 3896
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 10873 3927 10931 3933
rect 10873 3924 10885 3927
rect 10744 3896 10885 3924
rect 10744 3884 10750 3896
rect 10873 3893 10885 3896
rect 10919 3893 10931 3927
rect 10873 3887 10931 3893
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 11204 3896 11345 3924
rect 11204 3884 11210 3896
rect 11333 3893 11345 3896
rect 11379 3893 11391 3927
rect 11333 3887 11391 3893
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12526 3924 12532 3936
rect 11848 3896 11893 3924
rect 12487 3896 12532 3924
rect 11848 3884 11854 3896
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 12989 3927 13047 3933
rect 12989 3893 13001 3927
rect 13035 3924 13047 3927
rect 13357 3927 13415 3933
rect 13357 3924 13369 3927
rect 13035 3896 13369 3924
rect 13035 3893 13047 3896
rect 12989 3887 13047 3893
rect 13357 3893 13369 3896
rect 13403 3893 13415 3927
rect 13464 3924 13492 3964
rect 14737 3961 14749 3995
rect 14783 3992 14795 3995
rect 15197 3995 15255 4001
rect 15197 3992 15209 3995
rect 14783 3964 15209 3992
rect 14783 3961 14795 3964
rect 14737 3955 14795 3961
rect 15197 3961 15209 3964
rect 15243 3961 15255 3995
rect 15197 3955 15255 3961
rect 18506 3952 18512 4004
rect 18564 3952 18570 4004
rect 14369 3927 14427 3933
rect 14369 3924 14381 3927
rect 13464 3896 14381 3924
rect 13357 3887 13415 3893
rect 14369 3893 14381 3896
rect 14415 3893 14427 3927
rect 14369 3887 14427 3893
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 16206 3924 16212 3936
rect 15620 3896 16212 3924
rect 15620 3884 15626 3896
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 16390 3924 16396 3936
rect 16351 3896 16396 3924
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18874 3924 18880 3936
rect 18095 3896 18880 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 3476 3692 3525 3720
rect 3476 3680 3482 3692
rect 3513 3689 3525 3692
rect 3559 3689 3571 3723
rect 4614 3720 4620 3732
rect 4575 3692 4620 3720
rect 3513 3683 3571 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 4908 3692 6377 3720
rect 2958 3652 2964 3664
rect 2056 3624 2964 3652
rect 2056 3593 2084 3624
rect 2958 3612 2964 3624
rect 3016 3652 3022 3664
rect 4522 3652 4528 3664
rect 3016 3624 4292 3652
rect 4483 3624 4528 3652
rect 3016 3612 3022 3624
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 2308 3587 2366 3593
rect 2308 3553 2320 3587
rect 2354 3584 2366 3587
rect 2590 3584 2596 3596
rect 2354 3556 2596 3584
rect 2354 3553 2366 3556
rect 2308 3547 2366 3553
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 3970 3584 3976 3596
rect 2740 3556 3976 3584
rect 2740 3544 2746 3556
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4264 3584 4292 3624
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 4264 3556 4752 3584
rect 4724 3460 4752 3556
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 4908 3516 4936 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6365 3683 6423 3689
rect 6380 3652 6408 3683
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7800 3692 7941 3720
rect 7800 3680 7806 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 9824 3692 11069 3720
rect 9824 3680 9830 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11057 3683 11115 3689
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 11790 3720 11796 3732
rect 11563 3692 11796 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 11885 3723 11943 3729
rect 11885 3689 11897 3723
rect 11931 3720 11943 3723
rect 12066 3720 12072 3732
rect 11931 3692 12072 3720
rect 11931 3689 11943 3692
rect 11885 3683 11943 3689
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12584 3692 13001 3720
rect 12584 3680 12590 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 14550 3720 14556 3732
rect 12989 3683 13047 3689
rect 13556 3692 14556 3720
rect 13556 3664 13584 3692
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 14829 3723 14887 3729
rect 14829 3689 14841 3723
rect 14875 3689 14887 3723
rect 14829 3683 14887 3689
rect 15473 3723 15531 3729
rect 15473 3689 15485 3723
rect 15519 3720 15531 3723
rect 16850 3720 16856 3732
rect 15519 3692 16856 3720
rect 15519 3689 15531 3692
rect 15473 3683 15531 3689
rect 6730 3661 6736 3664
rect 6724 3652 6736 3661
rect 6380 3624 6736 3652
rect 6724 3615 6736 3624
rect 6730 3612 6736 3615
rect 6788 3612 6794 3664
rect 6822 3612 6828 3664
rect 6880 3652 6886 3664
rect 7650 3652 7656 3664
rect 6880 3624 7656 3652
rect 6880 3612 6886 3624
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8168 3624 8708 3652
rect 8168 3612 8174 3624
rect 5241 3587 5299 3593
rect 5241 3553 5253 3587
rect 5287 3584 5299 3587
rect 5718 3584 5724 3596
rect 5287 3556 5724 3584
rect 5287 3553 5299 3556
rect 5241 3547 5299 3553
rect 5718 3544 5724 3556
rect 5776 3584 5782 3596
rect 6178 3584 6184 3596
rect 5776 3556 6184 3584
rect 5776 3544 5782 3556
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3584 8355 3587
rect 8570 3584 8576 3596
rect 8343 3556 8576 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8680 3584 8708 3624
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 9217 3655 9275 3661
rect 9217 3652 9229 3655
rect 8996 3624 9229 3652
rect 8996 3612 9002 3624
rect 9217 3621 9229 3624
rect 9263 3621 9275 3655
rect 9217 3615 9275 3621
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 11977 3655 12035 3661
rect 11977 3652 11989 3655
rect 11756 3624 11989 3652
rect 11756 3612 11762 3624
rect 11977 3621 11989 3624
rect 12023 3621 12035 3655
rect 11977 3615 12035 3621
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8680 3556 9137 3584
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9223 3556 9444 3584
rect 4847 3488 4936 3516
rect 4985 3519 5043 3525
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 4985 3479 5043 3485
rect 4706 3448 4712 3460
rect 4619 3420 4712 3448
rect 4706 3408 4712 3420
rect 4764 3448 4770 3460
rect 5000 3448 5028 3479
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 8662 3516 8668 3528
rect 8527 3488 8668 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 8110 3448 8116 3460
rect 4764 3420 5028 3448
rect 7392 3420 8116 3448
rect 4764 3408 4770 3420
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3016 3352 3433 3380
rect 3016 3340 3022 3352
rect 3421 3349 3433 3352
rect 3467 3380 3479 3383
rect 3510 3380 3516 3392
rect 3467 3352 3516 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 7392 3380 7420 3420
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8404 3448 8432 3479
rect 8662 3476 8668 3488
rect 8720 3516 8726 3528
rect 9223 3516 9251 3556
rect 8720 3488 9251 3516
rect 9309 3519 9367 3525
rect 8720 3476 8726 3488
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9416 3516 9444 3556
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9640 3556 9689 3584
rect 9640 3544 9646 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 9766 3544 9772 3596
rect 9824 3544 9830 3596
rect 9944 3587 10002 3593
rect 9944 3553 9956 3587
rect 9990 3584 10002 3587
rect 10318 3584 10324 3596
rect 9990 3556 10324 3584
rect 9990 3553 10002 3556
rect 9944 3547 10002 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 11112 3556 11161 3584
rect 11112 3544 11118 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 11992 3584 12020 3615
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 13081 3655 13139 3661
rect 13081 3652 13093 3655
rect 12768 3624 13093 3652
rect 12768 3612 12774 3624
rect 13081 3621 13093 3624
rect 13127 3621 13139 3655
rect 13538 3652 13544 3664
rect 13081 3615 13139 3621
rect 13188 3624 13544 3652
rect 13188 3584 13216 3624
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13722 3661 13728 3664
rect 13716 3652 13728 3661
rect 13683 3624 13728 3652
rect 13716 3615 13728 3624
rect 13722 3612 13728 3615
rect 13780 3612 13786 3664
rect 14844 3584 14872 3683
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 17589 3723 17647 3729
rect 17589 3689 17601 3723
rect 17635 3689 17647 3723
rect 17589 3683 17647 3689
rect 18417 3723 18475 3729
rect 18417 3689 18429 3723
rect 18463 3720 18475 3723
rect 19705 3723 19763 3729
rect 19705 3720 19717 3723
rect 18463 3692 19717 3720
rect 18463 3689 18475 3692
rect 18417 3683 18475 3689
rect 19705 3689 19717 3692
rect 19751 3689 19763 3723
rect 19705 3683 19763 3689
rect 15838 3652 15844 3664
rect 15799 3624 15844 3652
rect 15838 3612 15844 3624
rect 15896 3612 15902 3664
rect 15933 3655 15991 3661
rect 15933 3621 15945 3655
rect 15979 3652 15991 3655
rect 16114 3652 16120 3664
rect 15979 3624 16120 3652
rect 15979 3621 15991 3624
rect 15933 3615 15991 3621
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 16482 3612 16488 3664
rect 16540 3652 16546 3664
rect 17129 3655 17187 3661
rect 17129 3652 17141 3655
rect 16540 3624 17141 3652
rect 16540 3612 16546 3624
rect 17129 3621 17141 3624
rect 17175 3621 17187 3655
rect 17129 3615 17187 3621
rect 17218 3612 17224 3664
rect 17276 3652 17282 3664
rect 17604 3652 17632 3683
rect 18785 3655 18843 3661
rect 18785 3652 18797 3655
rect 17276 3624 17321 3652
rect 17604 3624 18797 3652
rect 17276 3612 17282 3624
rect 18785 3621 18797 3624
rect 18831 3621 18843 3655
rect 18785 3615 18843 3621
rect 19518 3612 19524 3664
rect 19576 3652 19582 3664
rect 19613 3655 19671 3661
rect 19613 3652 19625 3655
rect 19576 3624 19625 3652
rect 19576 3612 19582 3624
rect 19613 3621 19625 3624
rect 19659 3621 19671 3655
rect 19613 3615 19671 3621
rect 11992 3556 13216 3584
rect 13280 3556 14872 3584
rect 15856 3584 15884 3612
rect 16301 3587 16359 3593
rect 16301 3584 16313 3587
rect 15856 3556 16313 3584
rect 11149 3547 11207 3553
rect 9784 3516 9812 3544
rect 13280 3528 13308 3556
rect 16301 3553 16313 3556
rect 16347 3553 16359 3587
rect 17954 3584 17960 3596
rect 17915 3556 17960 3584
rect 16301 3547 16359 3553
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18506 3584 18512 3596
rect 18095 3556 18512 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 12158 3516 12164 3528
rect 9416 3488 9812 3516
rect 12071 3488 12164 3516
rect 9309 3479 9367 3485
rect 8570 3448 8576 3460
rect 8404 3420 8576 3448
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 9324 3448 9352 3479
rect 12158 3476 12164 3488
rect 12216 3516 12222 3528
rect 13078 3516 13084 3528
rect 12216 3488 13084 3516
rect 12216 3476 12222 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13262 3516 13268 3528
rect 13175 3488 13268 3516
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16574 3516 16580 3528
rect 16163 3488 16580 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 8680 3420 9352 3448
rect 4203 3352 7420 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 7616 3352 7849 3380
rect 7616 3340 7622 3352
rect 7837 3349 7849 3352
rect 7883 3380 7895 3383
rect 8680 3380 8708 3420
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13170 3448 13176 3460
rect 12492 3420 13176 3448
rect 12492 3408 12498 3420
rect 13170 3408 13176 3420
rect 13228 3448 13234 3460
rect 13464 3448 13492 3479
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17126 3516 17132 3528
rect 16908 3488 17132 3516
rect 16908 3476 16914 3488
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17310 3476 17316 3528
rect 17368 3516 17374 3528
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17368 3488 18153 3516
rect 17368 3476 17374 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3485 18935 3519
rect 18877 3479 18935 3485
rect 13228 3420 13492 3448
rect 13228 3408 13234 3420
rect 16390 3408 16396 3460
rect 16448 3448 16454 3460
rect 18892 3448 18920 3479
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19024 3488 19069 3516
rect 19024 3476 19030 3488
rect 19702 3476 19708 3528
rect 19760 3516 19766 3528
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 19760 3488 19809 3516
rect 19760 3476 19766 3488
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 16448 3420 18920 3448
rect 19245 3451 19303 3457
rect 16448 3408 16454 3420
rect 19245 3417 19257 3451
rect 19291 3448 19303 3451
rect 20530 3448 20536 3460
rect 19291 3420 20536 3448
rect 19291 3417 19303 3420
rect 19245 3411 19303 3417
rect 20530 3408 20536 3420
rect 20588 3408 20594 3460
rect 7883 3352 8708 3380
rect 8757 3383 8815 3389
rect 7883 3349 7895 3352
rect 7837 3343 7895 3349
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 10870 3380 10876 3392
rect 8803 3352 10876 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 11333 3383 11391 3389
rect 11333 3349 11345 3383
rect 11379 3380 11391 3383
rect 11698 3380 11704 3392
rect 11379 3352 11704 3380
rect 11379 3349 11391 3352
rect 11333 3343 11391 3349
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 12621 3383 12679 3389
rect 12621 3380 12633 3383
rect 11848 3352 12633 3380
rect 11848 3340 11854 3352
rect 12621 3349 12633 3352
rect 12667 3349 12679 3383
rect 12621 3343 12679 3349
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 16485 3383 16543 3389
rect 16485 3380 16497 3383
rect 16356 3352 16497 3380
rect 16356 3340 16362 3352
rect 16485 3349 16497 3352
rect 16531 3349 16543 3383
rect 16485 3343 16543 3349
rect 16761 3383 16819 3389
rect 16761 3349 16773 3383
rect 16807 3380 16819 3383
rect 18598 3380 18604 3392
rect 16807 3352 18604 3380
rect 16807 3349 16819 3352
rect 16761 3343 16819 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 2004 3148 2237 3176
rect 2004 3136 2010 3148
rect 2225 3145 2237 3148
rect 2271 3145 2283 3179
rect 3694 3176 3700 3188
rect 2225 3139 2283 3145
rect 2700 3148 3700 3176
rect 566 3068 572 3120
rect 624 3108 630 3120
rect 2590 3108 2596 3120
rect 624 3080 2596 3108
rect 624 3068 630 3080
rect 2590 3068 2596 3080
rect 2648 3068 2654 3120
rect 2700 3049 2728 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 4764 3148 6132 3176
rect 4764 3136 4770 3148
rect 4433 3111 4491 3117
rect 4433 3077 4445 3111
rect 4479 3108 4491 3111
rect 4798 3108 4804 3120
rect 4479 3080 4804 3108
rect 4479 3077 4491 3080
rect 4433 3071 4491 3077
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 6104 3108 6132 3148
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 6273 3179 6331 3185
rect 6273 3176 6285 3179
rect 6236 3148 6285 3176
rect 6236 3136 6242 3148
rect 6273 3145 6285 3148
rect 6319 3145 6331 3179
rect 6273 3139 6331 3145
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 6604 3148 8432 3176
rect 6604 3136 6610 3148
rect 6454 3108 6460 3120
rect 6104 3080 6460 3108
rect 6454 3068 6460 3080
rect 6512 3068 6518 3120
rect 8404 3108 8432 3148
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 9582 3176 9588 3188
rect 8628 3148 9588 3176
rect 8628 3136 8634 3148
rect 9582 3136 9588 3148
rect 9640 3176 9646 3188
rect 10318 3176 10324 3188
rect 9640 3148 10180 3176
rect 10279 3148 10324 3176
rect 9640 3136 9646 3148
rect 8938 3108 8944 3120
rect 8404 3080 8944 3108
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 10152 3108 10180 3148
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13136 3148 13829 3176
rect 13136 3136 13142 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 13817 3139 13875 3145
rect 15013 3179 15071 3185
rect 15013 3145 15025 3179
rect 15059 3176 15071 3179
rect 17218 3176 17224 3188
rect 15059 3148 17224 3176
rect 15059 3145 15071 3148
rect 15013 3139 15071 3145
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17368 3148 17413 3176
rect 17368 3136 17374 3148
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 18012 3148 18061 3176
rect 18012 3136 18018 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 10152 3080 11928 3108
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 2958 3040 2964 3052
rect 2915 3012 2964 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10192 3012 10977 3040
rect 10192 3000 10198 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 2038 2932 2044 2984
rect 2096 2972 2102 2984
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 2096 2944 2605 2972
rect 2096 2932 2102 2944
rect 2593 2941 2605 2944
rect 2639 2941 2651 2975
rect 2593 2935 2651 2941
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2972 3111 2975
rect 4706 2972 4712 2984
rect 3099 2944 4712 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 4706 2932 4712 2944
rect 4764 2972 4770 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4764 2944 4905 2972
rect 4764 2932 4770 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 5994 2972 6000 2984
rect 5776 2944 6000 2972
rect 5776 2932 5782 2944
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7736 2975 7794 2981
rect 7736 2941 7748 2975
rect 7782 2972 7794 2975
rect 8662 2972 8668 2984
rect 7782 2944 8668 2972
rect 7782 2941 7794 2944
rect 7736 2935 7794 2941
rect 934 2864 940 2916
rect 992 2904 998 2916
rect 2958 2904 2964 2916
rect 992 2876 2964 2904
rect 992 2864 998 2876
rect 2958 2864 2964 2876
rect 3016 2864 3022 2916
rect 3142 2864 3148 2916
rect 3200 2904 3206 2916
rect 3298 2907 3356 2913
rect 3298 2904 3310 2907
rect 3200 2876 3310 2904
rect 3200 2864 3206 2876
rect 3298 2873 3310 2876
rect 3344 2873 3356 2907
rect 3298 2867 3356 2873
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 5166 2913 5172 2916
rect 5160 2904 5172 2913
rect 4028 2876 5028 2904
rect 5127 2876 5172 2904
rect 4028 2864 4034 2876
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 4890 2836 4896 2848
rect 256 2808 4896 2836
rect 256 2796 262 2808
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5000 2836 5028 2876
rect 5160 2867 5172 2876
rect 5166 2864 5172 2867
rect 5224 2864 5230 2916
rect 7484 2904 7512 2935
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 8941 2975 8999 2981
rect 8941 2972 8953 2975
rect 8904 2944 8953 2972
rect 8904 2932 8910 2944
rect 8941 2941 8953 2944
rect 8987 2941 8999 2975
rect 8941 2935 8999 2941
rect 9208 2975 9266 2981
rect 9208 2941 9220 2975
rect 9254 2972 9266 2975
rect 10152 2972 10180 3000
rect 9254 2944 10180 2972
rect 9254 2941 9266 2944
rect 9208 2935 9266 2941
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10928 2944 11253 2972
rect 10928 2932 10934 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11790 2972 11796 2984
rect 11751 2944 11796 2972
rect 11241 2935 11299 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 11900 2972 11928 3080
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 13780 3080 14105 3108
rect 13780 3068 13786 3080
rect 14093 3077 14105 3080
rect 14139 3077 14151 3111
rect 14093 3071 14151 3077
rect 16942 3068 16948 3120
rect 17000 3108 17006 3120
rect 17589 3111 17647 3117
rect 17589 3108 17601 3111
rect 17000 3080 17601 3108
rect 17000 3068 17006 3080
rect 17589 3077 17601 3080
rect 17635 3077 17647 3111
rect 17589 3071 17647 3077
rect 12434 3040 12440 3052
rect 12395 3012 12440 3040
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 15473 3043 15531 3049
rect 13688 3012 14412 3040
rect 13688 3000 13694 3012
rect 11900 2944 13391 2972
rect 8864 2904 8892 2932
rect 10686 2904 10692 2916
rect 7484 2876 8892 2904
rect 10336 2876 10692 2904
rect 7742 2836 7748 2848
rect 5000 2808 7748 2836
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 8846 2836 8852 2848
rect 8536 2808 8852 2836
rect 8536 2796 8542 2808
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 10336 2836 10364 2876
rect 10686 2864 10692 2876
rect 10744 2864 10750 2916
rect 10781 2907 10839 2913
rect 10781 2873 10793 2907
rect 10827 2904 10839 2907
rect 10962 2904 10968 2916
rect 10827 2876 10968 2904
rect 10827 2873 10839 2876
rect 10781 2867 10839 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 11517 2907 11575 2913
rect 11517 2873 11529 2907
rect 11563 2873 11575 2907
rect 11517 2867 11575 2873
rect 8996 2808 10364 2836
rect 8996 2796 9002 2808
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 10873 2839 10931 2845
rect 10468 2808 10513 2836
rect 10468 2796 10474 2808
rect 10873 2805 10885 2839
rect 10919 2836 10931 2839
rect 11146 2836 11152 2848
rect 10919 2808 11152 2836
rect 10919 2805 10931 2808
rect 10873 2799 10931 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11532 2836 11560 2867
rect 11882 2864 11888 2916
rect 11940 2904 11946 2916
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 11940 2876 12081 2904
rect 11940 2864 11946 2876
rect 12069 2873 12081 2876
rect 12115 2873 12127 2907
rect 12069 2867 12127 2873
rect 12704 2907 12762 2913
rect 12704 2873 12716 2907
rect 12750 2904 12762 2907
rect 13262 2904 13268 2916
rect 12750 2876 13268 2904
rect 12750 2873 12762 2876
rect 12704 2867 12762 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 13078 2836 13084 2848
rect 11532 2808 13084 2836
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 13363 2836 13391 2944
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 14384 2981 14412 3012
rect 15473 3009 15485 3043
rect 15519 3040 15531 3043
rect 15562 3040 15568 3052
rect 15519 3012 15568 3040
rect 15519 3009 15531 3012
rect 15473 3003 15531 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 15657 3043 15715 3049
rect 15657 3009 15669 3043
rect 15703 3009 15715 3043
rect 15930 3040 15936 3052
rect 15891 3012 15936 3040
rect 15657 3003 15715 3009
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 13596 2944 13921 2972
rect 13596 2932 13602 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2941 14427 2975
rect 15672 2972 15700 3003
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 17144 3012 18613 3040
rect 15672 2944 15976 2972
rect 14369 2935 14427 2941
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 15838 2904 15844 2916
rect 14691 2876 15844 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15838 2864 15844 2876
rect 15896 2864 15902 2916
rect 15948 2904 15976 2944
rect 16022 2932 16028 2984
rect 16080 2972 16086 2984
rect 16758 2972 16764 2984
rect 16080 2944 16764 2972
rect 16080 2932 16086 2944
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 16200 2907 16258 2913
rect 16200 2904 16212 2907
rect 15948 2876 16212 2904
rect 16200 2873 16212 2876
rect 16246 2904 16258 2907
rect 16574 2904 16580 2916
rect 16246 2876 16580 2904
rect 16246 2873 16258 2876
rect 16200 2867 16258 2873
rect 16574 2864 16580 2876
rect 16632 2904 16638 2916
rect 17144 2904 17172 3012
rect 18601 3009 18613 3012
rect 18647 3040 18659 3043
rect 18966 3040 18972 3052
rect 18647 3012 18972 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 17402 2972 17408 2984
rect 17363 2944 17408 2972
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 18414 2972 18420 2984
rect 18375 2944 18420 2972
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 18748 2944 18889 2972
rect 18748 2932 18754 2944
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 16632 2876 17172 2904
rect 16632 2864 16638 2876
rect 17954 2864 17960 2916
rect 18012 2904 18018 2916
rect 18012 2876 19104 2904
rect 18012 2864 18018 2876
rect 15381 2839 15439 2845
rect 15381 2836 15393 2839
rect 13363 2808 15393 2836
rect 15381 2805 15393 2808
rect 15427 2805 15439 2839
rect 15381 2799 15439 2805
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 16482 2836 16488 2848
rect 15712 2808 16488 2836
rect 15712 2796 15718 2808
rect 16482 2796 16488 2808
rect 16540 2796 16546 2848
rect 18509 2839 18567 2845
rect 18509 2805 18521 2839
rect 18555 2836 18567 2839
rect 18598 2836 18604 2848
rect 18555 2808 18604 2836
rect 18555 2805 18567 2808
rect 18509 2799 18567 2805
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 19076 2845 19104 2876
rect 19061 2839 19119 2845
rect 19061 2805 19073 2839
rect 19107 2805 19119 2839
rect 19061 2799 19119 2805
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 2924 2604 3157 2632
rect 2924 2592 2930 2604
rect 3145 2601 3157 2604
rect 3191 2601 3203 2635
rect 3145 2595 3203 2601
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 5350 2632 5356 2644
rect 4948 2604 5212 2632
rect 5311 2604 5356 2632
rect 4948 2592 4954 2604
rect 3605 2567 3663 2573
rect 3605 2533 3617 2567
rect 3651 2564 3663 2567
rect 4062 2564 4068 2576
rect 3651 2536 4068 2564
rect 3651 2533 3663 2536
rect 3605 2527 3663 2533
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 5074 2564 5080 2576
rect 5000 2536 5080 2564
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 3384 2468 3525 2496
rect 3384 2456 3390 2468
rect 3513 2465 3525 2468
rect 3559 2496 3571 2499
rect 3878 2496 3884 2508
rect 3559 2468 3884 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4890 2496 4896 2508
rect 4851 2468 4896 2496
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 5000 2437 5028 2536
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5184 2564 5212 2604
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 6454 2632 6460 2644
rect 5684 2604 6460 2632
rect 5684 2592 5690 2604
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7432 2604 7481 2632
rect 7432 2592 7438 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 7469 2595 7527 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 8757 2635 8815 2641
rect 8757 2632 8769 2635
rect 8628 2604 8769 2632
rect 8628 2592 8634 2604
rect 8757 2601 8769 2604
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2601 9827 2635
rect 9769 2595 9827 2601
rect 7558 2564 7564 2576
rect 5184 2536 7564 2564
rect 7558 2524 7564 2536
rect 7616 2564 7622 2576
rect 7929 2567 7987 2573
rect 7929 2564 7941 2567
rect 7616 2536 7941 2564
rect 7616 2524 7622 2536
rect 7929 2533 7941 2536
rect 7975 2533 7987 2567
rect 8662 2564 8668 2576
rect 8623 2536 8668 2564
rect 7929 2527 7987 2533
rect 8662 2524 8668 2536
rect 8720 2564 8726 2576
rect 9490 2564 9496 2576
rect 8720 2536 9496 2564
rect 8720 2524 8726 2536
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5684 2468 5733 2496
rect 5684 2456 5690 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 5868 2468 5913 2496
rect 5868 2456 5874 2468
rect 7742 2456 7748 2508
rect 7800 2496 7806 2508
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7800 2468 7849 2496
rect 7800 2456 7806 2468
rect 7837 2465 7849 2468
rect 7883 2496 7895 2499
rect 9674 2496 9680 2508
rect 7883 2468 9680 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 9784 2496 9812 2595
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 10100 2604 10149 2632
rect 10100 2592 10106 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10137 2595 10195 2601
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10410 2632 10416 2644
rect 10275 2604 10416 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 12952 2604 13860 2632
rect 12952 2592 12958 2604
rect 10873 2567 10931 2573
rect 10873 2533 10885 2567
rect 10919 2564 10931 2567
rect 11054 2564 11060 2576
rect 10919 2536 11060 2564
rect 10919 2533 10931 2536
rect 10873 2527 10931 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11425 2567 11483 2573
rect 11425 2533 11437 2567
rect 11471 2564 11483 2567
rect 13446 2564 13452 2576
rect 11471 2536 13452 2564
rect 11471 2533 11483 2536
rect 11425 2527 11483 2533
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 13832 2564 13860 2604
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14056 2604 14841 2632
rect 14056 2592 14062 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 16393 2635 16451 2641
rect 16393 2601 16405 2635
rect 16439 2601 16451 2635
rect 16393 2595 16451 2601
rect 13832 2536 14044 2564
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 9784 2468 10609 2496
rect 10597 2465 10609 2468
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2465 11207 2499
rect 11882 2496 11888 2508
rect 11843 2468 11888 2496
rect 11149 2459 11207 2465
rect 3697 2431 3755 2437
rect 3697 2428 3709 2431
rect 3660 2400 3709 2428
rect 3660 2388 3666 2400
rect 3697 2397 3709 2400
rect 3743 2397 3755 2431
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 3697 2391 3755 2397
rect 4264 2400 4997 2428
rect 2406 2320 2412 2372
rect 2464 2360 2470 2372
rect 4264 2360 4292 2400
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2428 5230 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5224 2400 5917 2428
rect 5224 2388 5230 2400
rect 5905 2397 5917 2400
rect 5951 2428 5963 2431
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 5951 2400 8033 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 8021 2397 8033 2400
rect 8067 2428 8079 2431
rect 8846 2428 8852 2440
rect 8067 2400 8852 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 2464 2332 4292 2360
rect 4525 2363 4583 2369
rect 2464 2320 2470 2332
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 5534 2360 5540 2372
rect 4571 2332 5540 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 5534 2320 5540 2332
rect 5592 2320 5598 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 11164 2360 11192 2459
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12667 2468 13032 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12894 2428 12900 2440
rect 12855 2400 12900 2428
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13004 2428 13032 2468
rect 13078 2456 13084 2508
rect 13136 2496 13142 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 13136 2468 13185 2496
rect 13136 2456 13142 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 13566 2499 13624 2505
rect 13566 2465 13578 2499
rect 13612 2496 13624 2499
rect 13814 2496 13820 2508
rect 13612 2468 13820 2496
rect 13612 2465 13624 2468
rect 13566 2459 13624 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 13354 2428 13360 2440
rect 13004 2400 13360 2428
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13446 2388 13452 2440
rect 13504 2428 13510 2440
rect 13924 2428 13952 2459
rect 13504 2400 13952 2428
rect 14016 2428 14044 2536
rect 14734 2524 14740 2576
rect 14792 2564 14798 2576
rect 16408 2564 16436 2595
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 17129 2635 17187 2641
rect 17129 2632 17141 2635
rect 16540 2604 17141 2632
rect 16540 2592 16546 2604
rect 17129 2601 17141 2604
rect 17175 2601 17187 2635
rect 17129 2595 17187 2601
rect 18325 2635 18383 2641
rect 18325 2601 18337 2635
rect 18371 2632 18383 2635
rect 18506 2632 18512 2644
rect 18371 2604 18512 2632
rect 18371 2601 18383 2604
rect 18325 2595 18383 2601
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 18782 2632 18788 2644
rect 18743 2604 18788 2632
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 14792 2536 16436 2564
rect 14792 2524 14798 2536
rect 16758 2524 16764 2576
rect 16816 2564 16822 2576
rect 16816 2536 17356 2564
rect 16816 2524 16822 2536
rect 14274 2496 14280 2508
rect 14235 2468 14280 2496
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14516 2468 14657 2496
rect 14516 2456 14522 2468
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 15013 2499 15071 2505
rect 15013 2465 15025 2499
rect 15059 2465 15071 2499
rect 15013 2459 15071 2465
rect 15028 2428 15056 2459
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 15657 2499 15715 2505
rect 15657 2496 15669 2499
rect 15528 2468 15669 2496
rect 15528 2456 15534 2468
rect 15657 2465 15669 2468
rect 15703 2465 15715 2499
rect 15657 2459 15715 2465
rect 15746 2456 15752 2508
rect 15804 2496 15810 2508
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 15804 2468 16221 2496
rect 15804 2456 15810 2468
rect 16209 2465 16221 2468
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2496 16635 2499
rect 16850 2496 16856 2508
rect 16623 2468 16856 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17034 2496 17040 2508
rect 16991 2468 17040 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 17328 2505 17356 2536
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 19720 2564 19748 2595
rect 17828 2536 19748 2564
rect 17828 2524 17834 2536
rect 17313 2499 17371 2505
rect 17313 2465 17325 2499
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17586 2456 17592 2508
rect 17644 2496 17650 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17644 2468 17693 2496
rect 17644 2456 17650 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 18690 2496 18696 2508
rect 18651 2468 18696 2496
rect 17681 2459 17739 2465
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 19153 2499 19211 2505
rect 19153 2496 19165 2499
rect 18800 2468 19165 2496
rect 14016 2400 15056 2428
rect 15933 2431 15991 2437
rect 13504 2388 13510 2400
rect 15933 2397 15945 2431
rect 15979 2428 15991 2431
rect 18800 2428 18828 2468
rect 19153 2465 19165 2468
rect 19199 2465 19211 2499
rect 19153 2459 19211 2465
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19521 2499 19579 2505
rect 19521 2496 19533 2499
rect 19392 2468 19533 2496
rect 19392 2456 19398 2468
rect 19521 2465 19533 2468
rect 19567 2465 19579 2499
rect 19521 2459 19579 2465
rect 19794 2456 19800 2508
rect 19852 2496 19858 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19852 2468 19901 2496
rect 19852 2456 19858 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 18966 2428 18972 2440
rect 15979 2400 18828 2428
rect 18927 2400 18972 2428
rect 15979 2397 15991 2400
rect 15933 2391 15991 2397
rect 18966 2388 18972 2400
rect 19024 2388 19030 2440
rect 8444 2332 11192 2360
rect 8444 2320 8450 2332
rect 12526 2320 12532 2372
rect 12584 2360 12590 2372
rect 12584 2332 13492 2360
rect 12584 2320 12590 2332
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 6638 2292 6644 2304
rect 3936 2264 6644 2292
rect 3936 2252 3942 2264
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 9398 2292 9404 2304
rect 8076 2264 9404 2292
rect 8076 2252 8082 2264
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 12069 2295 12127 2301
rect 12069 2292 12081 2295
rect 11664 2264 12081 2292
rect 11664 2252 11670 2264
rect 12069 2261 12081 2264
rect 12115 2261 12127 2295
rect 12069 2255 12127 2261
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 12216 2264 13369 2292
rect 12216 2252 12222 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13464 2292 13492 2332
rect 13630 2320 13636 2372
rect 13688 2360 13694 2372
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 13688 2332 14473 2360
rect 13688 2320 13694 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 14461 2323 14519 2329
rect 15102 2320 15108 2372
rect 15160 2360 15166 2372
rect 15160 2332 16528 2360
rect 15160 2320 15166 2332
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 13464 2264 13737 2292
rect 13357 2255 13415 2261
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 14090 2292 14096 2304
rect 14051 2264 14096 2292
rect 13725 2255 13783 2261
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 14366 2252 14372 2304
rect 14424 2292 14430 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 14424 2264 15209 2292
rect 14424 2252 14430 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 16500 2292 16528 2332
rect 16574 2320 16580 2372
rect 16632 2360 16638 2372
rect 17865 2363 17923 2369
rect 17865 2360 17877 2363
rect 16632 2332 17877 2360
rect 16632 2320 16638 2332
rect 17865 2329 17877 2332
rect 17911 2329 17923 2363
rect 17865 2323 17923 2329
rect 18506 2320 18512 2372
rect 18564 2360 18570 2372
rect 20073 2363 20131 2369
rect 20073 2360 20085 2363
rect 18564 2332 20085 2360
rect 18564 2320 18570 2332
rect 20073 2329 20085 2332
rect 20119 2329 20131 2363
rect 20073 2323 20131 2329
rect 16761 2295 16819 2301
rect 16761 2292 16773 2295
rect 16500 2264 16773 2292
rect 15197 2255 15255 2261
rect 16761 2261 16773 2264
rect 16807 2261 16819 2295
rect 17494 2292 17500 2304
rect 17455 2264 17500 2292
rect 16761 2255 16819 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 17586 2252 17592 2304
rect 17644 2292 17650 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 17644 2264 19349 2292
rect 17644 2252 17650 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2038 2048 2044 2100
rect 2096 2088 2102 2100
rect 2096 2060 3648 2088
rect 2096 2048 2102 2060
rect 3620 1952 3648 2060
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 8202 2088 8208 2100
rect 4120 2060 8208 2088
rect 4120 2048 4126 2060
rect 8202 2048 8208 2060
rect 8260 2048 8266 2100
rect 6546 1980 6552 2032
rect 6604 2020 6610 2032
rect 9306 2020 9312 2032
rect 6604 1992 9312 2020
rect 6604 1980 6610 1992
rect 9306 1980 9312 1992
rect 9364 1980 9370 2032
rect 5626 1952 5632 1964
rect 3620 1924 5632 1952
rect 5626 1912 5632 1924
rect 5684 1912 5690 1964
rect 1302 1776 1308 1828
rect 1360 1816 1366 1828
rect 8662 1816 8668 1828
rect 1360 1788 8668 1816
rect 1360 1776 1366 1788
rect 8662 1776 8668 1788
rect 8720 1776 8726 1828
rect 1670 1708 1676 1760
rect 1728 1748 1734 1760
rect 5810 1748 5816 1760
rect 1728 1720 5816 1748
rect 1728 1708 1734 1720
rect 5810 1708 5816 1720
rect 5868 1708 5874 1760
rect 13262 1436 13268 1488
rect 13320 1476 13326 1488
rect 13722 1476 13728 1488
rect 13320 1448 13728 1476
rect 13320 1436 13326 1448
rect 13722 1436 13728 1448
rect 13780 1436 13786 1488
rect 8386 1368 8392 1420
rect 8444 1408 8450 1420
rect 9214 1408 9220 1420
rect 8444 1380 9220 1408
rect 8444 1368 8450 1380
rect 9214 1368 9220 1380
rect 9272 1368 9278 1420
rect 9950 1368 9956 1420
rect 10008 1408 10014 1420
rect 10594 1408 10600 1420
rect 10008 1380 10600 1408
rect 10008 1368 10014 1380
rect 10594 1368 10600 1380
rect 10652 1368 10658 1420
rect 12894 1368 12900 1420
rect 12952 1408 12958 1420
rect 14090 1408 14096 1420
rect 12952 1380 14096 1408
rect 12952 1368 12958 1380
rect 14090 1368 14096 1380
rect 14148 1368 14154 1420
rect 15838 1368 15844 1420
rect 15896 1408 15902 1420
rect 17494 1408 17500 1420
rect 15896 1380 17500 1408
rect 15896 1368 15902 1380
rect 17494 1368 17500 1380
rect 17552 1368 17558 1420
rect 20714 892 20720 944
rect 20772 932 20778 944
rect 21542 932 21548 944
rect 20772 904 21548 932
rect 20772 892 20778 904
rect 21542 892 21548 904
rect 21600 892 21606 944
<< via1 >>
rect 7012 20544 7064 20596
rect 7564 20544 7616 20596
rect 4344 20340 4396 20392
rect 9036 20340 9088 20392
rect 7104 20272 7156 20324
rect 8116 20272 8168 20324
rect 4068 20204 4120 20256
rect 15200 20204 15252 20256
rect 19340 20204 19392 20256
rect 20628 20204 20680 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 4804 20000 4856 20052
rect 9772 20000 9824 20052
rect 13820 20000 13872 20052
rect 15752 20000 15804 20052
rect 16120 20000 16172 20052
rect 5172 19932 5224 19984
rect 10140 19932 10192 19984
rect 22192 20000 22244 20052
rect 5540 19864 5592 19916
rect 6828 19864 6880 19916
rect 7288 19864 7340 19916
rect 8208 19864 8260 19916
rect 13268 19907 13320 19916
rect 13268 19873 13277 19907
rect 13277 19873 13311 19907
rect 13311 19873 13320 19907
rect 13268 19864 13320 19873
rect 15844 19907 15896 19916
rect 4252 19839 4304 19848
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 7748 19796 7800 19848
rect 15844 19873 15853 19907
rect 15853 19873 15887 19907
rect 15887 19873 15896 19907
rect 15844 19864 15896 19873
rect 21456 19932 21508 19984
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 19524 19864 19576 19916
rect 19800 19864 19852 19916
rect 20444 19907 20496 19916
rect 16304 19796 16356 19848
rect 11612 19728 11664 19780
rect 5632 19703 5684 19712
rect 5632 19669 5641 19703
rect 5641 19669 5675 19703
rect 5675 19669 5684 19703
rect 5632 19660 5684 19669
rect 5816 19660 5868 19712
rect 9772 19660 9824 19712
rect 19156 19796 19208 19848
rect 20444 19873 20453 19907
rect 20453 19873 20487 19907
rect 20487 19873 20496 19907
rect 20444 19864 20496 19873
rect 21824 19796 21876 19848
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 4252 19456 4304 19508
rect 204 19252 256 19304
rect 4252 19320 4304 19372
rect 4620 19388 4672 19440
rect 5540 19456 5592 19508
rect 9680 19388 9732 19440
rect 9220 19363 9272 19372
rect 572 19184 624 19236
rect 4160 19184 4212 19236
rect 4804 19252 4856 19304
rect 4988 19252 5040 19304
rect 2964 19116 3016 19168
rect 3424 19116 3476 19168
rect 4068 19159 4120 19168
rect 4068 19125 4077 19159
rect 4077 19125 4111 19159
rect 4111 19125 4120 19159
rect 4068 19116 4120 19125
rect 4620 19116 4672 19168
rect 4988 19116 5040 19168
rect 6092 19184 6144 19236
rect 5264 19116 5316 19168
rect 5448 19116 5500 19168
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 9956 19252 10008 19304
rect 10140 19295 10192 19304
rect 10140 19261 10149 19295
rect 10149 19261 10183 19295
rect 10183 19261 10192 19295
rect 10140 19252 10192 19261
rect 13268 19320 13320 19372
rect 15200 19320 15252 19372
rect 10876 19252 10928 19304
rect 11888 19252 11940 19304
rect 12992 19252 13044 19304
rect 13452 19295 13504 19304
rect 8668 19184 8720 19236
rect 8760 19184 8812 19236
rect 7656 19116 7708 19168
rect 7748 19116 7800 19168
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 9128 19116 9180 19168
rect 9496 19116 9548 19168
rect 10784 19184 10836 19236
rect 11152 19116 11204 19168
rect 12348 19184 12400 19236
rect 12808 19184 12860 19236
rect 13452 19261 13461 19295
rect 13461 19261 13495 19295
rect 13495 19261 13504 19295
rect 13452 19252 13504 19261
rect 13820 19295 13872 19304
rect 13820 19261 13829 19295
rect 13829 19261 13863 19295
rect 13863 19261 13872 19295
rect 13820 19252 13872 19261
rect 13912 19252 13964 19304
rect 14372 19252 14424 19304
rect 13176 19184 13228 19236
rect 11980 19159 12032 19168
rect 11980 19125 11989 19159
rect 11989 19125 12023 19159
rect 12023 19125 12032 19159
rect 11980 19116 12032 19125
rect 12716 19116 12768 19168
rect 13544 19184 13596 19236
rect 14096 19184 14148 19236
rect 15108 19252 15160 19304
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 16488 19295 16540 19304
rect 16488 19261 16497 19295
rect 16497 19261 16531 19295
rect 16531 19261 16540 19295
rect 16488 19252 16540 19261
rect 16948 19252 17000 19304
rect 17684 19295 17736 19304
rect 17132 19227 17184 19236
rect 17132 19193 17141 19227
rect 17141 19193 17175 19227
rect 17175 19193 17184 19227
rect 17132 19184 17184 19193
rect 14188 19116 14240 19168
rect 14556 19116 14608 19168
rect 15016 19116 15068 19168
rect 15384 19116 15436 19168
rect 16856 19116 16908 19168
rect 17684 19261 17693 19295
rect 17693 19261 17727 19295
rect 17727 19261 17736 19295
rect 17684 19252 17736 19261
rect 18328 19295 18380 19304
rect 18328 19261 18337 19295
rect 18337 19261 18371 19295
rect 18371 19261 18380 19295
rect 18328 19252 18380 19261
rect 18788 19252 18840 19304
rect 19892 19252 19944 19304
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 20720 19295 20772 19304
rect 20720 19261 20729 19295
rect 20729 19261 20763 19295
rect 20763 19261 20772 19295
rect 20720 19252 20772 19261
rect 18604 19227 18656 19236
rect 18604 19193 18613 19227
rect 18613 19193 18647 19227
rect 18647 19193 18656 19227
rect 18604 19184 18656 19193
rect 19616 19184 19668 19236
rect 19340 19116 19392 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1676 18912 1728 18964
rect 3056 18912 3108 18964
rect 3240 18955 3292 18964
rect 3240 18921 3249 18955
rect 3249 18921 3283 18955
rect 3283 18921 3292 18955
rect 3240 18912 3292 18921
rect 940 18844 992 18896
rect 3792 18912 3844 18964
rect 4068 18912 4120 18964
rect 5448 18955 5500 18964
rect 5448 18921 5457 18955
rect 5457 18921 5491 18955
rect 5491 18921 5500 18955
rect 5448 18912 5500 18921
rect 5816 18955 5868 18964
rect 5816 18921 5825 18955
rect 5825 18921 5859 18955
rect 5859 18921 5868 18955
rect 5816 18912 5868 18921
rect 6000 18912 6052 18964
rect 9496 18912 9548 18964
rect 11704 18912 11756 18964
rect 3424 18844 3476 18896
rect 5172 18887 5224 18896
rect 2412 18776 2464 18828
rect 4068 18776 4120 18828
rect 5172 18853 5181 18887
rect 5181 18853 5215 18887
rect 5215 18853 5224 18887
rect 5172 18844 5224 18853
rect 5264 18844 5316 18896
rect 8760 18844 8812 18896
rect 8852 18844 8904 18896
rect 10876 18887 10928 18896
rect 2044 18708 2096 18760
rect 2872 18640 2924 18692
rect 3424 18708 3476 18760
rect 3792 18708 3844 18760
rect 4988 18776 5040 18828
rect 5356 18776 5408 18828
rect 7840 18776 7892 18828
rect 9220 18776 9272 18828
rect 10508 18776 10560 18828
rect 10876 18853 10885 18887
rect 10885 18853 10919 18887
rect 10919 18853 10928 18887
rect 10876 18844 10928 18853
rect 13452 18912 13504 18964
rect 17316 18912 17368 18964
rect 19156 18912 19208 18964
rect 10692 18776 10744 18828
rect 12164 18844 12216 18896
rect 13912 18844 13964 18896
rect 15108 18844 15160 18896
rect 16488 18844 16540 18896
rect 11612 18819 11664 18828
rect 11612 18785 11646 18819
rect 11646 18785 11664 18819
rect 11612 18776 11664 18785
rect 2780 18615 2832 18624
rect 2780 18581 2789 18615
rect 2789 18581 2823 18615
rect 2823 18581 2832 18615
rect 3240 18640 3292 18692
rect 3976 18640 4028 18692
rect 5264 18708 5316 18760
rect 5908 18751 5960 18760
rect 5908 18717 5917 18751
rect 5917 18717 5951 18751
rect 5951 18717 5960 18751
rect 5908 18708 5960 18717
rect 6092 18751 6144 18760
rect 6092 18717 6101 18751
rect 6101 18717 6135 18751
rect 6135 18717 6144 18751
rect 6092 18708 6144 18717
rect 7656 18708 7708 18760
rect 9588 18708 9640 18760
rect 4988 18640 5040 18692
rect 5632 18640 5684 18692
rect 2780 18572 2832 18581
rect 9220 18640 9272 18692
rect 8668 18572 8720 18624
rect 9404 18572 9456 18624
rect 10784 18572 10836 18624
rect 13820 18776 13872 18828
rect 14280 18819 14332 18828
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 15016 18776 15068 18828
rect 16764 18776 16816 18828
rect 18328 18776 18380 18828
rect 18144 18751 18196 18760
rect 18144 18717 18153 18751
rect 18153 18717 18187 18751
rect 18187 18717 18196 18751
rect 18144 18708 18196 18717
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 16948 18640 17000 18692
rect 19524 18912 19576 18964
rect 21088 18912 21140 18964
rect 20536 18887 20588 18896
rect 20536 18853 20545 18887
rect 20545 18853 20579 18887
rect 20579 18853 20588 18887
rect 20536 18844 20588 18853
rect 19432 18776 19484 18828
rect 19800 18776 19852 18828
rect 18972 18708 19024 18760
rect 19064 18640 19116 18692
rect 13452 18572 13504 18624
rect 13728 18572 13780 18624
rect 15936 18572 15988 18624
rect 20352 18572 20404 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18343 2004 18352
rect 1952 18309 1961 18343
rect 1961 18309 1995 18343
rect 1995 18309 2004 18343
rect 1952 18300 2004 18309
rect 2136 18232 2188 18284
rect 5908 18368 5960 18420
rect 11152 18368 11204 18420
rect 2872 18300 2924 18352
rect 4252 18300 4304 18352
rect 2872 18164 2924 18216
rect 4068 18232 4120 18284
rect 2412 18096 2464 18148
rect 2688 18096 2740 18148
rect 4436 18164 4488 18216
rect 3240 18139 3292 18148
rect 3240 18105 3274 18139
rect 3274 18105 3292 18139
rect 3240 18096 3292 18105
rect 3700 18096 3752 18148
rect 4712 18096 4764 18148
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 2872 18028 2924 18080
rect 3056 18028 3108 18080
rect 5724 18164 5776 18216
rect 6460 18232 6512 18284
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8576 18275 8628 18284
rect 8576 18241 8585 18275
rect 8585 18241 8619 18275
rect 8619 18241 8628 18275
rect 8576 18232 8628 18241
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 9864 18275 9916 18284
rect 8668 18232 8720 18241
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 11244 18300 11296 18352
rect 12992 18300 13044 18352
rect 13176 18368 13228 18420
rect 17592 18368 17644 18420
rect 9404 18164 9456 18216
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 9680 18164 9732 18216
rect 9772 18096 9824 18148
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 8760 18028 8812 18080
rect 11612 18232 11664 18284
rect 11060 18164 11112 18216
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 22560 18300 22612 18352
rect 20260 18232 20312 18284
rect 17500 18164 17552 18216
rect 19524 18164 19576 18216
rect 20352 18164 20404 18216
rect 20812 18232 20864 18284
rect 10968 18096 11020 18148
rect 12256 18096 12308 18148
rect 12992 18096 13044 18148
rect 19984 18096 20036 18148
rect 11428 18028 11480 18080
rect 11612 18071 11664 18080
rect 11612 18037 11621 18071
rect 11621 18037 11655 18071
rect 11655 18037 11664 18071
rect 11612 18028 11664 18037
rect 11796 18028 11848 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 4896 17824 4948 17876
rect 5448 17824 5500 17876
rect 7288 17824 7340 17876
rect 8208 17824 8260 17876
rect 11060 17824 11112 17876
rect 11152 17824 11204 17876
rect 11612 17824 11664 17876
rect 11888 17824 11940 17876
rect 12256 17824 12308 17876
rect 21088 17867 21140 17876
rect 21088 17833 21097 17867
rect 21097 17833 21131 17867
rect 21131 17833 21140 17867
rect 21088 17824 21140 17833
rect 2136 17799 2188 17808
rect 2136 17765 2170 17799
rect 2170 17765 2188 17799
rect 2136 17756 2188 17765
rect 2872 17756 2924 17808
rect 4068 17756 4120 17808
rect 4252 17756 4304 17808
rect 5264 17756 5316 17808
rect 9680 17756 9732 17808
rect 9864 17756 9916 17808
rect 11980 17756 12032 17808
rect 2412 17688 2464 17740
rect 2688 17688 2740 17740
rect 4068 17620 4120 17672
rect 4528 17663 4580 17672
rect 4528 17629 4537 17663
rect 4537 17629 4571 17663
rect 4571 17629 4580 17663
rect 4528 17620 4580 17629
rect 5540 17552 5592 17604
rect 6092 17552 6144 17604
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 5172 17484 5224 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 6000 17527 6052 17536
rect 6000 17493 6009 17527
rect 6009 17493 6043 17527
rect 6043 17493 6052 17527
rect 8116 17688 8168 17740
rect 8576 17688 8628 17740
rect 11152 17688 11204 17740
rect 12164 17731 12216 17740
rect 6460 17620 6512 17672
rect 7748 17620 7800 17672
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 11428 17620 11480 17672
rect 12164 17697 12173 17731
rect 12173 17697 12207 17731
rect 12207 17697 12216 17731
rect 12164 17688 12216 17697
rect 12348 17756 12400 17808
rect 18696 17756 18748 17808
rect 13728 17731 13780 17740
rect 11244 17552 11296 17604
rect 6000 17484 6052 17493
rect 8760 17484 8812 17536
rect 10876 17484 10928 17536
rect 10968 17484 11020 17536
rect 12072 17620 12124 17672
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 13728 17697 13762 17731
rect 13762 17697 13780 17731
rect 13728 17688 13780 17697
rect 19800 17688 19852 17740
rect 13452 17663 13504 17672
rect 13452 17629 13461 17663
rect 13461 17629 13495 17663
rect 13495 17629 13504 17663
rect 13452 17620 13504 17629
rect 21364 17620 21416 17672
rect 14556 17552 14608 17604
rect 20904 17552 20956 17604
rect 11888 17484 11940 17536
rect 12624 17527 12676 17536
rect 12624 17493 12633 17527
rect 12633 17493 12667 17527
rect 12667 17493 12676 17527
rect 12624 17484 12676 17493
rect 14464 17484 14516 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 4160 17280 4212 17332
rect 4804 17280 4856 17332
rect 6828 17323 6880 17332
rect 3332 17212 3384 17264
rect 3424 17212 3476 17264
rect 2228 17144 2280 17196
rect 3884 17212 3936 17264
rect 5264 17212 5316 17264
rect 5540 17212 5592 17264
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 8484 17280 8536 17332
rect 10692 17280 10744 17332
rect 10968 17323 11020 17332
rect 10968 17289 10977 17323
rect 10977 17289 11011 17323
rect 11011 17289 11020 17323
rect 10968 17280 11020 17289
rect 11796 17280 11848 17332
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 2780 17076 2832 17128
rect 3700 17144 3752 17196
rect 5172 17187 5224 17196
rect 5172 17153 5181 17187
rect 5181 17153 5215 17187
rect 5215 17153 5224 17187
rect 5172 17144 5224 17153
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 8944 17212 8996 17264
rect 9496 17212 9548 17264
rect 11520 17212 11572 17264
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 8116 17187 8168 17196
rect 8116 17153 8125 17187
rect 8125 17153 8159 17187
rect 8159 17153 8168 17187
rect 8116 17144 8168 17153
rect 9220 17144 9272 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 1860 16940 1912 16992
rect 2688 16940 2740 16992
rect 3056 17008 3108 17060
rect 4528 17008 4580 17060
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 3792 16983 3844 16992
rect 3792 16949 3801 16983
rect 3801 16949 3835 16983
rect 3835 16949 3844 16983
rect 3792 16940 3844 16949
rect 4252 16983 4304 16992
rect 4252 16949 4261 16983
rect 4261 16949 4295 16983
rect 4295 16949 4304 16983
rect 4252 16940 4304 16949
rect 4896 17076 4948 17128
rect 5632 17076 5684 17128
rect 9864 17119 9916 17128
rect 4712 17008 4764 17060
rect 6184 17008 6236 17060
rect 9864 17085 9898 17119
rect 9898 17085 9916 17119
rect 9864 17076 9916 17085
rect 11704 17076 11756 17128
rect 12992 17280 13044 17332
rect 15844 17280 15896 17332
rect 19892 17323 19944 17332
rect 19892 17289 19901 17323
rect 19901 17289 19935 17323
rect 19935 17289 19944 17323
rect 19892 17280 19944 17289
rect 20260 17323 20312 17332
rect 20260 17289 20269 17323
rect 20269 17289 20303 17323
rect 20303 17289 20312 17323
rect 20260 17280 20312 17289
rect 21180 17323 21232 17332
rect 21180 17289 21189 17323
rect 21189 17289 21223 17323
rect 21223 17289 21232 17323
rect 21180 17280 21232 17289
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 10508 17008 10560 17060
rect 6644 16940 6696 16992
rect 6920 16940 6972 16992
rect 8760 16983 8812 16992
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 8760 16940 8812 16949
rect 8944 16940 8996 16992
rect 11428 16940 11480 16992
rect 12532 17008 12584 17060
rect 12440 16940 12492 16992
rect 13268 17119 13320 17128
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 19432 17144 19484 17196
rect 14464 17008 14516 17060
rect 12900 16940 12952 16992
rect 14280 16940 14332 16992
rect 14556 16940 14608 16992
rect 16672 17076 16724 17128
rect 14832 17008 14884 17060
rect 19432 17008 19484 17060
rect 19800 17076 19852 17128
rect 20628 17076 20680 17128
rect 21272 17008 21324 17060
rect 15200 16940 15252 16992
rect 16120 16983 16172 16992
rect 16120 16949 16129 16983
rect 16129 16949 16163 16983
rect 16163 16949 16172 16983
rect 16120 16940 16172 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 1860 16736 1912 16788
rect 3608 16779 3660 16788
rect 3608 16745 3617 16779
rect 3617 16745 3651 16779
rect 3651 16745 3660 16779
rect 3608 16736 3660 16745
rect 4528 16779 4580 16788
rect 4528 16745 4537 16779
rect 4537 16745 4571 16779
rect 4571 16745 4580 16779
rect 4528 16736 4580 16745
rect 5724 16779 5776 16788
rect 5724 16745 5733 16779
rect 5733 16745 5767 16779
rect 5767 16745 5776 16779
rect 5724 16736 5776 16745
rect 6184 16779 6236 16788
rect 6184 16745 6193 16779
rect 6193 16745 6227 16779
rect 6227 16745 6236 16779
rect 6184 16736 6236 16745
rect 6644 16779 6696 16788
rect 6644 16745 6653 16779
rect 6653 16745 6687 16779
rect 6687 16745 6696 16779
rect 6644 16736 6696 16745
rect 10600 16736 10652 16788
rect 3792 16668 3844 16720
rect 4988 16668 5040 16720
rect 2688 16600 2740 16652
rect 2780 16600 2832 16652
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 3700 16532 3752 16584
rect 4804 16532 4856 16584
rect 5448 16600 5500 16652
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 7656 16668 7708 16720
rect 11336 16736 11388 16788
rect 11152 16668 11204 16720
rect 11796 16736 11848 16788
rect 12900 16736 12952 16788
rect 13544 16736 13596 16788
rect 16580 16736 16632 16788
rect 21088 16779 21140 16788
rect 21088 16745 21097 16779
rect 21097 16745 21131 16779
rect 21131 16745 21140 16779
rect 21088 16736 21140 16745
rect 14280 16668 14332 16720
rect 7472 16643 7524 16652
rect 7472 16609 7506 16643
rect 7506 16609 7524 16643
rect 7472 16600 7524 16609
rect 8208 16600 8260 16652
rect 3148 16464 3200 16516
rect 3424 16464 3476 16516
rect 4896 16464 4948 16516
rect 5632 16532 5684 16584
rect 5908 16575 5960 16584
rect 5908 16541 5917 16575
rect 5917 16541 5951 16575
rect 5951 16541 5960 16575
rect 5908 16532 5960 16541
rect 6644 16532 6696 16584
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 9220 16575 9272 16584
rect 9220 16541 9229 16575
rect 9229 16541 9263 16575
rect 9263 16541 9272 16575
rect 9220 16532 9272 16541
rect 5356 16439 5408 16448
rect 5356 16405 5365 16439
rect 5365 16405 5399 16439
rect 5399 16405 5408 16439
rect 5356 16396 5408 16405
rect 9404 16464 9456 16516
rect 9772 16600 9824 16652
rect 10692 16600 10744 16652
rect 11796 16600 11848 16652
rect 12532 16600 12584 16652
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 14648 16643 14700 16652
rect 14648 16609 14657 16643
rect 14657 16609 14691 16643
rect 14691 16609 14700 16643
rect 14648 16600 14700 16609
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 11520 16575 11572 16584
rect 9772 16464 9824 16516
rect 10416 16464 10468 16516
rect 8116 16396 8168 16448
rect 8668 16396 8720 16448
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 13268 16532 13320 16584
rect 14556 16532 14608 16584
rect 16120 16668 16172 16720
rect 15200 16600 15252 16652
rect 17224 16600 17276 16652
rect 19524 16600 19576 16652
rect 20812 16600 20864 16652
rect 20904 16643 20956 16652
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 20904 16600 20956 16609
rect 16672 16507 16724 16516
rect 16672 16473 16681 16507
rect 16681 16473 16715 16507
rect 16715 16473 16724 16507
rect 16672 16464 16724 16473
rect 10876 16396 10928 16448
rect 13636 16396 13688 16448
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 3700 16235 3752 16244
rect 3700 16201 3709 16235
rect 3709 16201 3743 16235
rect 3743 16201 3752 16235
rect 3700 16192 3752 16201
rect 4252 16192 4304 16244
rect 5172 16192 5224 16244
rect 6368 16192 6420 16244
rect 8208 16235 8260 16244
rect 1952 16167 2004 16176
rect 1952 16133 1961 16167
rect 1961 16133 1995 16167
rect 1995 16133 2004 16167
rect 1952 16124 2004 16133
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 10140 16192 10192 16244
rect 4896 16056 4948 16108
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 10140 16056 10192 16108
rect 10784 16056 10836 16108
rect 11980 16192 12032 16244
rect 13268 16192 13320 16244
rect 13820 16192 13872 16244
rect 14648 16192 14700 16244
rect 17960 16192 18012 16244
rect 20352 16235 20404 16244
rect 20352 16201 20361 16235
rect 20361 16201 20395 16235
rect 20395 16201 20404 16235
rect 20352 16192 20404 16201
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 13360 16124 13412 16176
rect 14096 16124 14148 16176
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 2228 15988 2280 16040
rect 3424 15988 3476 16040
rect 4068 15988 4120 16040
rect 7656 15988 7708 16040
rect 8668 15988 8720 16040
rect 12256 15988 12308 16040
rect 12624 16056 12676 16108
rect 14188 16056 14240 16108
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14004 15988 14056 16040
rect 2412 15920 2464 15972
rect 3884 15920 3936 15972
rect 5540 15963 5592 15972
rect 5540 15929 5574 15963
rect 5574 15929 5592 15963
rect 5540 15920 5592 15929
rect 2688 15852 2740 15904
rect 3516 15852 3568 15904
rect 4896 15895 4948 15904
rect 4896 15861 4905 15895
rect 4905 15861 4939 15895
rect 4939 15861 4948 15895
rect 6644 15895 6696 15904
rect 4896 15852 4948 15861
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 8576 15852 8628 15904
rect 11152 15963 11204 15972
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 11152 15929 11186 15963
rect 11186 15929 11204 15963
rect 11152 15920 11204 15929
rect 19524 16124 19576 16176
rect 16488 16056 16540 16108
rect 17132 16056 17184 16108
rect 14280 15963 14332 15972
rect 14280 15929 14289 15963
rect 14289 15929 14323 15963
rect 14323 15929 14332 15963
rect 19432 15988 19484 16040
rect 20628 16056 20680 16108
rect 20168 16031 20220 16040
rect 20168 15997 20177 16031
rect 20177 15997 20211 16031
rect 20211 15997 20220 16031
rect 20168 15988 20220 15997
rect 20904 16031 20956 16040
rect 14280 15920 14332 15929
rect 18604 15920 18656 15972
rect 19340 15920 19392 15972
rect 20904 15997 20913 16031
rect 20913 15997 20947 16031
rect 20947 15997 20956 16031
rect 20904 15988 20956 15997
rect 10416 15852 10468 15861
rect 11060 15852 11112 15904
rect 12532 15852 12584 15904
rect 13360 15852 13412 15904
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 15108 15895 15160 15904
rect 14372 15852 14424 15861
rect 15108 15861 15117 15895
rect 15117 15861 15151 15895
rect 15151 15861 15160 15895
rect 15108 15852 15160 15861
rect 16396 15895 16448 15904
rect 16396 15861 16405 15895
rect 16405 15861 16439 15895
rect 16439 15861 16448 15895
rect 16396 15852 16448 15861
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 17960 15852 18012 15904
rect 20628 15852 20680 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 2780 15648 2832 15700
rect 3056 15648 3108 15700
rect 5172 15648 5224 15700
rect 6552 15648 6604 15700
rect 8852 15648 8904 15700
rect 9956 15648 10008 15700
rect 12072 15691 12124 15700
rect 12072 15657 12081 15691
rect 12081 15657 12115 15691
rect 12115 15657 12124 15691
rect 12072 15648 12124 15657
rect 12808 15648 12860 15700
rect 13360 15691 13412 15700
rect 13360 15657 13369 15691
rect 13369 15657 13403 15691
rect 13403 15657 13412 15691
rect 13360 15648 13412 15657
rect 13636 15648 13688 15700
rect 14372 15648 14424 15700
rect 15108 15648 15160 15700
rect 16396 15648 16448 15700
rect 18512 15648 18564 15700
rect 20260 15691 20312 15700
rect 20260 15657 20269 15691
rect 20269 15657 20303 15691
rect 20303 15657 20312 15691
rect 20260 15648 20312 15657
rect 1768 15623 1820 15632
rect 1768 15589 1777 15623
rect 1777 15589 1811 15623
rect 1811 15589 1820 15623
rect 1768 15580 1820 15589
rect 8024 15580 8076 15632
rect 11980 15580 12032 15632
rect 2136 15512 2188 15564
rect 1308 15444 1360 15496
rect 6552 15512 6604 15564
rect 7196 15555 7248 15564
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 9128 15512 9180 15564
rect 9956 15512 10008 15564
rect 10140 15555 10192 15564
rect 10140 15521 10174 15555
rect 10174 15521 10192 15555
rect 10140 15512 10192 15521
rect 12164 15512 12216 15564
rect 12440 15512 12492 15564
rect 2412 15444 2464 15496
rect 3424 15487 3476 15496
rect 3424 15453 3433 15487
rect 3433 15453 3467 15487
rect 3467 15453 3476 15487
rect 3424 15444 3476 15453
rect 3884 15444 3936 15496
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 8392 15444 8444 15496
rect 6920 15376 6972 15428
rect 5540 15308 5592 15360
rect 7472 15308 7524 15360
rect 9588 15444 9640 15496
rect 12072 15444 12124 15496
rect 12900 15580 12952 15632
rect 14004 15580 14056 15632
rect 19156 15580 19208 15632
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 16488 15555 16540 15564
rect 16488 15521 16522 15555
rect 16522 15521 16540 15555
rect 16488 15512 16540 15521
rect 18972 15512 19024 15564
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 10876 15376 10928 15428
rect 13636 15444 13688 15496
rect 13728 15376 13780 15428
rect 14464 15444 14516 15496
rect 15200 15444 15252 15496
rect 18788 15487 18840 15496
rect 17592 15419 17644 15428
rect 17592 15385 17601 15419
rect 17601 15385 17635 15419
rect 17635 15385 17644 15419
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 19892 15444 19944 15496
rect 17592 15376 17644 15385
rect 11152 15308 11204 15360
rect 19248 15308 19300 15360
rect 20444 15308 20496 15360
rect 21088 15351 21140 15360
rect 21088 15317 21097 15351
rect 21097 15317 21131 15351
rect 21131 15317 21140 15351
rect 21088 15308 21140 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 2780 15104 2832 15156
rect 2872 15104 2924 15156
rect 7196 15147 7248 15156
rect 7196 15113 7205 15147
rect 7205 15113 7239 15147
rect 7239 15113 7248 15147
rect 7196 15104 7248 15113
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 9956 15104 10008 15156
rect 2044 14900 2096 14952
rect 3792 15036 3844 15088
rect 6184 15036 6236 15088
rect 7472 15036 7524 15088
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 4804 15011 4856 15020
rect 4804 14977 4813 15011
rect 4813 14977 4847 15011
rect 4847 14977 4856 15011
rect 4804 14968 4856 14977
rect 5908 15011 5960 15020
rect 5908 14977 5917 15011
rect 5917 14977 5951 15011
rect 5951 14977 5960 15011
rect 5908 14968 5960 14977
rect 6644 14968 6696 15020
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 8852 15011 8904 15020
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 10140 14968 10192 15020
rect 10692 15036 10744 15088
rect 15016 15036 15068 15088
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 4896 14832 4948 14884
rect 7288 14900 7340 14952
rect 7932 14900 7984 14952
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 10876 14900 10928 14952
rect 11428 14968 11480 15020
rect 13912 14968 13964 15020
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 13636 14900 13688 14952
rect 9312 14832 9364 14884
rect 14280 14832 14332 14884
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 2320 14807 2372 14816
rect 2320 14773 2329 14807
rect 2329 14773 2363 14807
rect 2363 14773 2372 14807
rect 2320 14764 2372 14773
rect 2964 14764 3016 14816
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 5724 14807 5776 14816
rect 5724 14773 5733 14807
rect 5733 14773 5767 14807
rect 5767 14773 5776 14807
rect 5724 14764 5776 14773
rect 6000 14764 6052 14816
rect 6276 14764 6328 14816
rect 8484 14764 8536 14816
rect 10784 14764 10836 14816
rect 10968 14764 11020 14816
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 11888 14807 11940 14816
rect 11152 14764 11204 14773
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 11980 14807 12032 14816
rect 11980 14773 11989 14807
rect 11989 14773 12023 14807
rect 12023 14773 12032 14807
rect 13176 14807 13228 14816
rect 11980 14764 12032 14773
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 13728 14764 13780 14816
rect 13820 14764 13872 14816
rect 14556 14764 14608 14816
rect 16856 15104 16908 15156
rect 18604 15104 18656 15156
rect 19708 15104 19760 15156
rect 16672 15036 16724 15088
rect 15200 14968 15252 15020
rect 16396 14900 16448 14952
rect 17500 14943 17552 14952
rect 17500 14909 17509 14943
rect 17509 14909 17543 14943
rect 17543 14909 17552 14943
rect 17500 14900 17552 14909
rect 17960 14900 18012 14952
rect 18880 15036 18932 15088
rect 18788 14968 18840 15020
rect 20536 15036 20588 15088
rect 20720 14900 20772 14952
rect 20260 14832 20312 14884
rect 15936 14764 15988 14816
rect 16028 14764 16080 14816
rect 16488 14764 16540 14816
rect 18420 14764 18472 14816
rect 18696 14764 18748 14816
rect 19708 14764 19760 14816
rect 20352 14807 20404 14816
rect 20352 14773 20361 14807
rect 20361 14773 20395 14807
rect 20395 14773 20404 14807
rect 20352 14764 20404 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 3792 14560 3844 14612
rect 4068 14560 4120 14612
rect 6000 14603 6052 14612
rect 2872 14492 2924 14544
rect 3056 14424 3108 14476
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 3240 14356 3292 14408
rect 3608 14399 3660 14408
rect 3608 14365 3617 14399
rect 3617 14365 3651 14399
rect 3651 14365 3660 14399
rect 3608 14356 3660 14365
rect 4804 14492 4856 14544
rect 6000 14569 6009 14603
rect 6009 14569 6043 14603
rect 6043 14569 6052 14603
rect 6000 14560 6052 14569
rect 6460 14560 6512 14612
rect 7196 14560 7248 14612
rect 7656 14603 7708 14612
rect 7656 14569 7665 14603
rect 7665 14569 7699 14603
rect 7699 14569 7708 14603
rect 7656 14560 7708 14569
rect 6736 14492 6788 14544
rect 7104 14424 7156 14476
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 6092 14356 6144 14408
rect 6276 14356 6328 14408
rect 6552 14399 6604 14408
rect 6552 14365 6561 14399
rect 6561 14365 6595 14399
rect 6595 14365 6604 14399
rect 7288 14399 7340 14408
rect 6552 14356 6604 14365
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 7472 14399 7524 14408
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 7472 14356 7524 14365
rect 7656 14424 7708 14476
rect 8852 14560 8904 14612
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 11060 14560 11112 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 14004 14560 14056 14612
rect 14188 14560 14240 14612
rect 15936 14560 15988 14612
rect 16488 14560 16540 14612
rect 8116 14492 8168 14544
rect 13636 14492 13688 14544
rect 17592 14492 17644 14544
rect 17684 14492 17736 14544
rect 19340 14492 19392 14544
rect 19892 14535 19944 14544
rect 19892 14501 19901 14535
rect 19901 14501 19935 14535
rect 19935 14501 19944 14535
rect 19892 14492 19944 14501
rect 20076 14492 20128 14544
rect 8208 14467 8260 14476
rect 8208 14433 8242 14467
rect 8242 14433 8260 14467
rect 8208 14424 8260 14433
rect 9404 14356 9456 14408
rect 7932 14288 7984 14340
rect 9312 14331 9364 14340
rect 9312 14297 9321 14331
rect 9321 14297 9355 14331
rect 9355 14297 9364 14331
rect 9312 14288 9364 14297
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 2780 14220 2832 14272
rect 3056 14220 3108 14272
rect 3332 14220 3384 14272
rect 5172 14220 5224 14272
rect 7748 14220 7800 14272
rect 8852 14220 8904 14272
rect 9036 14220 9088 14272
rect 9404 14220 9456 14272
rect 10048 14220 10100 14272
rect 11060 14356 11112 14408
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11612 14424 11664 14476
rect 12256 14424 12308 14476
rect 11336 14356 11388 14365
rect 11704 14356 11756 14408
rect 11980 14288 12032 14340
rect 10968 14220 11020 14272
rect 13820 14424 13872 14476
rect 14004 14424 14056 14476
rect 15568 14424 15620 14476
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 16028 14356 16080 14408
rect 16212 14399 16264 14408
rect 16212 14365 16221 14399
rect 16221 14365 16255 14399
rect 16255 14365 16264 14399
rect 16212 14356 16264 14365
rect 18512 14424 18564 14476
rect 19248 14424 19300 14476
rect 16580 14356 16632 14408
rect 16948 14356 17000 14408
rect 19892 14356 19944 14408
rect 17868 14220 17920 14272
rect 21180 14220 21232 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 4804 14016 4856 14068
rect 5448 14016 5500 14068
rect 5908 14059 5960 14068
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 6092 14016 6144 14068
rect 1860 13812 1912 13864
rect 2044 13812 2096 13864
rect 1676 13676 1728 13728
rect 3884 13812 3936 13864
rect 4068 13812 4120 13864
rect 3700 13744 3752 13796
rect 3884 13676 3936 13728
rect 5816 13812 5868 13864
rect 5540 13744 5592 13796
rect 6368 13948 6420 14000
rect 10416 14016 10468 14068
rect 11060 14016 11112 14068
rect 13176 14016 13228 14068
rect 16396 14016 16448 14068
rect 16580 14016 16632 14068
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10416 13880 10468 13932
rect 11888 13948 11940 14000
rect 13912 13948 13964 14000
rect 18512 13948 18564 14000
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 11612 13880 11664 13932
rect 6736 13812 6788 13864
rect 7104 13855 7156 13864
rect 7104 13821 7138 13855
rect 7138 13821 7156 13855
rect 7104 13812 7156 13821
rect 10232 13812 10284 13864
rect 10692 13812 10744 13864
rect 10876 13812 10928 13864
rect 11704 13812 11756 13864
rect 12072 13812 12124 13864
rect 12256 13812 12308 13864
rect 13820 13812 13872 13864
rect 15200 13880 15252 13932
rect 7656 13744 7708 13796
rect 6276 13676 6328 13728
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 10048 13744 10100 13796
rect 11152 13744 11204 13796
rect 12164 13744 12216 13796
rect 13084 13744 13136 13796
rect 13728 13744 13780 13796
rect 15660 13855 15712 13864
rect 15660 13821 15694 13855
rect 15694 13821 15712 13855
rect 15660 13812 15712 13821
rect 16028 13812 16080 13864
rect 17868 13880 17920 13932
rect 18420 13880 18472 13932
rect 19064 13880 19116 13932
rect 19892 14016 19944 14068
rect 20444 13880 20496 13932
rect 20720 13923 20772 13932
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 20720 13880 20772 13889
rect 18328 13812 18380 13864
rect 16948 13744 17000 13796
rect 17408 13787 17460 13796
rect 17408 13753 17417 13787
rect 17417 13753 17451 13787
rect 17451 13753 17460 13787
rect 17408 13744 17460 13753
rect 18696 13744 18748 13796
rect 10416 13676 10468 13728
rect 10692 13719 10744 13728
rect 10692 13685 10701 13719
rect 10701 13685 10735 13719
rect 10735 13685 10744 13719
rect 10692 13676 10744 13685
rect 10784 13719 10836 13728
rect 10784 13685 10793 13719
rect 10793 13685 10827 13719
rect 10827 13685 10836 13719
rect 10784 13676 10836 13685
rect 11704 13676 11756 13728
rect 13452 13676 13504 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 15016 13676 15068 13728
rect 17316 13676 17368 13728
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 18512 13719 18564 13728
rect 18512 13685 18521 13719
rect 18521 13685 18555 13719
rect 18555 13685 18564 13719
rect 18512 13676 18564 13685
rect 19984 13744 20036 13796
rect 20628 13812 20680 13864
rect 19340 13719 19392 13728
rect 19340 13685 19349 13719
rect 19349 13685 19383 13719
rect 19383 13685 19392 13719
rect 19340 13676 19392 13685
rect 19524 13676 19576 13728
rect 20352 13676 20404 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2872 13472 2924 13524
rect 3516 13472 3568 13524
rect 3608 13472 3660 13524
rect 4896 13515 4948 13524
rect 4896 13481 4905 13515
rect 4905 13481 4939 13515
rect 4939 13481 4948 13515
rect 4896 13472 4948 13481
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 5816 13472 5868 13524
rect 8760 13472 8812 13524
rect 1860 13447 1912 13456
rect 1860 13413 1869 13447
rect 1869 13413 1903 13447
rect 1903 13413 1912 13447
rect 1860 13404 1912 13413
rect 1952 13336 2004 13388
rect 2964 13336 3016 13388
rect 4712 13336 4764 13388
rect 6092 13379 6144 13388
rect 1860 13268 1912 13320
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 2780 13268 2832 13277
rect 5356 13311 5408 13320
rect 2504 13200 2556 13252
rect 3700 13200 3752 13252
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 6092 13345 6101 13379
rect 6101 13345 6135 13379
rect 6135 13345 6144 13379
rect 6092 13336 6144 13345
rect 5448 13268 5500 13277
rect 6276 13268 6328 13320
rect 6552 13268 6604 13320
rect 6092 13200 6144 13252
rect 6828 13336 6880 13388
rect 8208 13379 8260 13388
rect 8208 13345 8217 13379
rect 8217 13345 8251 13379
rect 8251 13345 8260 13379
rect 8208 13336 8260 13345
rect 8392 13404 8444 13456
rect 13268 13472 13320 13524
rect 13452 13515 13504 13524
rect 13452 13481 13461 13515
rect 13461 13481 13495 13515
rect 13495 13481 13504 13515
rect 13452 13472 13504 13481
rect 14096 13472 14148 13524
rect 14280 13515 14332 13524
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 16212 13472 16264 13524
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 18420 13472 18472 13524
rect 19064 13515 19116 13524
rect 19064 13481 19073 13515
rect 19073 13481 19107 13515
rect 19107 13481 19116 13515
rect 19064 13472 19116 13481
rect 20076 13472 20128 13524
rect 20904 13472 20956 13524
rect 10876 13404 10928 13456
rect 12808 13404 12860 13456
rect 17592 13404 17644 13456
rect 11060 13379 11112 13388
rect 6920 13200 6972 13252
rect 7748 13268 7800 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 8300 13200 8352 13252
rect 11060 13345 11069 13379
rect 11069 13345 11103 13379
rect 11103 13345 11112 13379
rect 11060 13336 11112 13345
rect 10416 13268 10468 13320
rect 11612 13268 11664 13320
rect 13360 13336 13412 13388
rect 13452 13336 13504 13388
rect 13820 13336 13872 13388
rect 14648 13379 14700 13388
rect 14648 13345 14657 13379
rect 14657 13345 14691 13379
rect 14691 13345 14700 13379
rect 14648 13336 14700 13345
rect 15660 13379 15712 13388
rect 13084 13268 13136 13320
rect 13268 13268 13320 13320
rect 13636 13268 13688 13320
rect 13728 13268 13780 13320
rect 14372 13268 14424 13320
rect 15016 13268 15068 13320
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 15844 13336 15896 13388
rect 16948 13336 17000 13388
rect 17960 13379 18012 13388
rect 17960 13345 17994 13379
rect 17994 13345 18012 13379
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 17960 13336 18012 13345
rect 19248 13336 19300 13388
rect 20904 13379 20956 13388
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 10600 13200 10652 13252
rect 3332 13132 3384 13184
rect 5080 13132 5132 13184
rect 5448 13132 5500 13184
rect 8760 13132 8812 13184
rect 10324 13132 10376 13184
rect 12440 13132 12492 13184
rect 15568 13200 15620 13252
rect 16396 13200 16448 13252
rect 12808 13132 12860 13184
rect 14004 13132 14056 13184
rect 17040 13132 17092 13184
rect 18788 13132 18840 13184
rect 20444 13132 20496 13184
rect 20628 13132 20680 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1768 12971 1820 12980
rect 1768 12937 1777 12971
rect 1777 12937 1811 12971
rect 1811 12937 1820 12971
rect 1768 12928 1820 12937
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 2596 12928 2648 12980
rect 2320 12792 2372 12844
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 3884 12928 3936 12980
rect 5356 12928 5408 12980
rect 5540 12928 5592 12980
rect 6828 12971 6880 12980
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 7656 12971 7708 12980
rect 7656 12937 7665 12971
rect 7665 12937 7699 12971
rect 7699 12937 7708 12971
rect 7656 12928 7708 12937
rect 8208 12928 8260 12980
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 11060 12928 11112 12980
rect 12440 12928 12492 12980
rect 6736 12860 6788 12912
rect 6920 12860 6972 12912
rect 7196 12860 7248 12912
rect 6552 12792 6604 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 11520 12860 11572 12912
rect 12256 12860 12308 12912
rect 14740 12928 14792 12980
rect 15292 12928 15344 12980
rect 15752 12928 15804 12980
rect 16120 12928 16172 12980
rect 18512 12928 18564 12980
rect 18696 12928 18748 12980
rect 19340 12928 19392 12980
rect 19984 12928 20036 12980
rect 14372 12860 14424 12912
rect 15108 12860 15160 12912
rect 15936 12860 15988 12912
rect 19892 12860 19944 12912
rect 9220 12792 9272 12844
rect 10784 12792 10836 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 15568 12792 15620 12844
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 16672 12792 16724 12844
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17960 12792 18012 12844
rect 18696 12792 18748 12844
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 7564 12724 7616 12776
rect 8116 12724 8168 12776
rect 9864 12724 9916 12776
rect 10600 12724 10652 12776
rect 15936 12724 15988 12776
rect 17684 12724 17736 12776
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 20352 12724 20404 12776
rect 2044 12656 2096 12708
rect 3516 12699 3568 12708
rect 3516 12665 3550 12699
rect 3550 12665 3568 12699
rect 3516 12656 3568 12665
rect 5724 12656 5776 12708
rect 7104 12656 7156 12708
rect 10232 12656 10284 12708
rect 10968 12656 11020 12708
rect 1768 12588 1820 12640
rect 8208 12588 8260 12640
rect 8484 12588 8536 12640
rect 11060 12588 11112 12640
rect 11152 12588 11204 12640
rect 12624 12588 12676 12640
rect 15108 12631 15160 12640
rect 15108 12597 15117 12631
rect 15117 12597 15151 12631
rect 15151 12597 15160 12631
rect 15108 12588 15160 12597
rect 16672 12656 16724 12708
rect 16856 12699 16908 12708
rect 16856 12665 16865 12699
rect 16865 12665 16899 12699
rect 16899 12665 16908 12699
rect 16856 12656 16908 12665
rect 17776 12656 17828 12708
rect 18788 12656 18840 12708
rect 19156 12656 19208 12708
rect 19432 12656 19484 12708
rect 16120 12588 16172 12640
rect 17316 12588 17368 12640
rect 17960 12588 18012 12640
rect 18604 12588 18656 12640
rect 18880 12588 18932 12640
rect 19340 12588 19392 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2780 12384 2832 12436
rect 3516 12384 3568 12436
rect 5540 12384 5592 12436
rect 7380 12384 7432 12436
rect 4804 12316 4856 12368
rect 4988 12316 5040 12368
rect 6736 12316 6788 12368
rect 6920 12316 6972 12368
rect 11612 12384 11664 12436
rect 11704 12384 11756 12436
rect 13360 12384 13412 12436
rect 14004 12384 14056 12436
rect 15108 12384 15160 12436
rect 16212 12384 16264 12436
rect 16396 12384 16448 12436
rect 16580 12384 16632 12436
rect 2136 12291 2188 12300
rect 2136 12257 2170 12291
rect 2170 12257 2188 12291
rect 2136 12248 2188 12257
rect 3332 12291 3384 12300
rect 3332 12257 3341 12291
rect 3341 12257 3375 12291
rect 3375 12257 3384 12291
rect 3332 12248 3384 12257
rect 6184 12248 6236 12300
rect 7380 12248 7432 12300
rect 8484 12248 8536 12300
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 1676 12087 1728 12096
rect 1676 12053 1685 12087
rect 1685 12053 1719 12087
rect 1719 12053 1728 12087
rect 1676 12044 1728 12053
rect 3976 12112 4028 12164
rect 2136 12044 2188 12096
rect 2596 12044 2648 12096
rect 4712 12044 4764 12096
rect 8208 12180 8260 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 7472 12155 7524 12164
rect 7472 12121 7481 12155
rect 7481 12121 7515 12155
rect 7515 12121 7524 12155
rect 7472 12112 7524 12121
rect 7840 12112 7892 12164
rect 6276 12044 6328 12096
rect 6828 12044 6880 12096
rect 8668 12044 8720 12096
rect 10784 12248 10836 12300
rect 12164 12316 12216 12368
rect 17868 12359 17920 12368
rect 17868 12325 17902 12359
rect 17902 12325 17920 12359
rect 17868 12316 17920 12325
rect 18696 12384 18748 12436
rect 19432 12384 19484 12436
rect 19800 12384 19852 12436
rect 20444 12316 20496 12368
rect 11704 12248 11756 12300
rect 13912 12291 13964 12300
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 13912 12248 13964 12257
rect 14372 12248 14424 12300
rect 9864 12180 9916 12232
rect 11520 12180 11572 12232
rect 15384 12248 15436 12300
rect 15568 12291 15620 12300
rect 15568 12257 15602 12291
rect 15602 12257 15620 12291
rect 15568 12248 15620 12257
rect 16396 12248 16448 12300
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 19248 12248 19300 12300
rect 20996 12291 21048 12300
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 10048 12044 10100 12096
rect 10508 12044 10560 12096
rect 10876 12044 10928 12096
rect 11152 12044 11204 12096
rect 15108 12180 15160 12232
rect 16304 12180 16356 12232
rect 16764 12180 16816 12232
rect 15200 12112 15252 12164
rect 16948 12112 17000 12164
rect 12348 12044 12400 12096
rect 12992 12087 13044 12096
rect 12992 12053 13001 12087
rect 13001 12053 13035 12087
rect 13035 12053 13044 12087
rect 12992 12044 13044 12053
rect 14096 12044 14148 12096
rect 14556 12044 14608 12096
rect 17316 12044 17368 12096
rect 18604 12044 18656 12096
rect 20536 12044 20588 12096
rect 21180 12087 21232 12096
rect 21180 12053 21189 12087
rect 21189 12053 21223 12087
rect 21223 12053 21232 12087
rect 21180 12044 21232 12053
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 2136 11840 2188 11892
rect 4160 11840 4212 11892
rect 5080 11840 5132 11892
rect 7104 11840 7156 11892
rect 7748 11840 7800 11892
rect 8300 11883 8352 11892
rect 8300 11849 8309 11883
rect 8309 11849 8343 11883
rect 8343 11849 8352 11883
rect 8300 11840 8352 11849
rect 8484 11840 8536 11892
rect 8944 11840 8996 11892
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 6184 11772 6236 11824
rect 3884 11704 3936 11756
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 3976 11636 4028 11688
rect 2136 11568 2188 11620
rect 3792 11568 3844 11620
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 7840 11704 7892 11756
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 11796 11840 11848 11892
rect 15384 11840 15436 11892
rect 16028 11840 16080 11892
rect 16396 11840 16448 11892
rect 17960 11840 18012 11892
rect 9772 11772 9824 11824
rect 10048 11772 10100 11824
rect 10784 11747 10836 11756
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 16764 11772 16816 11824
rect 19708 11840 19760 11892
rect 18420 11772 18472 11824
rect 19156 11772 19208 11824
rect 2320 11500 2372 11552
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 4068 11543 4120 11552
rect 4068 11509 4077 11543
rect 4077 11509 4111 11543
rect 4111 11509 4120 11543
rect 4068 11500 4120 11509
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 4344 11500 4396 11552
rect 4620 11500 4672 11552
rect 6460 11568 6512 11620
rect 6736 11568 6788 11620
rect 10692 11636 10744 11688
rect 9036 11568 9088 11620
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 17868 11704 17920 11756
rect 18696 11704 18748 11756
rect 19708 11704 19760 11756
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 20904 11704 20956 11756
rect 12348 11636 12400 11688
rect 12992 11636 13044 11688
rect 13268 11636 13320 11688
rect 15108 11636 15160 11688
rect 16028 11679 16080 11688
rect 16028 11645 16062 11679
rect 16062 11645 16080 11679
rect 16028 11636 16080 11645
rect 18972 11636 19024 11688
rect 15292 11568 15344 11620
rect 18420 11611 18472 11620
rect 18420 11577 18429 11611
rect 18429 11577 18463 11611
rect 18463 11577 18472 11611
rect 18420 11568 18472 11577
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 8944 11500 8996 11552
rect 9220 11500 9272 11552
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 12900 11500 12952 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 17408 11500 17460 11552
rect 17592 11500 17644 11552
rect 18512 11543 18564 11552
rect 18512 11509 18521 11543
rect 18521 11509 18555 11543
rect 18555 11509 18564 11543
rect 18512 11500 18564 11509
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 19248 11500 19300 11509
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 1860 11296 1912 11348
rect 3700 11296 3752 11348
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 4160 11296 4212 11348
rect 5632 11296 5684 11348
rect 3240 11228 3292 11280
rect 3608 11228 3660 11280
rect 2596 11160 2648 11212
rect 3148 11160 3200 11212
rect 3976 11160 4028 11212
rect 6828 11160 6880 11212
rect 11612 11296 11664 11348
rect 13360 11296 13412 11348
rect 14372 11339 14424 11348
rect 8852 11228 8904 11280
rect 9128 11228 9180 11280
rect 9496 11228 9548 11280
rect 7840 11203 7892 11212
rect 7840 11169 7874 11203
rect 7874 11169 7892 11203
rect 7840 11160 7892 11169
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 3976 11024 4028 11076
rect 6184 11092 6236 11144
rect 6920 11092 6972 11144
rect 8944 11092 8996 11144
rect 9772 11092 9824 11144
rect 7196 11024 7248 11076
rect 7472 11024 7524 11076
rect 9496 11024 9548 11076
rect 10140 11024 10192 11076
rect 11612 11160 11664 11212
rect 12716 11160 12768 11212
rect 13820 11228 13872 11280
rect 14372 11305 14381 11339
rect 14381 11305 14415 11339
rect 14415 11305 14424 11339
rect 14372 11296 14424 11305
rect 15200 11296 15252 11348
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 16304 11296 16356 11348
rect 17684 11296 17736 11348
rect 19248 11296 19300 11348
rect 21088 11339 21140 11348
rect 21088 11305 21097 11339
rect 21097 11305 21131 11339
rect 21131 11305 21140 11339
rect 21088 11296 21140 11305
rect 17040 11228 17092 11280
rect 19432 11228 19484 11280
rect 19892 11228 19944 11280
rect 20352 11228 20404 11280
rect 14556 11160 14608 11212
rect 12440 11092 12492 11144
rect 14372 11092 14424 11144
rect 15292 11160 15344 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 15016 11092 15068 11144
rect 4988 10956 5040 11008
rect 5448 10956 5500 11008
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 9128 10956 9180 11008
rect 11980 10956 12032 11008
rect 13636 10956 13688 11008
rect 15292 11024 15344 11076
rect 16396 11092 16448 11144
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 17316 11092 17368 11144
rect 19340 11203 19392 11212
rect 19340 11169 19349 11203
rect 19349 11169 19383 11203
rect 19383 11169 19392 11203
rect 19340 11160 19392 11169
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 17868 11024 17920 11076
rect 18512 11092 18564 11144
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 19156 11092 19208 11144
rect 19616 10956 19668 11008
rect 20720 10999 20772 11008
rect 20720 10965 20729 10999
rect 20729 10965 20763 10999
rect 20763 10965 20772 10999
rect 20720 10956 20772 10965
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1768 10752 1820 10804
rect 3240 10795 3292 10804
rect 3240 10761 3249 10795
rect 3249 10761 3283 10795
rect 3283 10761 3292 10795
rect 3240 10752 3292 10761
rect 3792 10752 3844 10804
rect 3976 10684 4028 10736
rect 5264 10752 5316 10804
rect 7196 10752 7248 10804
rect 7380 10752 7432 10804
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 3148 10616 3200 10668
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 9128 10684 9180 10736
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 6000 10616 6052 10668
rect 8944 10616 8996 10668
rect 10784 10752 10836 10804
rect 11152 10752 11204 10804
rect 13360 10752 13412 10804
rect 15016 10752 15068 10804
rect 15660 10752 15712 10804
rect 16672 10752 16724 10804
rect 19892 10795 19944 10804
rect 12716 10684 12768 10736
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 4252 10548 4304 10600
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 2228 10412 2280 10464
rect 3240 10480 3292 10532
rect 4712 10480 4764 10532
rect 4988 10480 5040 10532
rect 6644 10480 6696 10532
rect 10876 10548 10928 10600
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 13268 10616 13320 10668
rect 13636 10616 13688 10668
rect 11152 10548 11204 10600
rect 12440 10548 12492 10600
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 13084 10548 13136 10600
rect 14280 10548 14332 10600
rect 15568 10616 15620 10668
rect 17316 10684 17368 10736
rect 18236 10684 18288 10736
rect 19892 10761 19901 10795
rect 19901 10761 19935 10795
rect 19935 10761 19944 10795
rect 19892 10752 19944 10761
rect 20720 10684 20772 10736
rect 20812 10684 20864 10736
rect 22560 10684 22612 10736
rect 16856 10548 16908 10600
rect 16948 10548 17000 10600
rect 11060 10480 11112 10532
rect 11796 10523 11848 10532
rect 11796 10489 11805 10523
rect 11805 10489 11839 10523
rect 11839 10489 11848 10523
rect 11796 10480 11848 10489
rect 11888 10480 11940 10532
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 2780 10412 2832 10421
rect 3792 10412 3844 10464
rect 5264 10412 5316 10464
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 5908 10412 5960 10464
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 7012 10455 7064 10464
rect 6184 10412 6236 10421
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 8208 10455 8260 10464
rect 7472 10412 7524 10421
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 8576 10455 8628 10464
rect 8576 10421 8585 10455
rect 8585 10421 8619 10455
rect 8619 10421 8628 10455
rect 8576 10412 8628 10421
rect 9036 10412 9088 10464
rect 11152 10412 11204 10464
rect 15108 10523 15160 10532
rect 15108 10489 15117 10523
rect 15117 10489 15151 10523
rect 15151 10489 15160 10523
rect 15108 10480 15160 10489
rect 16396 10480 16448 10532
rect 20996 10659 21048 10668
rect 17500 10480 17552 10532
rect 19892 10548 19944 10600
rect 20168 10548 20220 10600
rect 20352 10591 20404 10600
rect 20352 10557 20361 10591
rect 20361 10557 20395 10591
rect 20395 10557 20404 10591
rect 20352 10548 20404 10557
rect 18696 10480 18748 10532
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 20812 10591 20864 10600
rect 20812 10557 20821 10591
rect 20821 10557 20855 10591
rect 20855 10557 20864 10591
rect 20812 10548 20864 10557
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 13912 10412 13964 10464
rect 15016 10455 15068 10464
rect 15016 10421 15025 10455
rect 15025 10421 15059 10455
rect 15059 10421 15068 10455
rect 15016 10412 15068 10421
rect 15384 10412 15436 10464
rect 16764 10412 16816 10464
rect 19708 10412 19760 10464
rect 20444 10455 20496 10464
rect 20444 10421 20453 10455
rect 20453 10421 20487 10455
rect 20487 10421 20496 10455
rect 20444 10412 20496 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1952 10208 2004 10260
rect 2780 10208 2832 10260
rect 3516 10208 3568 10260
rect 3792 10208 3844 10260
rect 4068 10208 4120 10260
rect 6644 10208 6696 10260
rect 7472 10208 7524 10260
rect 3700 10140 3752 10192
rect 4344 10183 4396 10192
rect 4344 10149 4378 10183
rect 4378 10149 4396 10183
rect 4344 10140 4396 10149
rect 5448 10140 5500 10192
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 3148 10004 3200 10056
rect 3424 10072 3476 10124
rect 6276 10115 6328 10124
rect 3516 10004 3568 10056
rect 3884 10004 3936 10056
rect 6276 10081 6285 10115
rect 6285 10081 6319 10115
rect 6319 10081 6328 10115
rect 6276 10072 6328 10081
rect 6736 10140 6788 10192
rect 10692 10208 10744 10260
rect 11152 10208 11204 10260
rect 11980 10208 12032 10260
rect 13728 10208 13780 10260
rect 2412 9936 2464 9988
rect 2780 9936 2832 9988
rect 5908 9979 5960 9988
rect 5908 9945 5917 9979
rect 5917 9945 5951 9979
rect 5951 9945 5960 9979
rect 5908 9936 5960 9945
rect 3976 9868 4028 9920
rect 7472 10004 7524 10056
rect 8484 10140 8536 10192
rect 9220 10140 9272 10192
rect 10600 10140 10652 10192
rect 11704 10183 11756 10192
rect 11704 10149 11713 10183
rect 11713 10149 11747 10183
rect 11747 10149 11756 10183
rect 11704 10140 11756 10149
rect 14096 10208 14148 10260
rect 15752 10208 15804 10260
rect 16304 10208 16356 10260
rect 16396 10208 16448 10260
rect 18696 10208 18748 10260
rect 20352 10208 20404 10260
rect 16028 10140 16080 10192
rect 17960 10140 18012 10192
rect 19156 10140 19208 10192
rect 8944 10072 8996 10124
rect 10324 10072 10376 10124
rect 10968 10072 11020 10124
rect 11152 10072 11204 10124
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 12808 10072 12860 10124
rect 13728 10072 13780 10124
rect 14372 10072 14424 10124
rect 14740 10115 14792 10124
rect 14740 10081 14749 10115
rect 14749 10081 14783 10115
rect 14783 10081 14792 10115
rect 14740 10072 14792 10081
rect 15568 10115 15620 10124
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 9772 10004 9824 10056
rect 10784 10004 10836 10056
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 12624 10004 12676 10056
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13636 10004 13688 10056
rect 13820 10004 13872 10056
rect 14004 10004 14056 10056
rect 8484 9868 8536 9920
rect 11796 9868 11848 9920
rect 12532 9936 12584 9988
rect 14096 9936 14148 9988
rect 15568 10081 15602 10115
rect 15602 10081 15620 10115
rect 15568 10072 15620 10081
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 17500 10047 17552 10056
rect 15200 9936 15252 9988
rect 11980 9868 12032 9920
rect 15108 9868 15160 9920
rect 15660 9868 15712 9920
rect 17500 10013 17509 10047
rect 17509 10013 17543 10047
rect 17543 10013 17552 10047
rect 17500 10004 17552 10013
rect 20076 10047 20128 10056
rect 20076 10013 20085 10047
rect 20085 10013 20119 10047
rect 20119 10013 20128 10047
rect 20076 10004 20128 10013
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 1952 9664 2004 9716
rect 3148 9664 3200 9716
rect 4252 9664 4304 9716
rect 6000 9664 6052 9716
rect 8300 9664 8352 9716
rect 12808 9664 12860 9716
rect 8484 9596 8536 9648
rect 6276 9571 6328 9580
rect 6276 9537 6285 9571
rect 6285 9537 6319 9571
rect 6319 9537 6328 9571
rect 6276 9528 6328 9537
rect 2044 9460 2096 9512
rect 2504 9503 2556 9512
rect 2504 9469 2513 9503
rect 2513 9469 2547 9503
rect 2547 9469 2556 9503
rect 2504 9460 2556 9469
rect 3056 9392 3108 9444
rect 3884 9392 3936 9444
rect 4068 9392 4120 9444
rect 6000 9460 6052 9512
rect 7564 9460 7616 9512
rect 6736 9392 6788 9444
rect 10324 9596 10376 9648
rect 10968 9596 11020 9648
rect 15200 9664 15252 9716
rect 17500 9664 17552 9716
rect 8944 9528 8996 9580
rect 9864 9528 9916 9580
rect 11336 9571 11388 9580
rect 11336 9537 11345 9571
rect 11345 9537 11379 9571
rect 11379 9537 11388 9571
rect 11336 9528 11388 9537
rect 11428 9528 11480 9580
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 14004 9528 14056 9580
rect 14924 9528 14976 9580
rect 9496 9460 9548 9512
rect 8944 9435 8996 9444
rect 2688 9324 2740 9376
rect 2964 9324 3016 9376
rect 6000 9324 6052 9376
rect 6828 9324 6880 9376
rect 8944 9401 8953 9435
rect 8953 9401 8987 9435
rect 8987 9401 8996 9435
rect 8944 9392 8996 9401
rect 10508 9392 10560 9444
rect 8208 9324 8260 9376
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 9496 9324 9548 9333
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 10876 9324 10928 9376
rect 11888 9503 11940 9512
rect 11428 9392 11480 9444
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 17684 9596 17736 9648
rect 18880 9596 18932 9648
rect 19432 9639 19484 9648
rect 19432 9605 19441 9639
rect 19441 9605 19475 9639
rect 19475 9605 19484 9639
rect 19432 9596 19484 9605
rect 19984 9664 20036 9716
rect 15476 9528 15528 9580
rect 16764 9528 16816 9580
rect 19340 9528 19392 9580
rect 11980 9392 12032 9444
rect 13268 9392 13320 9444
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 14464 9392 14516 9444
rect 17316 9460 17368 9512
rect 18788 9460 18840 9512
rect 19800 9460 19852 9512
rect 21364 9596 21416 9648
rect 21548 9528 21600 9580
rect 16120 9392 16172 9444
rect 15200 9324 15252 9376
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 16580 9324 16632 9376
rect 19248 9392 19300 9444
rect 19984 9392 20036 9444
rect 16948 9324 17000 9376
rect 17224 9324 17276 9376
rect 19800 9367 19852 9376
rect 19800 9333 19809 9367
rect 19809 9333 19843 9367
rect 19843 9333 19852 9367
rect 19800 9324 19852 9333
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 20168 9324 20220 9376
rect 20536 9324 20588 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2228 9120 2280 9172
rect 3332 9120 3384 9172
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 6184 9120 6236 9172
rect 6828 9120 6880 9172
rect 7380 9120 7432 9172
rect 2964 9052 3016 9104
rect 3424 9052 3476 9104
rect 7012 9052 7064 9104
rect 7564 9052 7616 9104
rect 9588 9120 9640 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11704 9120 11756 9172
rect 8576 9095 8628 9104
rect 8576 9061 8585 9095
rect 8585 9061 8619 9095
rect 8619 9061 8628 9095
rect 8576 9052 8628 9061
rect 3148 8916 3200 8968
rect 3516 8984 3568 9036
rect 7104 8984 7156 9036
rect 8300 8984 8352 9036
rect 10968 9052 11020 9104
rect 12164 9052 12216 9104
rect 13820 9052 13872 9104
rect 14372 9095 14424 9104
rect 3608 8916 3660 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6736 8916 6788 8968
rect 8852 8916 8904 8968
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 10876 8984 10928 9036
rect 13452 8984 13504 9036
rect 11060 8916 11112 8968
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 12808 8916 12860 8968
rect 12900 8916 12952 8968
rect 14004 8916 14056 8968
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 15016 9120 15068 9172
rect 15200 9120 15252 9172
rect 15476 9120 15528 9172
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 17960 9120 18012 9172
rect 18604 9120 18656 9172
rect 18880 9120 18932 9172
rect 20076 9120 20128 9172
rect 16672 9052 16724 9104
rect 16764 9052 16816 9104
rect 15016 8984 15068 9036
rect 15200 8984 15252 9036
rect 14832 8916 14884 8968
rect 19432 9052 19484 9104
rect 20536 9052 20588 9104
rect 18512 8984 18564 9036
rect 19248 8984 19300 9036
rect 20628 8984 20680 9036
rect 4712 8848 4764 8900
rect 6644 8848 6696 8900
rect 7932 8848 7984 8900
rect 15476 8848 15528 8900
rect 15660 8848 15712 8900
rect 17776 8916 17828 8968
rect 19340 8916 19392 8968
rect 19984 8916 20036 8968
rect 3424 8780 3476 8832
rect 6828 8780 6880 8832
rect 7012 8780 7064 8832
rect 8116 8780 8168 8832
rect 8668 8780 8720 8832
rect 10876 8780 10928 8832
rect 12808 8780 12860 8832
rect 12992 8780 13044 8832
rect 13728 8780 13780 8832
rect 13820 8780 13872 8832
rect 14464 8780 14516 8832
rect 20260 8848 20312 8900
rect 18512 8780 18564 8832
rect 18604 8780 18656 8832
rect 19156 8823 19208 8832
rect 19156 8789 19165 8823
rect 19165 8789 19199 8823
rect 19199 8789 19208 8823
rect 19156 8780 19208 8789
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2872 8576 2924 8628
rect 7288 8576 7340 8628
rect 7932 8576 7984 8628
rect 10508 8576 10560 8628
rect 11060 8576 11112 8628
rect 11704 8576 11756 8628
rect 12440 8576 12492 8628
rect 14372 8576 14424 8628
rect 16856 8576 16908 8628
rect 17132 8576 17184 8628
rect 18604 8576 18656 8628
rect 20812 8576 20864 8628
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 6920 8508 6972 8560
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 5540 8440 5592 8492
rect 6828 8440 6880 8492
rect 3332 8372 3384 8424
rect 6644 8372 6696 8424
rect 3976 8304 4028 8356
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 2780 8236 2832 8245
rect 3148 8236 3200 8288
rect 3792 8236 3844 8288
rect 5080 8236 5132 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 7472 8304 7524 8356
rect 9864 8508 9916 8560
rect 8116 8440 8168 8492
rect 12164 8508 12216 8560
rect 7748 8372 7800 8424
rect 9680 8372 9732 8424
rect 8576 8304 8628 8356
rect 9588 8304 9640 8356
rect 11152 8440 11204 8492
rect 12992 8440 13044 8492
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 13452 8508 13504 8560
rect 14740 8508 14792 8560
rect 15844 8508 15896 8560
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 16396 8440 16448 8492
rect 13728 8372 13780 8424
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 14372 8372 14424 8424
rect 17684 8508 17736 8560
rect 17408 8440 17460 8492
rect 17960 8440 18012 8492
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 19708 8440 19760 8492
rect 19800 8440 19852 8492
rect 20168 8440 20220 8492
rect 17776 8372 17828 8424
rect 10508 8304 10560 8356
rect 14464 8304 14516 8356
rect 14556 8304 14608 8356
rect 17040 8304 17092 8356
rect 7564 8236 7616 8288
rect 8392 8236 8444 8288
rect 9680 8236 9732 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 12808 8236 12860 8288
rect 13820 8236 13872 8288
rect 14280 8236 14332 8288
rect 15016 8279 15068 8288
rect 15016 8245 15025 8279
rect 15025 8245 15059 8279
rect 15059 8245 15068 8279
rect 15016 8236 15068 8245
rect 15384 8236 15436 8288
rect 15752 8236 15804 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 18512 8372 18564 8424
rect 19340 8415 19392 8424
rect 19340 8381 19349 8415
rect 19349 8381 19383 8415
rect 19383 8381 19392 8415
rect 19340 8372 19392 8381
rect 20628 8372 20680 8424
rect 19892 8304 19944 8356
rect 20536 8304 20588 8356
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3056 8032 3108 8084
rect 3608 8032 3660 8084
rect 3792 8032 3844 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 5908 8032 5960 8084
rect 7564 8032 7616 8084
rect 8944 8032 8996 8084
rect 3424 7896 3476 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 3884 7964 3936 8016
rect 6828 7964 6880 8016
rect 4068 7896 4120 7948
rect 4252 7896 4304 7948
rect 6276 7896 6328 7948
rect 9496 7964 9548 8016
rect 9956 8032 10008 8084
rect 11612 8032 11664 8084
rect 9772 7964 9824 8016
rect 10508 7964 10560 8016
rect 14096 8032 14148 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 14464 8032 14516 8084
rect 15384 8032 15436 8084
rect 17408 8032 17460 8084
rect 19156 8032 19208 8084
rect 20260 8032 20312 8084
rect 12992 7964 13044 8016
rect 13084 7964 13136 8016
rect 13728 7964 13780 8016
rect 17684 7964 17736 8016
rect 18696 7964 18748 8016
rect 19432 8007 19484 8016
rect 19432 7973 19466 8007
rect 19466 7973 19484 8007
rect 19432 7964 19484 7973
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 8392 7896 8444 7948
rect 5908 7760 5960 7812
rect 6184 7760 6236 7812
rect 7840 7828 7892 7880
rect 7196 7760 7248 7812
rect 8760 7828 8812 7880
rect 3240 7692 3292 7744
rect 4068 7692 4120 7744
rect 8300 7692 8352 7744
rect 8944 7760 8996 7812
rect 10692 7896 10744 7948
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 12256 7896 12308 7948
rect 14004 7896 14056 7948
rect 9864 7828 9916 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 9772 7760 9824 7812
rect 12440 7828 12492 7880
rect 9588 7692 9640 7744
rect 11244 7760 11296 7812
rect 10692 7692 10744 7744
rect 11060 7692 11112 7744
rect 12348 7692 12400 7744
rect 13636 7828 13688 7880
rect 15108 7896 15160 7948
rect 16672 7896 16724 7948
rect 16856 7896 16908 7948
rect 18512 7896 18564 7948
rect 13636 7692 13688 7744
rect 15660 7692 15712 7744
rect 16396 7692 16448 7744
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 18972 7760 19024 7812
rect 16764 7692 16816 7744
rect 17684 7692 17736 7744
rect 20168 7692 20220 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 3608 7488 3660 7540
rect 4068 7488 4120 7540
rect 12348 7488 12400 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 14280 7488 14332 7540
rect 15476 7488 15528 7540
rect 1492 7352 1544 7404
rect 2780 7352 2832 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 2964 7148 3016 7200
rect 3240 7148 3292 7200
rect 3792 7420 3844 7472
rect 3884 7420 3936 7472
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 4436 7420 4488 7472
rect 6828 7420 6880 7472
rect 7196 7420 7248 7472
rect 7748 7420 7800 7472
rect 8116 7420 8168 7472
rect 8392 7463 8444 7472
rect 8392 7429 8401 7463
rect 8401 7429 8435 7463
rect 8435 7429 8444 7463
rect 8392 7420 8444 7429
rect 9956 7420 10008 7472
rect 10416 7420 10468 7472
rect 12072 7420 12124 7472
rect 18604 7488 18656 7540
rect 19892 7531 19944 7540
rect 19892 7497 19901 7531
rect 19901 7497 19935 7531
rect 19935 7497 19944 7531
rect 19892 7488 19944 7497
rect 17040 7463 17092 7472
rect 17040 7429 17049 7463
rect 17049 7429 17083 7463
rect 17083 7429 17092 7463
rect 17040 7420 17092 7429
rect 19432 7420 19484 7472
rect 3424 7352 3476 7361
rect 4344 7352 4396 7404
rect 3700 7284 3752 7336
rect 7840 7352 7892 7404
rect 4436 7216 4488 7268
rect 7196 7216 7248 7268
rect 3792 7148 3844 7200
rect 7564 7284 7616 7336
rect 9588 7352 9640 7404
rect 10232 7352 10284 7404
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 14556 7352 14608 7404
rect 17684 7395 17736 7404
rect 8208 7284 8260 7336
rect 10508 7327 10560 7336
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 10508 7284 10560 7293
rect 12440 7284 12492 7336
rect 13452 7284 13504 7336
rect 13820 7284 13872 7336
rect 13912 7284 13964 7336
rect 7932 7216 7984 7268
rect 7656 7148 7708 7200
rect 8944 7216 8996 7268
rect 8668 7148 8720 7200
rect 9496 7148 9548 7200
rect 9772 7148 9824 7200
rect 10600 7216 10652 7268
rect 11152 7259 11204 7268
rect 11152 7225 11186 7259
rect 11186 7225 11204 7259
rect 11152 7216 11204 7225
rect 11336 7216 11388 7268
rect 11520 7216 11572 7268
rect 12164 7148 12216 7200
rect 15016 7216 15068 7268
rect 15384 7216 15436 7268
rect 12348 7148 12400 7200
rect 12900 7148 12952 7200
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 14464 7148 14516 7200
rect 17684 7361 17693 7395
rect 17693 7361 17727 7395
rect 17727 7361 17736 7395
rect 17684 7352 17736 7361
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 16396 7284 16448 7336
rect 15936 7216 15988 7268
rect 18512 7284 18564 7336
rect 19708 7284 19760 7336
rect 15752 7148 15804 7200
rect 17224 7148 17276 7200
rect 18880 7216 18932 7268
rect 18144 7148 18196 7200
rect 18604 7148 18656 7200
rect 19248 7148 19300 7200
rect 19524 7148 19576 7200
rect 19800 7148 19852 7200
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 2320 6944 2372 6996
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 4896 6944 4948 6996
rect 7012 6944 7064 6996
rect 8484 6944 8536 6996
rect 8760 6987 8812 6996
rect 8760 6953 8769 6987
rect 8769 6953 8803 6987
rect 8803 6953 8812 6987
rect 8760 6944 8812 6953
rect 11060 6944 11112 6996
rect 11152 6944 11204 6996
rect 2044 6919 2096 6928
rect 2044 6885 2053 6919
rect 2053 6885 2087 6919
rect 2087 6885 2096 6919
rect 2044 6876 2096 6885
rect 1584 6808 1636 6860
rect 3608 6876 3660 6928
rect 4988 6876 5040 6928
rect 5172 6876 5224 6928
rect 7196 6876 7248 6928
rect 2780 6851 2832 6860
rect 2780 6817 2814 6851
rect 2814 6817 2832 6851
rect 2780 6808 2832 6817
rect 3976 6808 4028 6860
rect 4344 6808 4396 6860
rect 6000 6808 6052 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 6644 6715 6696 6724
rect 6644 6681 6653 6715
rect 6653 6681 6687 6715
rect 6687 6681 6696 6715
rect 6644 6672 6696 6681
rect 7656 6808 7708 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8024 6876 8076 6928
rect 8944 6876 8996 6928
rect 9312 6876 9364 6928
rect 10140 6919 10192 6928
rect 10140 6885 10149 6919
rect 10149 6885 10183 6919
rect 10183 6885 10192 6919
rect 10140 6876 10192 6885
rect 10508 6876 10560 6928
rect 10968 6876 11020 6928
rect 11520 6876 11572 6928
rect 12716 6944 12768 6996
rect 12992 6944 13044 6996
rect 15844 6944 15896 6996
rect 19156 6944 19208 6996
rect 19708 6987 19760 6996
rect 19708 6953 19717 6987
rect 19717 6953 19751 6987
rect 19751 6953 19760 6987
rect 19708 6944 19760 6953
rect 20260 6944 20312 6996
rect 7196 6783 7248 6792
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 7932 6783 7984 6792
rect 7012 6672 7064 6724
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 9772 6808 9824 6860
rect 9956 6808 10008 6860
rect 11060 6808 11112 6860
rect 13268 6851 13320 6860
rect 9588 6740 9640 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10968 6740 11020 6792
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 7472 6715 7524 6724
rect 7472 6681 7481 6715
rect 7481 6681 7515 6715
rect 7515 6681 7524 6715
rect 7472 6672 7524 6681
rect 7564 6672 7616 6724
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 13636 6876 13688 6928
rect 14096 6919 14148 6928
rect 14096 6885 14105 6919
rect 14105 6885 14139 6919
rect 14139 6885 14148 6919
rect 14096 6876 14148 6885
rect 14648 6876 14700 6928
rect 15108 6876 15160 6928
rect 16396 6876 16448 6928
rect 17960 6876 18012 6928
rect 18144 6876 18196 6928
rect 17868 6808 17920 6860
rect 18420 6808 18472 6860
rect 19432 6808 19484 6860
rect 19708 6808 19760 6860
rect 20168 6851 20220 6860
rect 20168 6817 20177 6851
rect 20177 6817 20211 6851
rect 20211 6817 20220 6851
rect 20168 6808 20220 6817
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 14924 6740 14976 6792
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16028 6740 16080 6792
rect 2872 6604 2924 6656
rect 6184 6647 6236 6656
rect 6184 6613 6193 6647
rect 6193 6613 6227 6647
rect 6227 6613 6236 6647
rect 6184 6604 6236 6613
rect 6736 6604 6788 6656
rect 8484 6604 8536 6656
rect 9956 6604 10008 6656
rect 10508 6647 10560 6656
rect 10508 6613 10517 6647
rect 10517 6613 10551 6647
rect 10551 6613 10560 6647
rect 10508 6604 10560 6613
rect 13820 6672 13872 6724
rect 15016 6672 15068 6724
rect 12440 6604 12492 6656
rect 12532 6604 12584 6656
rect 14556 6604 14608 6656
rect 17040 6647 17092 6656
rect 17040 6613 17049 6647
rect 17049 6613 17083 6647
rect 17083 6613 17092 6647
rect 17040 6604 17092 6613
rect 19524 6740 19576 6792
rect 19248 6604 19300 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 3976 6400 4028 6452
rect 6276 6400 6328 6452
rect 2780 6332 2832 6384
rect 4068 6332 4120 6384
rect 6736 6332 6788 6384
rect 2964 6264 3016 6316
rect 4252 6264 4304 6316
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 6184 6264 6236 6316
rect 7472 6400 7524 6452
rect 7748 6400 7800 6452
rect 1584 6196 1636 6248
rect 4160 6196 4212 6248
rect 4620 6196 4672 6248
rect 5816 6196 5868 6248
rect 12440 6400 12492 6452
rect 15384 6400 15436 6452
rect 17040 6400 17092 6452
rect 19156 6400 19208 6452
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 20444 6400 20496 6452
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 7748 6128 7800 6180
rect 7840 6128 7892 6180
rect 10508 6196 10560 6248
rect 8852 6128 8904 6180
rect 10232 6128 10284 6180
rect 10600 6128 10652 6180
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 5724 6060 5776 6112
rect 6552 6060 6604 6112
rect 8668 6060 8720 6112
rect 9588 6060 9640 6112
rect 10140 6060 10192 6112
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 13912 6332 13964 6384
rect 14004 6332 14056 6384
rect 12256 6264 12308 6316
rect 12716 6196 12768 6248
rect 15660 6264 15712 6316
rect 20168 6264 20220 6316
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 11704 6128 11756 6180
rect 12900 6171 12952 6180
rect 11980 6060 12032 6112
rect 12900 6137 12909 6171
rect 12909 6137 12943 6171
rect 12943 6137 12952 6171
rect 12900 6128 12952 6137
rect 17224 6196 17276 6248
rect 16672 6128 16724 6180
rect 17868 6128 17920 6180
rect 19616 6196 19668 6248
rect 20628 6196 20680 6248
rect 19248 6128 19300 6180
rect 20168 6128 20220 6180
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 14372 6060 14424 6112
rect 15016 6060 15068 6112
rect 15936 6060 15988 6112
rect 19616 6060 19668 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 2964 5899 3016 5908
rect 2964 5865 2973 5899
rect 2973 5865 3007 5899
rect 3007 5865 3016 5899
rect 2964 5856 3016 5865
rect 3516 5856 3568 5908
rect 4068 5856 4120 5908
rect 1768 5788 1820 5840
rect 5080 5788 5132 5840
rect 6184 5788 6236 5840
rect 6368 5856 6420 5908
rect 6920 5856 6972 5908
rect 7564 5856 7616 5908
rect 7748 5856 7800 5908
rect 8208 5856 8260 5908
rect 9496 5856 9548 5908
rect 10232 5856 10284 5908
rect 10692 5856 10744 5908
rect 11796 5856 11848 5908
rect 12072 5856 12124 5908
rect 14188 5856 14240 5908
rect 15384 5856 15436 5908
rect 17868 5856 17920 5908
rect 17960 5856 18012 5908
rect 18788 5856 18840 5908
rect 20076 5856 20128 5908
rect 6736 5788 6788 5840
rect 6828 5788 6880 5840
rect 10784 5788 10836 5840
rect 11704 5788 11756 5840
rect 12256 5788 12308 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 2688 5720 2740 5772
rect 4068 5720 4120 5772
rect 4712 5720 4764 5772
rect 5356 5720 5408 5772
rect 6552 5720 6604 5772
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7748 5763 7800 5772
rect 7196 5720 7248 5729
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9220 5720 9272 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 3700 5695 3752 5704
rect 3700 5661 3709 5695
rect 3709 5661 3743 5695
rect 3743 5661 3752 5695
rect 3700 5652 3752 5661
rect 5540 5652 5592 5704
rect 5816 5652 5868 5704
rect 6736 5695 6788 5704
rect 5172 5584 5224 5636
rect 6736 5661 6745 5695
rect 6745 5661 6779 5695
rect 6779 5661 6788 5695
rect 6736 5652 6788 5661
rect 8392 5652 8444 5704
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 5080 5516 5132 5568
rect 5264 5559 5316 5568
rect 5264 5525 5273 5559
rect 5273 5525 5307 5559
rect 5307 5525 5316 5559
rect 5264 5516 5316 5525
rect 6276 5516 6328 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 7564 5516 7616 5568
rect 9956 5652 10008 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 9496 5584 9548 5636
rect 13728 5720 13780 5772
rect 15200 5720 15252 5772
rect 10876 5652 10928 5704
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11244 5652 11296 5704
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 14188 5652 14240 5704
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 10508 5559 10560 5568
rect 10508 5525 10517 5559
rect 10517 5525 10551 5559
rect 10551 5525 10560 5559
rect 10508 5516 10560 5525
rect 10692 5516 10744 5568
rect 10876 5516 10928 5568
rect 11704 5516 11756 5568
rect 11980 5516 12032 5568
rect 15108 5584 15160 5636
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 15844 5720 15896 5772
rect 16028 5720 16080 5772
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 15660 5584 15712 5636
rect 16672 5584 16724 5636
rect 17960 5652 18012 5704
rect 19432 5788 19484 5840
rect 19616 5831 19668 5840
rect 19616 5797 19625 5831
rect 19625 5797 19659 5831
rect 19659 5797 19668 5831
rect 19616 5788 19668 5797
rect 19248 5652 19300 5704
rect 20260 5652 20312 5704
rect 20536 5788 20588 5840
rect 20720 5584 20772 5636
rect 20076 5516 20128 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 3516 5312 3568 5364
rect 4160 5312 4212 5364
rect 4988 5312 5040 5364
rect 8852 5355 8904 5364
rect 6368 5244 6420 5296
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 9128 5312 9180 5364
rect 9404 5312 9456 5364
rect 10232 5312 10284 5364
rect 12992 5312 13044 5364
rect 14004 5312 14056 5364
rect 14096 5312 14148 5364
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 18880 5355 18932 5364
rect 18880 5321 18889 5355
rect 18889 5321 18923 5355
rect 18923 5321 18932 5355
rect 18880 5312 18932 5321
rect 19340 5312 19392 5364
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 5080 5219 5132 5228
rect 5080 5185 5089 5219
rect 5089 5185 5123 5219
rect 5123 5185 5132 5219
rect 5080 5176 5132 5185
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 5632 5176 5684 5228
rect 6184 5176 6236 5228
rect 6736 5176 6788 5228
rect 6828 5176 6880 5228
rect 7288 5176 7340 5228
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 10048 5176 10100 5228
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 2504 5151 2556 5160
rect 2504 5117 2513 5151
rect 2513 5117 2547 5151
rect 2547 5117 2556 5151
rect 2504 5108 2556 5117
rect 3056 5108 3108 5160
rect 2872 5040 2924 5092
rect 3700 5108 3752 5160
rect 5264 5108 5316 5160
rect 9956 5151 10008 5160
rect 3608 5040 3660 5092
rect 4068 5040 4120 5092
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 10968 5108 11020 5160
rect 2228 4972 2280 5024
rect 2688 4972 2740 5024
rect 5172 4972 5224 5024
rect 6184 4972 6236 5024
rect 6552 4972 6604 5024
rect 7564 4972 7616 5024
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 10324 4972 10376 5024
rect 11060 5040 11112 5092
rect 12808 5244 12860 5296
rect 11888 5176 11940 5228
rect 13268 5176 13320 5228
rect 13912 5176 13964 5228
rect 16120 5244 16172 5296
rect 17408 5244 17460 5296
rect 19524 5244 19576 5296
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 15936 5176 15988 5228
rect 16580 5176 16632 5228
rect 17592 5176 17644 5228
rect 18512 5176 18564 5228
rect 19248 5176 19300 5228
rect 15660 5151 15712 5160
rect 15660 5117 15669 5151
rect 15669 5117 15703 5151
rect 15703 5117 15712 5151
rect 15660 5108 15712 5117
rect 16120 5108 16172 5160
rect 16948 5108 17000 5160
rect 17684 5108 17736 5160
rect 19156 5108 19208 5160
rect 20444 5176 20496 5228
rect 20904 5176 20956 5228
rect 20076 5151 20128 5160
rect 20076 5117 20085 5151
rect 20085 5117 20119 5151
rect 20119 5117 20128 5151
rect 20076 5108 20128 5117
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 11520 5040 11572 5092
rect 17960 5040 18012 5092
rect 18052 5040 18104 5092
rect 13268 4972 13320 5024
rect 13544 5015 13596 5024
rect 13544 4981 13553 5015
rect 13553 4981 13587 5015
rect 13587 4981 13596 5015
rect 13544 4972 13596 4981
rect 13912 5015 13964 5024
rect 13912 4981 13921 5015
rect 13921 4981 13955 5015
rect 13955 4981 13964 5015
rect 13912 4972 13964 4981
rect 14004 4972 14056 5024
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 16764 4972 16816 5024
rect 16856 4972 16908 5024
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 18604 4972 18656 5024
rect 18788 4972 18840 5024
rect 19156 4972 19208 5024
rect 19432 4972 19484 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2044 4768 2096 4820
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 6000 4768 6052 4820
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 6828 4768 6880 4820
rect 9588 4768 9640 4820
rect 10324 4811 10376 4820
rect 10324 4777 10333 4811
rect 10333 4777 10367 4811
rect 10367 4777 10376 4811
rect 10324 4768 10376 4777
rect 10508 4768 10560 4820
rect 5724 4700 5776 4752
rect 2964 4632 3016 4684
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 7288 4700 7340 4752
rect 8300 4700 8352 4752
rect 7472 4632 7524 4684
rect 8668 4700 8720 4752
rect 9680 4700 9732 4752
rect 12348 4768 12400 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 14372 4768 14424 4820
rect 18052 4768 18104 4820
rect 18420 4768 18472 4820
rect 18788 4768 18840 4820
rect 19984 4768 20036 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 10692 4675 10744 4684
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 2688 4564 2740 4616
rect 3332 4564 3384 4616
rect 3700 4607 3752 4616
rect 3700 4573 3709 4607
rect 3709 4573 3743 4607
rect 3743 4573 3752 4607
rect 3700 4564 3752 4573
rect 4712 4564 4764 4616
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 5724 4564 5776 4616
rect 6828 4564 6880 4616
rect 7748 4564 7800 4616
rect 8484 4564 8536 4616
rect 4068 4496 4120 4548
rect 10692 4641 10701 4675
rect 10701 4641 10735 4675
rect 10735 4641 10744 4675
rect 10692 4632 10744 4641
rect 11152 4632 11204 4684
rect 11980 4632 12032 4684
rect 17040 4700 17092 4752
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 13912 4632 13964 4684
rect 14096 4632 14148 4684
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 9220 4496 9272 4548
rect 10600 4564 10652 4616
rect 11060 4564 11112 4616
rect 11612 4564 11664 4616
rect 16212 4632 16264 4684
rect 16396 4632 16448 4684
rect 16948 4632 17000 4684
rect 18880 4675 18932 4684
rect 18880 4641 18889 4675
rect 18889 4641 18923 4675
rect 18923 4641 18932 4675
rect 18880 4632 18932 4641
rect 10140 4496 10192 4548
rect 11796 4496 11848 4548
rect 2780 4428 2832 4480
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 8208 4428 8260 4480
rect 10048 4428 10100 4480
rect 11060 4428 11112 4480
rect 12716 4428 12768 4480
rect 16028 4564 16080 4616
rect 16672 4564 16724 4616
rect 16856 4564 16908 4616
rect 13728 4428 13780 4480
rect 18512 4564 18564 4616
rect 18972 4607 19024 4616
rect 18972 4573 18981 4607
rect 18981 4573 19015 4607
rect 19015 4573 19024 4607
rect 18972 4564 19024 4573
rect 19616 4675 19668 4684
rect 19616 4641 19650 4675
rect 19650 4641 19668 4675
rect 19616 4632 19668 4641
rect 21272 4632 21324 4684
rect 22192 4632 22244 4684
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 4896 4224 4948 4276
rect 6736 4224 6788 4276
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 2780 4020 2832 4072
rect 3700 4020 3752 4072
rect 4068 4020 4120 4072
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 6828 4156 6880 4208
rect 7656 4224 7708 4276
rect 5724 4131 5776 4140
rect 4988 4020 5040 4072
rect 5448 4020 5500 4072
rect 5724 4097 5733 4131
rect 5733 4097 5767 4131
rect 5767 4097 5776 4131
rect 5724 4088 5776 4097
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 8668 4224 8720 4276
rect 11888 4224 11940 4276
rect 12164 4224 12216 4276
rect 18972 4224 19024 4276
rect 19616 4224 19668 4276
rect 9956 4156 10008 4208
rect 10232 4156 10284 4208
rect 11152 4156 11204 4208
rect 11796 4156 11848 4208
rect 6920 4020 6972 4072
rect 9772 4088 9824 4140
rect 10876 4088 10928 4140
rect 11612 4088 11664 4140
rect 13728 4156 13780 4208
rect 13912 4156 13964 4208
rect 8852 4020 8904 4072
rect 10140 4020 10192 4072
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 13544 4088 13596 4140
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15016 4131 15068 4140
rect 15016 4097 15025 4131
rect 15025 4097 15059 4131
rect 15059 4097 15068 4131
rect 15016 4088 15068 4097
rect 15936 4088 15988 4140
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 17316 4088 17368 4140
rect 12164 4020 12216 4072
rect 5356 3952 5408 4004
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 2872 3884 2924 3936
rect 3700 3884 3752 3936
rect 4620 3884 4672 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 8300 3952 8352 4004
rect 9496 3952 9548 4004
rect 13452 4020 13504 4072
rect 13912 4020 13964 4072
rect 16488 4020 16540 4072
rect 16672 4020 16724 4072
rect 16856 4020 16908 4072
rect 18972 4020 19024 4072
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 8944 3884 8996 3936
rect 9404 3884 9456 3936
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 10692 3884 10744 3936
rect 11152 3884 11204 3936
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 12532 3927 12584 3936
rect 11796 3884 11848 3893
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 18512 3952 18564 4004
rect 15568 3884 15620 3936
rect 16212 3884 16264 3936
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 18880 3884 18932 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3424 3680 3476 3732
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 2964 3612 3016 3664
rect 4528 3655 4580 3664
rect 2596 3544 2648 3596
rect 2688 3544 2740 3596
rect 3976 3544 4028 3596
rect 4528 3621 4537 3655
rect 4537 3621 4571 3655
rect 4571 3621 4580 3655
rect 4528 3612 4580 3621
rect 7748 3680 7800 3732
rect 9772 3680 9824 3732
rect 11796 3680 11848 3732
rect 12072 3680 12124 3732
rect 12532 3680 12584 3732
rect 14556 3680 14608 3732
rect 6736 3655 6788 3664
rect 6736 3621 6770 3655
rect 6770 3621 6788 3655
rect 6736 3612 6788 3621
rect 6828 3612 6880 3664
rect 7656 3612 7708 3664
rect 8116 3612 8168 3664
rect 5724 3544 5776 3596
rect 6184 3544 6236 3596
rect 8576 3544 8628 3596
rect 8944 3612 8996 3664
rect 11704 3612 11756 3664
rect 6460 3519 6512 3528
rect 4712 3408 4764 3460
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 2964 3340 3016 3392
rect 3516 3340 3568 3392
rect 8116 3408 8168 3460
rect 8668 3476 8720 3528
rect 9588 3544 9640 3596
rect 9772 3544 9824 3596
rect 10324 3544 10376 3596
rect 11060 3544 11112 3596
rect 12716 3612 12768 3664
rect 13544 3612 13596 3664
rect 13728 3655 13780 3664
rect 13728 3621 13762 3655
rect 13762 3621 13780 3655
rect 13728 3612 13780 3621
rect 16856 3680 16908 3732
rect 15844 3655 15896 3664
rect 15844 3621 15853 3655
rect 15853 3621 15887 3655
rect 15887 3621 15896 3655
rect 15844 3612 15896 3621
rect 16120 3612 16172 3664
rect 16488 3612 16540 3664
rect 17224 3655 17276 3664
rect 17224 3621 17233 3655
rect 17233 3621 17267 3655
rect 17267 3621 17276 3655
rect 17224 3612 17276 3621
rect 19524 3612 19576 3664
rect 17960 3587 18012 3596
rect 17960 3553 17969 3587
rect 17969 3553 18003 3587
rect 18003 3553 18012 3587
rect 17960 3544 18012 3553
rect 18512 3544 18564 3596
rect 12164 3519 12216 3528
rect 8576 3408 8628 3460
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 13084 3476 13136 3528
rect 13268 3519 13320 3528
rect 13268 3485 13277 3519
rect 13277 3485 13311 3519
rect 13311 3485 13320 3519
rect 13268 3476 13320 3485
rect 7564 3340 7616 3392
rect 12440 3408 12492 3460
rect 13176 3408 13228 3460
rect 16580 3476 16632 3528
rect 16856 3476 16908 3528
rect 17132 3476 17184 3528
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 16396 3408 16448 3460
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 19708 3476 19760 3528
rect 20536 3408 20588 3460
rect 10876 3340 10928 3392
rect 11704 3340 11756 3392
rect 11796 3340 11848 3392
rect 16304 3340 16356 3392
rect 18604 3340 18656 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 1952 3136 2004 3188
rect 572 3068 624 3120
rect 2596 3068 2648 3120
rect 3700 3136 3752 3188
rect 4712 3136 4764 3188
rect 4804 3068 4856 3120
rect 6184 3136 6236 3188
rect 6552 3136 6604 3188
rect 6460 3068 6512 3120
rect 8576 3136 8628 3188
rect 9588 3136 9640 3188
rect 10324 3179 10376 3188
rect 8944 3068 8996 3120
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 13084 3136 13136 3188
rect 17224 3136 17276 3188
rect 17316 3179 17368 3188
rect 17316 3145 17325 3179
rect 17325 3145 17359 3179
rect 17359 3145 17368 3179
rect 17316 3136 17368 3145
rect 17960 3136 18012 3188
rect 2964 3000 3016 3052
rect 10140 3000 10192 3052
rect 2044 2932 2096 2984
rect 4712 2932 4764 2984
rect 5724 2932 5776 2984
rect 6000 2932 6052 2984
rect 940 2864 992 2916
rect 2964 2864 3016 2916
rect 3148 2864 3200 2916
rect 3976 2864 4028 2916
rect 5172 2907 5224 2916
rect 204 2796 256 2848
rect 4896 2796 4948 2848
rect 5172 2873 5206 2907
rect 5206 2873 5224 2907
rect 5172 2864 5224 2873
rect 8668 2932 8720 2984
rect 8852 2932 8904 2984
rect 10876 2932 10928 2984
rect 11796 2975 11848 2984
rect 11796 2941 11805 2975
rect 11805 2941 11839 2975
rect 11839 2941 11848 2975
rect 11796 2932 11848 2941
rect 13728 3068 13780 3120
rect 16948 3068 17000 3120
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 13636 3000 13688 3052
rect 7748 2796 7800 2848
rect 8484 2796 8536 2848
rect 8852 2839 8904 2848
rect 8852 2805 8861 2839
rect 8861 2805 8895 2839
rect 8895 2805 8904 2839
rect 8852 2796 8904 2805
rect 8944 2796 8996 2848
rect 10692 2864 10744 2916
rect 10968 2864 11020 2916
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 11152 2796 11204 2848
rect 11888 2864 11940 2916
rect 13268 2864 13320 2916
rect 13084 2796 13136 2848
rect 13544 2932 13596 2984
rect 15568 3000 15620 3052
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 15844 2864 15896 2916
rect 16028 2932 16080 2984
rect 16764 2932 16816 2984
rect 16580 2864 16632 2916
rect 18972 3000 19024 3052
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 18696 2932 18748 2984
rect 17960 2864 18012 2916
rect 15660 2796 15712 2848
rect 16488 2796 16540 2848
rect 18604 2796 18656 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2872 2592 2924 2644
rect 4896 2592 4948 2644
rect 5356 2635 5408 2644
rect 4068 2524 4120 2576
rect 3332 2456 3384 2508
rect 3884 2456 3936 2508
rect 4896 2499 4948 2508
rect 4896 2465 4905 2499
rect 4905 2465 4939 2499
rect 4939 2465 4948 2499
rect 4896 2456 4948 2465
rect 3608 2388 3660 2440
rect 5080 2524 5132 2576
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 5632 2592 5684 2644
rect 6460 2592 6512 2644
rect 7380 2592 7432 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 8576 2592 8628 2644
rect 7564 2524 7616 2576
rect 8668 2567 8720 2576
rect 8668 2533 8677 2567
rect 8677 2533 8711 2567
rect 8711 2533 8720 2567
rect 8668 2524 8720 2533
rect 9496 2524 9548 2576
rect 5632 2456 5684 2508
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 7748 2456 7800 2508
rect 9680 2456 9732 2508
rect 10048 2592 10100 2644
rect 10416 2592 10468 2644
rect 12900 2592 12952 2644
rect 11060 2524 11112 2576
rect 13452 2524 13504 2576
rect 14004 2592 14056 2644
rect 11888 2499 11940 2508
rect 2412 2320 2464 2372
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 8852 2431 8904 2440
rect 8852 2397 8861 2431
rect 8861 2397 8895 2431
rect 8895 2397 8904 2431
rect 8852 2388 8904 2397
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 5540 2320 5592 2372
rect 8392 2320 8444 2372
rect 11888 2465 11897 2499
rect 11897 2465 11931 2499
rect 11931 2465 11940 2499
rect 11888 2456 11940 2465
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13084 2456 13136 2508
rect 13820 2456 13872 2508
rect 13360 2388 13412 2440
rect 13452 2388 13504 2440
rect 14740 2524 14792 2576
rect 16488 2592 16540 2644
rect 18512 2592 18564 2644
rect 18788 2635 18840 2644
rect 18788 2601 18797 2635
rect 18797 2601 18831 2635
rect 18831 2601 18840 2635
rect 18788 2592 18840 2601
rect 16764 2524 16816 2576
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 14464 2456 14516 2508
rect 15476 2456 15528 2508
rect 15752 2456 15804 2508
rect 16856 2456 16908 2508
rect 17040 2456 17092 2508
rect 17776 2524 17828 2576
rect 17592 2456 17644 2508
rect 18696 2499 18748 2508
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 19340 2456 19392 2508
rect 19800 2456 19852 2508
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 12532 2320 12584 2372
rect 3884 2252 3936 2304
rect 6644 2252 6696 2304
rect 8024 2252 8076 2304
rect 9404 2252 9456 2304
rect 11612 2252 11664 2304
rect 12164 2252 12216 2304
rect 13636 2320 13688 2372
rect 15108 2320 15160 2372
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 14372 2252 14424 2304
rect 16580 2320 16632 2372
rect 18512 2320 18564 2372
rect 17500 2295 17552 2304
rect 17500 2261 17509 2295
rect 17509 2261 17543 2295
rect 17543 2261 17552 2295
rect 17500 2252 17552 2261
rect 17592 2252 17644 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2044 2048 2096 2100
rect 4068 2048 4120 2100
rect 8208 2048 8260 2100
rect 6552 1980 6604 2032
rect 9312 1980 9364 2032
rect 5632 1912 5684 1964
rect 1308 1776 1360 1828
rect 8668 1776 8720 1828
rect 1676 1708 1728 1760
rect 5816 1708 5868 1760
rect 13268 1436 13320 1488
rect 13728 1436 13780 1488
rect 8392 1368 8444 1420
rect 9220 1368 9272 1420
rect 9956 1368 10008 1420
rect 10600 1368 10652 1420
rect 12900 1368 12952 1420
rect 14096 1368 14148 1420
rect 15844 1368 15896 1420
rect 17500 1368 17552 1420
rect 20720 892 20772 944
rect 21548 892 21600 944
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 938 22000 994 22800
rect 1306 22000 1362 22800
rect 1674 22000 1730 22800
rect 2042 22000 2098 22800
rect 2410 22000 2466 22800
rect 2778 22000 2834 22800
rect 3238 22000 3294 22800
rect 3606 22000 3662 22800
rect 3974 22000 4030 22800
rect 4342 22000 4398 22800
rect 4710 22000 4766 22800
rect 5078 22000 5134 22800
rect 5446 22000 5502 22800
rect 5906 22000 5962 22800
rect 6274 22000 6330 22800
rect 6642 22000 6698 22800
rect 7010 22000 7066 22800
rect 7378 22000 7434 22800
rect 7746 22000 7802 22800
rect 8114 22000 8170 22800
rect 8482 22000 8538 22800
rect 8942 22000 8998 22800
rect 9310 22000 9366 22800
rect 9678 22000 9734 22800
rect 10046 22000 10102 22800
rect 10414 22000 10470 22800
rect 10782 22000 10838 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12346 22000 12402 22800
rect 12714 22000 12770 22800
rect 13082 22000 13138 22800
rect 13450 22000 13506 22800
rect 13818 22000 13874 22800
rect 14186 22000 14242 22800
rect 14646 22000 14702 22800
rect 15014 22000 15070 22800
rect 15382 22000 15438 22800
rect 15750 22000 15806 22800
rect 16118 22000 16174 22800
rect 16486 22000 16542 22800
rect 16854 22000 16910 22800
rect 17314 22000 17370 22800
rect 17682 22000 17738 22800
rect 18050 22000 18106 22800
rect 18418 22000 18474 22800
rect 18786 22000 18842 22800
rect 18970 22672 19026 22681
rect 18970 22607 19026 22616
rect 216 19310 244 22000
rect 204 19304 256 19310
rect 204 19246 256 19252
rect 584 19242 612 22000
rect 572 19236 624 19242
rect 572 19178 624 19184
rect 952 18902 980 22000
rect 940 18896 992 18902
rect 940 18838 992 18844
rect 1320 18193 1348 22000
rect 1688 18970 1716 22000
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 2056 18766 2084 22000
rect 2424 18834 2452 22000
rect 2792 20754 2820 22000
rect 2792 20726 3188 20754
rect 2962 20632 3018 20641
rect 2962 20567 3018 20576
rect 2976 19281 3004 20567
rect 2962 19272 3018 19281
rect 2962 19207 3018 19216
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2044 18760 2096 18766
rect 1674 18728 1730 18737
rect 2044 18702 2096 18708
rect 1674 18663 1730 18672
rect 2872 18692 2924 18698
rect 1306 18184 1362 18193
rect 1306 18119 1362 18128
rect 1688 17882 1716 18663
rect 2872 18634 2924 18640
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2410 18456 2466 18465
rect 2410 18391 2466 18400
rect 1952 18352 2004 18358
rect 1950 18320 1952 18329
rect 2004 18320 2006 18329
rect 1950 18255 2006 18264
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 2148 17814 2176 18226
rect 2424 18154 2452 18391
rect 2412 18148 2464 18154
rect 2412 18090 2464 18096
rect 2688 18148 2740 18154
rect 2688 18090 2740 18096
rect 2136 17808 2188 17814
rect 2136 17750 2188 17756
rect 1950 17504 2006 17513
rect 1950 17439 2006 17448
rect 1964 17338 1992 17439
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2148 17218 2176 17750
rect 2700 17746 2728 18090
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2148 17202 2268 17218
rect 2148 17196 2280 17202
rect 2148 17190 2228 17196
rect 2228 17138 2280 17144
rect 1768 17128 1820 17134
rect 1582 17096 1638 17105
rect 1768 17070 1820 17076
rect 1582 17031 1638 17040
rect 1596 16794 1624 17031
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1398 16552 1454 16561
rect 1398 16487 1454 16496
rect 1412 16046 1440 16487
rect 1596 16250 1624 16623
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1780 15638 1808 17070
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1872 16794 1900 16934
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1950 16280 2006 16289
rect 1950 16215 2006 16224
rect 1964 16182 1992 16215
rect 1952 16176 2004 16182
rect 1952 16118 2004 16124
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 1308 15496 1360 15502
rect 1308 15438 1360 15444
rect 1582 15464 1638 15473
rect 1320 8809 1348 15438
rect 1582 15399 1638 15408
rect 1596 15162 1624 15399
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14385 1992 14758
rect 1950 14376 2006 14385
rect 1950 14311 2006 14320
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1780 13977 1808 14214
rect 1766 13968 1822 13977
rect 1766 13903 1822 13912
rect 2056 13870 2084 14894
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1596 12782 1624 12815
rect 1584 12776 1636 12782
rect 1688 12753 1716 13670
rect 1872 13462 1900 13806
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1766 13152 1822 13161
rect 1766 13087 1822 13096
rect 1780 12986 1808 13087
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1584 12718 1636 12724
rect 1674 12744 1730 12753
rect 1674 12679 1730 12688
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1596 11898 1624 12271
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11937 1716 12038
rect 1674 11928 1730 11937
rect 1584 11892 1636 11898
rect 1674 11863 1730 11872
rect 1584 11834 1636 11840
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11121 1440 11630
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1780 10810 1808 12582
rect 1872 11354 1900 13262
rect 1964 12986 1992 13330
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 2056 12594 2084 12650
rect 1964 12566 2084 12594
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1964 10266 1992 12566
rect 2148 12458 2176 15506
rect 2240 15473 2268 15982
rect 2424 15978 2452 17682
rect 2792 17134 2820 18566
rect 2884 18465 2912 18634
rect 2870 18456 2926 18465
rect 2870 18391 2926 18400
rect 2872 18352 2924 18358
rect 2872 18294 2924 18300
rect 2884 18222 2912 18294
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17814 2912 18022
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2688 16992 2740 16998
rect 2976 16946 3004 19110
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3068 18086 3096 18906
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 3160 17592 3188 20726
rect 3252 19258 3280 22000
rect 3252 19230 3556 19258
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3238 19000 3294 19009
rect 3238 18935 3240 18944
rect 3292 18935 3294 18944
rect 3240 18906 3292 18912
rect 3252 18698 3280 18906
rect 3436 18902 3464 19110
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3436 18601 3464 18702
rect 3422 18592 3478 18601
rect 3422 18527 3478 18536
rect 3240 18148 3292 18154
rect 3240 18090 3292 18096
rect 3068 17564 3188 17592
rect 3068 17066 3096 17564
rect 3252 17542 3280 18090
rect 3240 17536 3292 17542
rect 3160 17496 3240 17524
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 2688 16934 2740 16940
rect 2700 16810 2728 16934
rect 2792 16918 3004 16946
rect 2792 16810 2820 16918
rect 2700 16782 2820 16810
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2700 15910 2728 16594
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2792 15706 2820 16594
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2870 15872 2926 15881
rect 2870 15807 2926 15816
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2412 15496 2464 15502
rect 2226 15464 2282 15473
rect 2412 15438 2464 15444
rect 2226 15399 2282 15408
rect 2320 14816 2372 14822
rect 2318 14784 2320 14793
rect 2372 14784 2374 14793
rect 2318 14719 2374 14728
rect 2424 13433 2452 15438
rect 2778 15192 2834 15201
rect 2884 15162 2912 15807
rect 3068 15706 3096 16526
rect 3160 16522 3188 17496
rect 3240 17478 3292 17484
rect 3436 17270 3464 18527
rect 3332 17264 3384 17270
rect 3330 17232 3332 17241
rect 3424 17264 3476 17270
rect 3384 17232 3386 17241
rect 3424 17206 3476 17212
rect 3330 17167 3386 17176
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 2778 15127 2780 15136
rect 2832 15127 2834 15136
rect 2872 15156 2924 15162
rect 2780 15098 2832 15104
rect 2872 15098 2924 15104
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14550 2912 14894
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13569 2820 14214
rect 2778 13560 2834 13569
rect 2976 13546 3004 14758
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3068 14278 3096 14418
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 2884 13530 3004 13546
rect 2778 13495 2834 13504
rect 2872 13524 3004 13530
rect 2924 13518 3004 13524
rect 2872 13466 2924 13472
rect 2410 13424 2466 13433
rect 2410 13359 2466 13368
rect 2964 13388 3016 13394
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2056 12430 2176 12458
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1964 9722 1992 10066
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 2056 9602 2084 12430
rect 2332 12322 2360 12786
rect 2148 12306 2360 12322
rect 2136 12300 2360 12306
rect 2188 12294 2360 12300
rect 2136 12242 2188 12248
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 11898 2176 12038
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2148 10674 2176 11562
rect 2332 11558 2360 12294
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 11150 2360 11494
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 10062 2176 10610
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 1964 9574 2084 9602
rect 1306 8800 1362 8809
rect 1306 8735 1362 8744
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1504 7410 1532 8366
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1596 6866 1624 7822
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6254 1624 6802
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5778 1624 6190
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 572 3120 624 3126
rect 572 3062 624 3068
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 800 244 2790
rect 584 800 612 3062
rect 940 2916 992 2922
rect 940 2858 992 2864
rect 952 800 980 2858
rect 1308 1828 1360 1834
rect 1308 1770 1360 1776
rect 1320 800 1348 1770
rect 1676 1760 1728 1766
rect 1676 1702 1728 1708
rect 1688 800 1716 1702
rect 1780 921 1808 5782
rect 1964 3194 1992 9574
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2056 8498 2084 9454
rect 2240 9178 2268 10406
rect 2424 9994 2452 13359
rect 2964 13330 3016 13336
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2516 9518 2544 13194
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2608 12102 2636 12922
rect 2792 12442 2820 13262
rect 2976 12850 3004 13330
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11218 2636 12038
rect 3054 11656 3110 11665
rect 3054 11591 3110 11600
rect 2870 11248 2926 11257
rect 2596 11212 2648 11218
rect 2870 11183 2926 11192
rect 2596 11154 2648 11160
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10266 2820 10406
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2504 9512 2556 9518
rect 2792 9489 2820 9930
rect 2504 9454 2556 9460
rect 2778 9480 2834 9489
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2332 7002 2360 7142
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 2056 4826 2084 6870
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 5370 2176 6734
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2516 5166 2544 9454
rect 2778 9415 2834 9424
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 7177 2728 9318
rect 2884 8634 2912 11183
rect 3068 9602 3096 11591
rect 3252 11370 3280 14350
rect 3344 14278 3372 16934
rect 3436 16522 3464 17206
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 3436 16046 3464 16458
rect 3528 16130 3556 19230
rect 3620 18057 3648 22000
rect 3698 21040 3754 21049
rect 3698 20975 3754 20984
rect 3712 18329 3740 20975
rect 3988 19530 4016 22000
rect 4356 20398 4384 22000
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4068 20256 4120 20262
rect 4066 20224 4068 20233
rect 4120 20224 4122 20233
rect 4066 20159 4122 20168
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 3896 19502 4016 19530
rect 4264 19514 4292 19790
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4252 19508 4304 19514
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3804 18766 3832 18906
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3698 18320 3754 18329
rect 3698 18255 3754 18264
rect 3698 18184 3754 18193
rect 3698 18119 3700 18128
rect 3752 18119 3754 18128
rect 3700 18090 3752 18096
rect 3606 18048 3662 18057
rect 3606 17983 3662 17992
rect 3606 17912 3662 17921
rect 3606 17847 3662 17856
rect 3620 16794 3648 17847
rect 3896 17270 3924 19502
rect 4252 19450 4304 19456
rect 4620 19440 4672 19446
rect 3974 19408 4030 19417
rect 4620 19382 4672 19388
rect 3974 19343 4030 19352
rect 4252 19372 4304 19378
rect 3988 18873 4016 19343
rect 4252 19314 4304 19320
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18970 4108 19110
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 3974 18864 4030 18873
rect 3974 18799 4030 18808
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3988 18601 4016 18634
rect 3974 18592 4030 18601
rect 3974 18527 4030 18536
rect 4080 18290 4108 18770
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4068 17808 4120 17814
rect 4066 17776 4068 17785
rect 4120 17776 4122 17785
rect 4066 17711 4122 17720
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3700 17196 3752 17202
rect 3700 17138 3752 17144
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3712 16590 3740 17138
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3804 16726 3832 16934
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3712 16250 3740 16526
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3528 16102 4016 16130
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3436 15502 3464 15982
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3528 14600 3556 15846
rect 3896 15502 3924 15914
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3792 15088 3844 15094
rect 3790 15056 3792 15065
rect 3844 15056 3846 15065
rect 3790 14991 3846 15000
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 14618 3832 14758
rect 3436 14572 3556 14600
rect 3792 14612 3844 14618
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3344 12306 3372 13126
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3252 11342 3372 11370
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3160 10674 3188 11154
rect 3252 10810 3280 11222
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10062 3188 10610
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3160 9722 3188 9998
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 2976 9574 3096 9602
rect 2976 9382 3004 9574
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7546 2820 8230
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2686 7168 2742 7177
rect 2686 7103 2742 7112
rect 2792 6866 2820 7346
rect 2976 7290 3004 9046
rect 3068 8498 3096 9386
rect 3160 8974 3188 9658
rect 3252 9058 3280 10474
rect 3344 9178 3372 11342
rect 3436 10577 3464 14572
rect 3792 14554 3844 14560
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3528 13530 3556 14418
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3620 13530 3648 14350
rect 3896 13870 3924 15438
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3700 13796 3752 13802
rect 3700 13738 3752 13744
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3712 13258 3740 13738
rect 3896 13734 3924 13806
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3896 12986 3924 13670
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3528 12442 3556 12650
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3988 12322 4016 16102
rect 4080 16046 4108 17614
rect 4172 17338 4200 19178
rect 4264 18358 4292 19314
rect 4632 19174 4660 19382
rect 4620 19168 4672 19174
rect 4724 19145 4752 22000
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4816 19825 4844 19994
rect 4802 19816 4858 19825
rect 4802 19751 4858 19760
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4620 19110 4672 19116
rect 4710 19136 4766 19145
rect 4710 19071 4766 19080
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4252 18352 4304 18358
rect 4252 18294 4304 18300
rect 4264 17814 4292 18294
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 4342 18048 4398 18057
rect 4342 17983 4398 17992
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 4356 17524 4384 17983
rect 4448 17762 4476 18158
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4724 18057 4752 18090
rect 4710 18048 4766 18057
rect 4710 17983 4766 17992
rect 4816 17898 4844 19246
rect 5000 19174 5028 19246
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5000 18834 5028 19110
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 5000 18290 5028 18634
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4816 17882 4936 17898
rect 4816 17876 4948 17882
rect 4816 17870 4896 17876
rect 4896 17818 4948 17824
rect 4448 17734 4752 17762
rect 4528 17672 4580 17678
rect 4526 17640 4528 17649
rect 4580 17640 4582 17649
rect 4526 17575 4582 17584
rect 4264 17496 4384 17524
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4264 17082 4292 17496
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4172 17054 4292 17082
rect 4724 17066 4752 17734
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4528 17060 4580 17066
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14618 4108 14962
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 13870 4108 14350
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3528 12294 4016 12322
rect 3422 10568 3478 10577
rect 3422 10503 3478 10512
rect 3528 10266 3556 12294
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3712 11354 3740 11494
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3436 9110 3464 10066
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3424 9104 3476 9110
rect 3252 9030 3372 9058
rect 3424 9046 3476 9052
rect 3528 9042 3556 9998
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3068 8090 3096 8434
rect 3344 8430 3372 9030
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3332 8424 3384 8430
rect 3436 8401 3464 8774
rect 3332 8366 3384 8372
rect 3422 8392 3478 8401
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3160 7342 3188 8230
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7410 3280 7686
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 7336 3200 7342
rect 2976 7262 3096 7290
rect 3148 7278 3200 7284
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2792 6390 2820 6802
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2884 6304 2912 6598
rect 2976 6458 3004 7142
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2964 6316 3016 6322
rect 2884 6276 2964 6304
rect 2964 6258 3016 6264
rect 2976 5914 3004 6258
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2700 5545 2728 5714
rect 3068 5658 3096 7262
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 2976 5630 3096 5658
rect 2686 5536 2742 5545
rect 2686 5471 2742 5480
rect 2700 5234 2728 5471
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 4826 2268 4966
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2056 2990 2084 3878
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2332 2553 2360 4558
rect 2318 2544 2374 2553
rect 2318 2479 2374 2488
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 1766 912 1822 921
rect 1766 847 1822 856
rect 2056 800 2084 2042
rect 2424 800 2452 2314
rect 2516 1737 2544 5102
rect 2700 5030 2728 5170
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2700 4622 2728 4966
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2608 3602 2636 4082
rect 2792 4078 2820 4422
rect 2884 4146 2912 5034
rect 2976 4690 3004 5630
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5166 3096 5510
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2872 4140 2924 4146
rect 2924 4100 3004 4128
rect 2872 4082 2924 4088
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2700 3210 2728 3538
rect 2608 3182 2728 3210
rect 2608 3126 2636 3182
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2884 2650 2912 3878
rect 2976 3670 3004 4100
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3058 3004 3334
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2962 2952 3018 2961
rect 2962 2887 2964 2896
rect 3016 2887 3018 2896
rect 3148 2916 3200 2922
rect 2964 2858 3016 2864
rect 3148 2858 3200 2864
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2778 2544 2834 2553
rect 2778 2479 2834 2488
rect 2502 1728 2558 1737
rect 2502 1663 2558 1672
rect 2792 800 2820 2479
rect 3160 800 3188 2858
rect 3252 2145 3280 7142
rect 3344 4622 3372 8366
rect 3422 8327 3478 8336
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3436 7449 3464 7890
rect 3422 7440 3478 7449
rect 3422 7375 3424 7384
rect 3476 7375 3478 7384
rect 3424 7346 3476 7352
rect 3528 5914 3556 8978
rect 3620 8974 3648 11222
rect 3804 11098 3832 11562
rect 3896 11354 3924 11698
rect 3988 11694 4016 12106
rect 4172 11898 4200 17054
rect 4528 17002 4580 17008
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4264 16250 4292 16934
rect 4540 16794 4568 17002
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4816 16590 4844 17274
rect 4894 17232 4950 17241
rect 4894 17167 4950 17176
rect 4908 17134 4936 17167
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4816 15201 4844 16526
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4908 16114 4936 16458
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4896 15904 4948 15910
rect 4894 15872 4896 15881
rect 4948 15872 4950 15881
rect 4894 15807 4950 15816
rect 4802 15192 4858 15201
rect 4802 15127 4858 15136
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4816 14550 4844 14962
rect 4896 14884 4948 14890
rect 4896 14826 4948 14832
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4816 14074 4844 14486
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4908 13530 4936 14826
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4724 12322 4752 13330
rect 5000 12374 5028 16662
rect 5092 13190 5120 22000
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5184 18902 5212 19926
rect 5460 19258 5488 22000
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5552 19514 5580 19858
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5460 19230 5580 19258
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5276 18902 5304 19110
rect 5460 18970 5488 19110
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5276 17814 5304 18702
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5368 17649 5396 18770
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5354 17640 5410 17649
rect 5354 17575 5410 17584
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5184 17202 5212 17478
rect 5264 17264 5316 17270
rect 5264 17206 5316 17212
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5184 15706 5212 16186
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4804 12368 4856 12374
rect 4724 12316 4804 12322
rect 4724 12310 4856 12316
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4724 12294 4844 12310
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 4618 11656 4674 11665
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3712 11070 3832 11098
rect 3712 10198 3740 11070
rect 3790 10840 3846 10849
rect 3790 10775 3792 10784
rect 3844 10775 3846 10784
rect 3792 10746 3844 10752
rect 3790 10704 3846 10713
rect 3896 10674 3924 11290
rect 3988 11218 4016 11630
rect 4618 11591 4674 11600
rect 4632 11558 4660 11591
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4160 11552 4212 11558
rect 4344 11552 4396 11558
rect 4160 11494 4212 11500
rect 4264 11512 4344 11540
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3988 11082 4016 11154
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3988 10742 4016 11018
rect 4080 10849 4108 11494
rect 4172 11354 4200 11494
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3790 10639 3846 10648
rect 3884 10668 3936 10674
rect 3804 10470 3832 10639
rect 3884 10610 3936 10616
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 8090 3648 8910
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3620 7546 3648 7822
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3712 7342 3740 10134
rect 3804 8294 3832 10202
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3896 9450 3924 9998
rect 3988 9926 4016 10678
rect 4264 10606 4292 11512
rect 4344 11494 4396 11500
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4252 10600 4304 10606
rect 4436 10600 4488 10606
rect 4252 10542 4304 10548
rect 4434 10568 4436 10577
rect 4488 10568 4490 10577
rect 4724 10538 4752 12038
rect 4434 10503 4490 10512
rect 4712 10532 4764 10538
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 10033 4108 10202
rect 4344 10192 4396 10198
rect 4264 10152 4344 10180
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 4264 9722 4292 10152
rect 4344 10134 4396 10140
rect 4448 9908 4476 10503
rect 4712 10474 4764 10480
rect 4448 9880 4752 9908
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3804 7478 3832 8026
rect 3896 8022 3924 8434
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3528 5273 3556 5306
rect 3514 5264 3570 5273
rect 3514 5199 3570 5208
rect 3620 5098 3648 6870
rect 3712 6746 3740 7278
rect 3792 7200 3844 7206
rect 3790 7168 3792 7177
rect 3844 7168 3846 7177
rect 3790 7103 3846 7112
rect 3804 6882 3832 7103
rect 3896 7002 3924 7414
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3804 6854 3924 6882
rect 3988 6866 4016 8298
rect 4080 7954 4108 9386
rect 4724 8906 4752 9880
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4618 8392 4674 8401
rect 4618 8327 4674 8336
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4068 7744 4120 7750
rect 4066 7712 4068 7721
rect 4120 7712 4122 7721
rect 4066 7647 4122 7656
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4080 7313 4108 7482
rect 4264 7426 4292 7890
rect 4632 7732 4660 8327
rect 4632 7704 4752 7732
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4436 7472 4488 7478
rect 4264 7410 4384 7426
rect 4436 7414 4488 7420
rect 4264 7404 4396 7410
rect 4264 7398 4344 7404
rect 4344 7346 4396 7352
rect 4066 7304 4122 7313
rect 4066 7239 4122 7248
rect 4356 6866 4384 7346
rect 4448 7274 4476 7414
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 3712 6718 3832 6746
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3712 5166 3740 5646
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3344 3097 3372 4558
rect 3436 3738 3464 4626
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4078 3740 4558
rect 3700 4072 3752 4078
rect 3620 4032 3700 4060
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3330 3088 3386 3097
rect 3330 3023 3386 3032
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3238 2136 3294 2145
rect 3238 2071 3294 2080
rect 3344 1329 3372 2450
rect 3330 1320 3386 1329
rect 3330 1255 3386 1264
rect 3528 800 3556 3334
rect 3620 2446 3648 4032
rect 3700 4014 3752 4020
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3712 3194 3740 3878
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3804 513 3832 6718
rect 3896 2514 3924 6854
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4066 6488 4122 6497
rect 3976 6452 4028 6458
rect 4388 6480 4684 6500
rect 4066 6423 4122 6432
rect 3976 6394 4028 6400
rect 3988 5681 4016 6394
rect 4080 6390 4108 6423
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4066 6080 4122 6089
rect 4066 6015 4122 6024
rect 4080 5914 4108 6015
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3974 5672 4030 5681
rect 3974 5607 4030 5616
rect 4080 5216 4108 5714
rect 4172 5370 4200 6190
rect 4264 5545 4292 6258
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4632 6089 4660 6190
rect 4618 6080 4674 6089
rect 4618 6015 4674 6024
rect 4724 5896 4752 7704
rect 4632 5868 4752 5896
rect 4632 5658 4660 5868
rect 4712 5772 4764 5778
rect 4816 5760 4844 12294
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11665 5028 11698
rect 4986 11656 5042 11665
rect 4986 11591 5042 11600
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5000 10538 5028 10950
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 9897 5028 10474
rect 4986 9888 5042 9897
rect 4986 9823 5042 9832
rect 5092 9489 5120 11834
rect 5184 10452 5212 14214
rect 5276 12866 5304 17206
rect 5460 16658 5488 17818
rect 5552 17610 5580 19230
rect 5644 18698 5672 19654
rect 5828 18970 5856 19654
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5920 18850 5948 22000
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 5998 19000 6054 19009
rect 5998 18935 6000 18944
rect 6052 18935 6054 18944
rect 6000 18906 6052 18912
rect 5920 18822 6040 18850
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5920 18426 5948 18702
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5368 15201 5396 16390
rect 5552 15978 5580 17206
rect 5644 17134 5672 18022
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5736 16794 5764 18158
rect 6012 17649 6040 18822
rect 6104 18766 6132 19178
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 5998 17640 6054 17649
rect 5998 17575 6054 17584
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5920 16590 5948 17478
rect 6012 17202 6040 17478
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5552 15366 5580 15914
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5354 15192 5410 15201
rect 5354 15127 5410 15136
rect 5644 14521 5672 16526
rect 5814 15464 5870 15473
rect 5814 15399 5870 15408
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5630 14512 5686 14521
rect 5630 14447 5686 14456
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5460 13326 5488 14010
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5368 12986 5396 13262
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5276 12838 5396 12866
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5276 10810 5304 11086
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5262 10704 5318 10713
rect 5262 10639 5318 10648
rect 5276 10606 5304 10639
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5264 10464 5316 10470
rect 5184 10424 5264 10452
rect 5264 10406 5316 10412
rect 5170 10296 5226 10305
rect 5170 10231 5226 10240
rect 5078 9480 5134 9489
rect 5078 9415 5134 9424
rect 5092 8401 5120 9415
rect 5078 8392 5134 8401
rect 5078 8327 5134 8336
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4764 5732 4844 5760
rect 4712 5714 4764 5720
rect 4908 5658 4936 6938
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 5000 5953 5028 6870
rect 5092 6633 5120 8230
rect 5184 6934 5212 10231
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5078 6624 5134 6633
rect 5078 6559 5134 6568
rect 4986 5944 5042 5953
rect 4986 5879 5042 5888
rect 5092 5846 5120 6559
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4632 5630 4752 5658
rect 4250 5536 4306 5545
rect 4250 5471 4306 5480
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4250 5264 4306 5273
rect 4080 5188 4200 5216
rect 4250 5199 4306 5208
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4080 4865 4108 5034
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4080 4457 4108 4490
rect 4066 4448 4122 4457
rect 4066 4383 4122 4392
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3988 2922 4016 3538
rect 4080 3369 4108 4014
rect 4066 3360 4122 3369
rect 4066 3295 4122 3304
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 800 3924 2246
rect 4080 2106 4108 2518
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 3790 504 3846 513
rect 3790 439 3846 448
rect 3882 0 3938 800
rect 4172 241 4200 5188
rect 4264 800 4292 5199
rect 4724 4622 4752 5630
rect 4816 5630 4936 5658
rect 5184 5642 5212 6258
rect 5276 5658 5304 10406
rect 5368 5778 5396 12838
rect 5460 11014 5488 13126
rect 5552 12986 5580 13738
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5644 12832 5672 14447
rect 5736 13530 5764 14758
rect 5828 13954 5856 15399
rect 6104 15178 6132 17546
rect 6288 17354 6316 22000
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6472 17678 6500 18226
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6288 17326 6408 17354
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 6196 16794 6224 17002
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6380 16425 6408 17326
rect 6366 16416 6422 16425
rect 6366 16351 6422 16360
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6104 15150 6316 15178
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5920 14074 5948 14962
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 14618 6040 14758
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6104 14074 6132 14350
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 5828 13926 5948 13954
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5828 13530 5856 13806
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5920 13410 5948 13926
rect 5828 13382 5948 13410
rect 6104 13394 6132 14010
rect 6092 13388 6144 13394
rect 5724 12844 5776 12850
rect 5644 12804 5724 12832
rect 5724 12786 5776 12792
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10198 5488 10610
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5552 10044 5580 12378
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11354 5672 11494
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5736 11234 5764 12650
rect 5644 11206 5764 11234
rect 5644 10169 5672 11206
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5630 10160 5686 10169
rect 5630 10095 5686 10104
rect 5460 10016 5580 10044
rect 5460 7188 5488 10016
rect 5644 9058 5672 10095
rect 5736 9178 5764 10406
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5644 9030 5764 9058
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5552 8090 5580 8434
rect 5736 8378 5764 9030
rect 5644 8350 5764 8378
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5552 7449 5580 8026
rect 5538 7440 5594 7449
rect 5538 7375 5594 7384
rect 5460 7160 5580 7188
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5172 5636 5224 5642
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4526 4176 4582 4185
rect 4526 4111 4582 4120
rect 4540 3670 4568 4111
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 3738 4660 3878
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4724 3194 4752 3402
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4724 2990 4752 3130
rect 4816 3126 4844 5630
rect 5276 5630 5396 5658
rect 5172 5578 5224 5584
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5000 4570 5028 5306
rect 5092 5234 5120 5510
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5184 5030 5212 5170
rect 5276 5166 5304 5510
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5368 4865 5396 5630
rect 5354 4856 5410 4865
rect 5354 4791 5410 4800
rect 5000 4542 5120 4570
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4908 4146 4936 4218
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5000 4078 5028 4422
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4986 3768 5042 3777
rect 4986 3703 5042 3712
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4908 2650 4936 2790
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4894 2544 4950 2553
rect 4894 2479 4896 2488
rect 4948 2479 4950 2488
rect 4896 2450 4948 2456
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4618 2000 4674 2009
rect 4618 1935 4674 1944
rect 4632 800 4660 1935
rect 5000 800 5028 3703
rect 5092 2582 5120 4542
rect 5460 4078 5488 6054
rect 5552 5710 5580 7160
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5644 5522 5672 8350
rect 5828 7449 5856 13382
rect 6092 13330 6144 13336
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 9994 5948 10406
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 6012 9722 6040 10610
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6012 9518 6040 9658
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6012 8974 6040 9318
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 8090 5948 8230
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5814 7440 5870 7449
rect 5814 7375 5870 7384
rect 5828 6254 5856 7375
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5552 5494 5672 5522
rect 5552 4468 5580 5494
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5644 4622 5672 5170
rect 5736 4758 5764 6054
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5724 4616 5776 4622
rect 5828 4593 5856 5646
rect 5920 4706 5948 7754
rect 6012 6866 6040 8910
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5998 6488 6054 6497
rect 5998 6423 6054 6432
rect 6012 4826 6040 6423
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5920 4678 6040 4706
rect 5724 4558 5776 4564
rect 5814 4584 5870 4593
rect 5552 4440 5672 4468
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5184 2446 5212 2858
rect 5368 2650 5396 3946
rect 5540 3936 5592 3942
rect 5446 3904 5502 3913
rect 5540 3878 5592 3884
rect 5446 3839 5502 3848
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5460 898 5488 3839
rect 5552 2378 5580 3878
rect 5644 3777 5672 4440
rect 5736 4146 5764 4558
rect 5814 4519 5870 4528
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 4185 5856 4422
rect 5906 4312 5962 4321
rect 5906 4247 5962 4256
rect 5814 4176 5870 4185
rect 5724 4140 5776 4146
rect 5814 4111 5870 4120
rect 5724 4082 5776 4088
rect 5630 3768 5686 3777
rect 5630 3703 5686 3712
rect 5736 3602 5764 4082
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5644 2514 5672 2586
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 5644 1970 5672 2450
rect 5632 1964 5684 1970
rect 5632 1906 5684 1912
rect 5368 870 5488 898
rect 5368 800 5396 870
rect 5736 800 5764 2926
rect 5816 2508 5868 2514
rect 5920 2496 5948 4247
rect 6012 2990 6040 4678
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6104 2904 6132 13194
rect 6196 12481 6224 15030
rect 6288 14822 6316 15150
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6288 14414 6316 14758
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6380 14090 6408 16186
rect 6472 15586 6500 17614
rect 6656 17105 6684 22000
rect 7024 20602 7052 22000
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7392 20482 7420 22000
rect 7760 20754 7788 22000
rect 7024 20454 7420 20482
rect 7484 20726 7788 20754
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 17338 6868 19858
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6642 17096 6698 17105
rect 7024 17082 7052 20454
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 6642 17031 6698 17040
rect 6748 17054 7052 17082
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6656 16794 6684 16934
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6564 15706 6592 16594
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6656 15910 6684 16526
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6472 15570 6592 15586
rect 6472 15564 6604 15570
rect 6472 15558 6552 15564
rect 6552 15506 6604 15512
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 14618 6500 15438
rect 6564 15008 6592 15506
rect 6656 15502 6684 15846
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6644 15020 6696 15026
rect 6564 14980 6644 15008
rect 6644 14962 6696 14968
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6380 14062 6500 14090
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6288 13326 6316 13670
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6380 13172 6408 13942
rect 6288 13144 6408 13172
rect 6182 12472 6238 12481
rect 6182 12407 6238 12416
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11830 6224 12242
rect 6288 12102 6316 13144
rect 6472 13002 6500 14062
rect 6564 13326 6592 14350
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6380 12974 6500 13002
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6196 11150 6224 11766
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 9178 6224 10406
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 9586 6316 10066
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6182 8800 6238 8809
rect 6182 8735 6238 8744
rect 6196 7818 6224 8735
rect 6274 8392 6330 8401
rect 6274 8327 6330 8336
rect 6288 7954 6316 8327
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6274 7576 6330 7585
rect 6274 7511 6330 7520
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6196 6322 6224 6598
rect 6288 6458 6316 7511
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6184 6316 6236 6322
rect 6236 6276 6316 6304
rect 6184 6258 6236 6264
rect 6184 5840 6236 5846
rect 6182 5808 6184 5817
rect 6236 5808 6238 5817
rect 6182 5743 6238 5752
rect 6288 5658 6316 6276
rect 6380 5914 6408 12974
rect 6564 12850 6592 13262
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6550 12336 6606 12345
rect 6550 12271 6606 12280
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6472 8809 6500 11562
rect 6458 8800 6514 8809
rect 6458 8735 6514 8744
rect 6458 8528 6514 8537
rect 6458 8463 6514 8472
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6196 5630 6316 5658
rect 6196 5234 6224 5630
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 4826 6224 4966
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6288 4690 6316 5510
rect 6380 5302 6408 5850
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6472 5012 6500 8463
rect 6564 7313 6592 12271
rect 6656 11608 6684 14962
rect 6748 14550 6776 17054
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6932 15434 6960 16934
rect 7116 16810 7144 20266
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7300 17882 7328 19858
rect 7484 18578 7512 20726
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 7392 18550 7512 18578
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7024 16782 7144 16810
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6748 14385 6776 14486
rect 6734 14376 6790 14385
rect 6734 14311 6790 14320
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6748 12918 6776 13806
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6840 12986 6868 13330
rect 6918 13288 6974 13297
rect 6918 13223 6920 13232
rect 6972 13223 6974 13232
rect 6920 13194 6972 13200
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6932 12374 6960 12854
rect 7024 12617 7052 16782
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7208 15162 7236 15506
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14793 7328 14894
rect 7286 14784 7342 14793
rect 7286 14719 7342 14728
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7116 13870 7144 14418
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7208 12918 7236 14554
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7010 12608 7066 12617
rect 7010 12543 7066 12552
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6748 11937 6776 12310
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6734 11928 6790 11937
rect 6734 11863 6790 11872
rect 6840 11762 6868 12038
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6736 11620 6788 11626
rect 6656 11580 6736 11608
rect 6736 11562 6788 11568
rect 6748 10996 6776 11562
rect 6826 11248 6882 11257
rect 6826 11183 6828 11192
rect 6880 11183 6882 11192
rect 6828 11154 6880 11160
rect 6932 11150 6960 12310
rect 7116 11898 7144 12650
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7102 11792 7158 11801
rect 7102 11727 7158 11736
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6748 10968 6960 10996
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6656 10266 6684 10474
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6748 9450 6776 10134
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6748 8974 6776 9386
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 9178 6868 9318
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6656 8786 6684 8842
rect 6828 8832 6880 8838
rect 6826 8800 6828 8809
rect 6932 8820 6960 10968
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 9110 7052 10406
rect 7116 9217 7144 11727
rect 7208 11082 7236 12718
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7102 9208 7158 9217
rect 7102 9143 7158 9152
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7012 8832 7064 8838
rect 6880 8800 6882 8809
rect 6656 8758 6776 8786
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6564 6118 6592 7239
rect 6656 6730 6684 8366
rect 6748 6746 6776 8758
rect 6932 8792 7012 8820
rect 7012 8774 7064 8780
rect 6826 8735 6882 8744
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6840 8022 6868 8434
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6840 7478 6868 7958
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6644 6724 6696 6730
rect 6748 6718 6868 6746
rect 6644 6666 6696 6672
rect 6736 6656 6788 6662
rect 6656 6604 6736 6610
rect 6656 6598 6788 6604
rect 6656 6582 6776 6598
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 5137 6592 5714
rect 6550 5128 6606 5137
rect 6550 5063 6606 5072
rect 6552 5024 6604 5030
rect 6472 4984 6552 5012
rect 6552 4966 6604 4972
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6196 3194 6224 3538
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6472 3126 6500 3470
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6564 2938 6592 3130
rect 6472 2910 6592 2938
rect 6104 2876 6224 2904
rect 5868 2468 5948 2496
rect 5816 2450 5868 2456
rect 5828 1766 5856 2450
rect 5816 1760 5868 1766
rect 5816 1702 5868 1708
rect 6196 800 6224 2876
rect 6472 2650 6500 2910
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6656 2310 6684 6582
rect 6736 6384 6788 6390
rect 6734 6352 6736 6361
rect 6788 6352 6790 6361
rect 6734 6287 6790 6296
rect 6734 6216 6790 6225
rect 6734 6151 6790 6160
rect 6748 5846 6776 6151
rect 6840 5846 6868 6718
rect 6932 5914 6960 8502
rect 7024 7002 7052 8774
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5234 6776 5646
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6748 4729 6776 5170
rect 6840 4826 6868 5170
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6734 4720 6790 4729
rect 6734 4655 6790 4664
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6748 3670 6776 4218
rect 6840 4214 6868 4558
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6932 4078 6960 5850
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 7024 3913 7052 6666
rect 7010 3904 7066 3913
rect 7010 3839 7066 3848
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6840 2553 6868 3606
rect 7116 3097 7144 8978
rect 7208 7936 7236 10746
rect 7300 8634 7328 14350
rect 7392 12442 7420 18550
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7484 16658 7512 17138
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7484 15366 7512 15438
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 15094 7512 15302
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7484 14414 7512 15030
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7576 12866 7604 20538
rect 8128 20330 8156 22000
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7760 19174 7788 19790
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7668 18766 7696 19110
rect 7760 18952 7788 19110
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7760 18924 7880 18952
rect 7852 18834 7880 18924
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7668 16726 7696 18702
rect 7852 18290 7880 18770
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17882 8248 19858
rect 8496 17921 8524 22000
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18290 8616 19110
rect 8680 18630 8708 19178
rect 8772 18902 8800 19178
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8680 18290 8708 18566
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8482 17912 8538 17921
rect 8208 17876 8260 17882
rect 8482 17847 8538 17856
rect 8208 17818 8260 17824
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7668 16046 7696 16662
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7668 14618 7696 15982
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7668 13802 7696 14418
rect 7760 14278 7788 17614
rect 8128 17202 8156 17682
rect 8484 17672 8536 17678
rect 8588 17649 8616 17682
rect 8680 17678 8708 18226
rect 8772 18086 8800 18838
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8668 17672 8720 17678
rect 8484 17614 8536 17620
rect 8574 17640 8630 17649
rect 8496 17338 8524 17614
rect 8668 17614 8720 17620
rect 8574 17575 8630 17584
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8128 15960 8156 16390
rect 8220 16250 8248 16594
rect 8680 16454 8708 17614
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8772 17105 8800 17478
rect 8758 17096 8814 17105
rect 8758 17031 8814 17040
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8772 16697 8800 16934
rect 8758 16688 8814 16697
rect 8758 16623 8814 16632
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8758 16416 8814 16425
rect 8758 16351 8814 16360
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8128 15932 8248 15960
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 7930 15464 7986 15473
rect 7930 15399 7986 15408
rect 7944 14958 7972 15399
rect 8036 15162 8064 15574
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8116 14544 8168 14550
rect 7944 14504 8116 14532
rect 7944 14346 7972 14504
rect 8116 14486 8168 14492
rect 8220 14482 8248 15932
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8482 15464 8538 15473
rect 8404 14958 8432 15438
rect 8482 15399 8538 15408
rect 8496 15026 8524 15399
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8484 14816 8536 14822
rect 8390 14784 8446 14793
rect 8484 14758 8536 14764
rect 8390 14719 8446 14728
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7668 12986 7696 13738
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8220 13512 8248 13670
rect 8128 13484 8248 13512
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7472 12844 7524 12850
rect 7576 12838 7696 12866
rect 7472 12786 7524 12792
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 10810 7420 12242
rect 7484 12170 7512 12786
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7472 11076 7524 11082
rect 7576 11064 7604 12718
rect 7668 12209 7696 12838
rect 7654 12200 7710 12209
rect 7654 12135 7710 12144
rect 7654 12064 7710 12073
rect 7654 11999 7710 12008
rect 7524 11036 7604 11064
rect 7472 11018 7524 11024
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7392 9178 7420 10406
rect 7484 10266 7512 10406
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7472 10056 7524 10062
rect 7470 10024 7472 10033
rect 7524 10024 7526 10033
rect 7470 9959 7526 9968
rect 7470 9888 7526 9897
rect 7470 9823 7526 9832
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7484 8945 7512 9823
rect 7576 9518 7604 11036
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7470 8936 7526 8945
rect 7470 8871 7526 8880
rect 7576 8786 7604 9046
rect 7392 8758 7604 8786
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7208 7908 7328 7936
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7478 7236 7754
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7208 6934 7236 7210
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7208 6798 7236 6870
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7194 5944 7250 5953
rect 7194 5879 7250 5888
rect 7208 5778 7236 5879
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7300 5658 7328 7908
rect 7208 5630 7328 5658
rect 7102 3088 7158 3097
rect 7102 3023 7158 3032
rect 7208 2972 7236 5630
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5234 7328 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7286 4856 7342 4865
rect 7286 4791 7342 4800
rect 7300 4758 7328 4791
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7392 4604 7420 8758
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 6730 7512 8298
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 8090 7604 8230
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7562 7984 7618 7993
rect 7562 7919 7564 7928
rect 7616 7919 7618 7928
rect 7564 7890 7616 7896
rect 7668 7562 7696 11999
rect 7760 11898 7788 13262
rect 8128 13161 8156 13484
rect 8404 13462 8432 14719
rect 8496 14657 8524 14758
rect 8482 14648 8538 14657
rect 8482 14583 8538 14592
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8114 13152 8170 13161
rect 8114 13087 8170 13096
rect 8128 12782 8156 13087
rect 8220 12986 8248 13330
rect 8392 13320 8444 13326
rect 8444 13280 8524 13308
rect 8392 13262 8444 13268
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8220 12238 8248 12582
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7760 11200 7788 11834
rect 7852 11762 7880 12106
rect 8312 11898 8340 13194
rect 8390 12744 8446 12753
rect 8390 12679 8446 12688
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7840 11212 7892 11218
rect 7760 11172 7840 11200
rect 7840 11154 7892 11160
rect 8298 10568 8354 10577
rect 8298 10503 8354 10512
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7748 10056 7800 10062
rect 8220 10033 8248 10406
rect 7748 9998 7800 10004
rect 8206 10024 8262 10033
rect 7760 8430 7788 9998
rect 8206 9959 8262 9968
rect 8312 9722 8340 10503
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8298 9616 8354 9625
rect 8298 9551 8354 9560
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7944 8634 7972 8842
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8128 8498 8156 8774
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 8114 8392 8170 8401
rect 7576 7534 7696 7562
rect 7576 7342 7604 7534
rect 7760 7478 7788 8366
rect 8220 8378 8248 9318
rect 8312 9042 8340 9551
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8298 8664 8354 8673
rect 8298 8599 8354 8608
rect 8312 8401 8340 8599
rect 8170 8350 8248 8378
rect 8114 8327 8170 8336
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7562 6896 7618 6905
rect 7668 6866 7696 7142
rect 7562 6831 7618 6840
rect 7656 6860 7708 6866
rect 7576 6730 7604 6831
rect 7656 6802 7708 6808
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7760 6458 7788 7414
rect 7852 7410 7880 7822
rect 7930 7712 7986 7721
rect 7930 7647 7986 7656
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7944 7274 7972 7647
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 8128 7188 8156 7414
rect 8220 7342 8248 8350
rect 8298 8392 8354 8401
rect 8298 8327 8354 8336
rect 8404 8294 8432 12679
rect 8496 12646 8524 13280
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8482 12472 8538 12481
rect 8482 12407 8538 12416
rect 8496 12306 8524 12407
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8496 10198 8524 11834
rect 8588 11098 8616 15846
rect 8680 12753 8708 15982
rect 8772 13530 8800 16351
rect 8864 15706 8892 18838
rect 8956 17270 8984 22000
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8850 15328 8906 15337
rect 8850 15263 8906 15272
rect 8864 15026 8892 15263
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8864 14618 8892 14962
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8666 12744 8722 12753
rect 8666 12679 8722 12688
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11694 8708 12038
rect 8772 11762 8800 13126
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8864 11286 8892 14214
rect 8956 14090 8984 16934
rect 9048 14278 9076 20334
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9140 18193 9168 19110
rect 9232 18834 9260 19314
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9232 18698 9260 18770
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9126 18184 9182 18193
rect 9126 18119 9182 18128
rect 9232 17202 9260 18634
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9232 16590 9260 17138
rect 9128 16584 9180 16590
rect 9126 16552 9128 16561
rect 9220 16584 9272 16590
rect 9180 16552 9182 16561
rect 9220 16526 9272 16532
rect 9126 16487 9182 16496
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 8956 14062 9076 14090
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8956 11898 8984 12242
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9048 11778 9076 14062
rect 9140 11898 9168 15506
rect 9324 15042 9352 22000
rect 9692 19446 9720 22000
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9784 19718 9812 19994
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18970 9536 19110
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9416 18222 9444 18566
rect 9600 18222 9628 18702
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 18034 9720 18158
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9600 18006 9720 18034
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16114 9444 16458
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9402 15192 9458 15201
rect 9402 15127 9458 15136
rect 9232 15014 9352 15042
rect 9232 13410 9260 15014
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 9324 14346 9352 14826
rect 9416 14414 9444 15127
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9232 13382 9352 13410
rect 9220 13320 9272 13326
rect 9324 13297 9352 13382
rect 9220 13262 9272 13268
rect 9310 13288 9366 13297
rect 9232 13161 9260 13262
rect 9310 13223 9366 13232
rect 9218 13152 9274 13161
rect 9218 13087 9274 13096
rect 9232 12850 9260 13087
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9232 12238 9260 12786
rect 9324 12617 9352 13223
rect 9310 12608 9366 12617
rect 9310 12543 9366 12552
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9048 11750 9352 11778
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8956 11150 8984 11494
rect 8944 11144 8996 11150
rect 8588 11070 8800 11098
rect 8944 11086 8996 11092
rect 8574 10840 8630 10849
rect 8574 10775 8630 10784
rect 8588 10470 8616 10775
rect 8668 10600 8720 10606
rect 8666 10568 8668 10577
rect 8720 10568 8722 10577
rect 8666 10503 8722 10512
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8666 10432 8722 10441
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8588 10033 8616 10406
rect 8666 10367 8722 10376
rect 8574 10024 8630 10033
rect 8574 9959 8630 9968
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9654 8524 9862
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8574 9208 8630 9217
rect 8574 9143 8630 9152
rect 8588 9110 8616 9143
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8680 8838 8708 10367
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8480 8708 8774
rect 8496 8452 8708 8480
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8128 7160 8248 7188
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8220 7041 8248 7160
rect 8206 7032 8262 7041
rect 8206 6967 8262 6976
rect 8024 6928 8076 6934
rect 7852 6876 8024 6882
rect 7852 6870 8076 6876
rect 7852 6866 8064 6870
rect 7840 6860 8064 6866
rect 7892 6854 8064 6860
rect 7840 6802 7892 6808
rect 7932 6792 7984 6798
rect 7930 6760 7932 6769
rect 7984 6760 7986 6769
rect 7930 6695 7986 6704
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7484 5273 7512 6394
rect 7760 6304 7788 6394
rect 7760 6276 7880 6304
rect 7852 6186 7880 6276
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7760 5914 7788 6122
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7576 5574 7604 5850
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7760 5681 7788 5714
rect 7746 5672 7802 5681
rect 7746 5607 7802 5616
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7470 5264 7526 5273
rect 7470 5199 7472 5208
rect 7524 5199 7526 5208
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 7472 5170 7524 5176
rect 7484 5139 7512 5170
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 6932 2944 7236 2972
rect 7300 4576 7420 4604
rect 6826 2544 6882 2553
rect 6826 2479 6882 2488
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6564 800 6592 1974
rect 6932 800 6960 2944
rect 7300 800 7328 4576
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 2650 7420 3878
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7484 2428 7512 4626
rect 7576 3398 7604 4966
rect 7668 4282 7696 5199
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8220 4808 8248 5850
rect 8312 5250 8340 7686
rect 8404 7478 8432 7890
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8496 7002 8524 8452
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8404 5352 8432 5646
rect 8496 5556 8524 6598
rect 8588 5778 8616 8298
rect 8772 7970 8800 11070
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10674 8984 10950
rect 9048 10810 9076 11562
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9140 11014 9168 11222
rect 9128 11008 9180 11014
rect 9232 10985 9260 11494
rect 9128 10950 9180 10956
rect 9218 10976 9274 10985
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 9140 10742 9168 10950
rect 9218 10911 9274 10920
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8956 10130 8984 10610
rect 9232 10588 9260 10911
rect 9140 10560 9260 10588
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8956 9602 8984 10066
rect 8864 9586 8984 9602
rect 8864 9580 8996 9586
rect 8864 9574 8944 9580
rect 8864 8974 8892 9574
rect 8944 9522 8996 9528
rect 8942 9480 8998 9489
rect 8942 9415 8944 9424
rect 8996 9415 8998 9424
rect 8944 9386 8996 9392
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8772 7942 8892 7970
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6848 8708 7142
rect 8772 7002 8800 7822
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8864 6905 8892 7942
rect 8956 7818 8984 8026
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8942 7304 8998 7313
rect 8942 7239 8944 7248
rect 8996 7239 8998 7248
rect 8944 7210 8996 7216
rect 8944 6928 8996 6934
rect 8850 6896 8906 6905
rect 8680 6820 8800 6848
rect 8944 6870 8996 6876
rect 8850 6831 8906 6840
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8680 5710 8708 6054
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8496 5528 8708 5556
rect 8404 5324 8524 5352
rect 8312 5222 8432 5250
rect 8298 4992 8354 5001
rect 8298 4927 8354 4936
rect 8128 4780 8248 4808
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7654 4176 7710 4185
rect 7654 4111 7710 4120
rect 7668 3670 7696 4111
rect 7760 3738 7788 4558
rect 8128 4026 8156 4780
rect 8312 4758 8340 4927
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4146 8248 4422
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8128 3998 8248 4026
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7668 3210 7696 3470
rect 8128 3466 8156 3606
rect 8220 3534 8248 3998
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8206 3360 8262 3369
rect 8206 3295 8262 3304
rect 7576 3182 7696 3210
rect 7576 2582 7604 3182
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7760 2514 7788 2790
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7484 2400 7696 2428
rect 7668 800 7696 2400
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8036 800 8064 2246
rect 8220 2106 8248 3295
rect 8312 2650 8340 3946
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2378 8432 5222
rect 8496 4729 8524 5324
rect 8574 5264 8630 5273
rect 8574 5199 8630 5208
rect 8482 4720 8538 4729
rect 8482 4655 8538 4664
rect 8496 4622 8524 4655
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8496 2854 8524 4558
rect 8588 3602 8616 5199
rect 8680 4758 8708 5528
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8666 4312 8722 4321
rect 8772 4298 8800 6820
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8864 5370 8892 6122
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8956 4593 8984 6870
rect 8942 4584 8998 4593
rect 8942 4519 8998 4528
rect 8722 4270 8800 4298
rect 8666 4247 8668 4256
rect 8720 4247 8722 4256
rect 8668 4218 8720 4224
rect 8666 4176 8722 4185
rect 8956 4162 8984 4519
rect 8666 4111 8722 4120
rect 8772 4134 8984 4162
rect 8680 3913 8708 4111
rect 8666 3904 8722 3913
rect 8666 3839 8722 3848
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8668 3528 8720 3534
rect 8574 3496 8630 3505
rect 8668 3470 8720 3476
rect 8574 3431 8576 3440
rect 8628 3431 8630 3440
rect 8576 3402 8628 3408
rect 8574 3360 8630 3369
rect 8574 3295 8630 3304
rect 8588 3194 8616 3295
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8680 2990 8708 3470
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8574 2816 8630 2825
rect 8574 2751 8630 2760
rect 8588 2650 8616 2751
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 8680 1834 8708 2518
rect 8668 1828 8720 1834
rect 8668 1770 8720 1776
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8404 800 8432 1362
rect 8772 800 8800 4134
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8864 3777 8892 4014
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8850 3768 8906 3777
rect 8850 3703 8906 3712
rect 8864 2990 8892 3703
rect 8956 3670 8984 3878
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8944 3120 8996 3126
rect 9048 3108 9076 10406
rect 9140 5817 9168 10560
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9232 9353 9260 10134
rect 9218 9344 9274 9353
rect 9218 9279 9274 9288
rect 9232 6372 9260 9279
rect 9324 6934 9352 11750
rect 9416 10577 9444 14214
rect 9508 11286 9536 17206
rect 9600 17202 9628 18006
rect 9678 17912 9734 17921
rect 9678 17847 9734 17856
rect 9692 17814 9720 17847
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 15502 9628 17138
rect 9784 16658 9812 18090
rect 9876 17814 9904 18226
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9876 17134 9904 17750
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9600 15337 9628 15438
rect 9586 15328 9642 15337
rect 9586 15263 9642 15272
rect 9678 12336 9734 12345
rect 9600 12294 9678 12322
rect 9496 11280 9548 11286
rect 9494 11248 9496 11257
rect 9548 11248 9550 11257
rect 9494 11183 9550 11192
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9402 10568 9458 10577
rect 9402 10503 9458 10512
rect 9508 9518 9536 11018
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9402 8120 9458 8129
rect 9402 8055 9458 8064
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9232 6344 9352 6372
rect 9126 5808 9182 5817
rect 9126 5743 9182 5752
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8996 3080 9076 3108
rect 8944 3062 8996 3068
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8956 2854 8984 3062
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8864 2446 8892 2790
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 9140 800 9168 5306
rect 9232 4554 9260 5714
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9232 1426 9260 4490
rect 9324 2038 9352 6344
rect 9416 5370 9444 8055
rect 9508 8022 9536 9318
rect 9600 9178 9628 12294
rect 9678 12271 9734 12280
rect 9784 11830 9812 16458
rect 9968 15994 9996 19246
rect 9876 15966 9996 15994
rect 9876 12782 9904 15966
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15706 9996 15846
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15162 9996 15506
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10060 14906 10088 22000
rect 10140 19984 10192 19990
rect 10140 19926 10192 19932
rect 10152 19310 10180 19926
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16250 10180 16526
rect 10428 16522 10456 22000
rect 10796 19242 10824 22000
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10888 18902 10916 19246
rect 11164 19174 11192 22000
rect 11624 19786 11652 22000
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 10520 17066 10548 18770
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17060 10560 17066
rect 10508 17002 10560 17008
rect 10612 16794 10640 17614
rect 10704 17338 10732 18770
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10152 15570 10180 16050
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10152 15026 10180 15506
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10060 14878 10180 14906
rect 9954 14648 10010 14657
rect 9954 14583 9956 14592
rect 10008 14583 10010 14592
rect 9956 14554 10008 14560
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13938 10088 14214
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9770 11248 9826 11257
rect 9770 11183 9826 11192
rect 9784 11150 9812 11183
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9784 10062 9812 11086
rect 9876 10674 9904 12174
rect 10060 12102 10088 13738
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8430 9720 8910
rect 9770 8664 9826 8673
rect 9770 8599 9826 8608
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9600 7750 9628 8298
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7410 9628 7686
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 5914 9536 7142
rect 9600 6798 9628 7346
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9600 6118 9628 6734
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9692 5953 9720 8230
rect 9784 8022 9812 8599
rect 9876 8566 9904 9522
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9876 7886 9904 8502
rect 9968 8090 9996 9318
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10060 7993 10088 11766
rect 10152 11082 10180 14878
rect 10428 14074 10456 15846
rect 10704 15094 10732 16594
rect 10796 16114 10824 18566
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10980 17542 11008 18090
rect 11072 17882 11100 18158
rect 11164 17882 11192 18362
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10888 16454 10916 17478
rect 10980 17338 11008 17478
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11164 16726 11192 17682
rect 11256 17610 11284 18294
rect 11624 18290 11652 18770
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11624 18086 11652 18226
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11612 18080 11664 18086
rect 11716 18057 11744 18906
rect 11796 18080 11848 18086
rect 11612 18022 11664 18028
rect 11702 18048 11758 18057
rect 11440 17678 11468 18022
rect 11796 18022 11848 18028
rect 11702 17983 11758 17992
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11520 17264 11572 17270
rect 11520 17206 11572 17212
rect 11426 17096 11482 17105
rect 11426 17031 11482 17040
rect 11440 16998 11468 17031
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11334 16824 11390 16833
rect 11334 16759 11336 16768
rect 11388 16759 11390 16768
rect 11336 16730 11388 16736
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11532 16590 11560 17206
rect 11624 16640 11652 17818
rect 11808 17338 11836 18022
rect 11900 17882 11928 19246
rect 11992 19174 12020 22000
rect 12360 19242 12388 22000
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12728 19174 12756 22000
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12164 18896 12216 18902
rect 12164 18838 12216 18844
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11980 17808 12032 17814
rect 11980 17750 12032 17756
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11900 17202 11928 17478
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11716 16776 11744 17070
rect 11796 16788 11848 16794
rect 11716 16748 11796 16776
rect 11796 16730 11848 16736
rect 11796 16652 11848 16658
rect 11624 16612 11744 16640
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11610 16552 11666 16561
rect 11610 16487 11666 16496
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 10966 16144 11022 16153
rect 10784 16108 10836 16114
rect 10966 16079 11022 16088
rect 10784 16050 10836 16056
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10232 13864 10284 13870
rect 10230 13832 10232 13841
rect 10284 13832 10286 13841
rect 10230 13767 10286 13776
rect 10428 13734 10456 13874
rect 10704 13870 10732 15030
rect 10888 14958 10916 15370
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10980 14822 11008 16079
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10796 13734 10824 14758
rect 10980 14498 11008 14758
rect 11072 14618 11100 15846
rect 11164 15366 11192 15914
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11440 14906 11468 14962
rect 11348 14878 11468 14906
rect 11152 14816 11204 14822
rect 11150 14784 11152 14793
rect 11204 14784 11206 14793
rect 11150 14719 11206 14728
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10980 14470 11192 14498
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10980 13938 11008 14214
rect 11072 14074 11100 14350
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10876 13864 10928 13870
rect 10928 13812 11008 13818
rect 10876 13806 11008 13812
rect 10888 13790 11008 13806
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10230 13424 10286 13433
rect 10414 13424 10470 13433
rect 10230 13359 10286 13368
rect 10336 13382 10414 13410
rect 10244 12714 10272 13359
rect 10336 13190 10364 13382
rect 10414 13359 10470 13368
rect 10416 13320 10468 13326
rect 10704 13297 10732 13670
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 10416 13262 10468 13268
rect 10690 13288 10746 13297
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10230 12064 10286 12073
rect 10230 11999 10286 12008
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10138 10432 10194 10441
rect 10138 10367 10194 10376
rect 10046 7984 10102 7993
rect 10046 7919 10102 7928
rect 10152 7886 10180 10367
rect 10244 8265 10272 11999
rect 10336 10130 10364 13126
rect 10428 12986 10456 13262
rect 10600 13252 10652 13258
rect 10520 13212 10600 13240
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10520 12866 10548 13212
rect 10652 13232 10690 13240
rect 10652 13223 10746 13232
rect 10652 13212 10732 13223
rect 10600 13194 10652 13200
rect 10428 12838 10548 12866
rect 10784 12844 10836 12850
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10230 8256 10286 8265
rect 10230 8191 10286 8200
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7585 9812 7754
rect 9770 7576 9826 7585
rect 9770 7511 9826 7520
rect 9956 7472 10008 7478
rect 9876 7420 9956 7426
rect 9876 7414 10008 7420
rect 9876 7398 9996 7414
rect 10232 7404 10284 7410
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6866 9812 7142
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9678 5944 9734 5953
rect 9496 5908 9548 5914
rect 9678 5879 9734 5888
rect 9496 5850 9548 5856
rect 9508 5642 9536 5850
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4826 9628 4966
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9692 4758 9720 5510
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9416 3942 9444 4558
rect 9772 4140 9824 4146
rect 9692 4100 9772 4128
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9402 3088 9458 3097
rect 9402 3023 9458 3032
rect 9416 2310 9444 3023
rect 9508 2582 9536 3946
rect 9586 3768 9642 3777
rect 9586 3703 9642 3712
rect 9600 3602 9628 3703
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9312 2032 9364 2038
rect 9312 1974 9364 1980
rect 9600 1442 9628 3130
rect 9692 2514 9720 4100
rect 9772 4082 9824 4088
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9784 3602 9812 3674
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9220 1420 9272 1426
rect 9220 1362 9272 1368
rect 9508 1414 9628 1442
rect 9508 800 9536 1414
rect 9876 800 9904 7398
rect 10232 7346 10284 7352
rect 10140 6928 10192 6934
rect 10138 6896 10140 6905
rect 10192 6896 10194 6905
rect 9956 6860 10008 6866
rect 10138 6831 10194 6840
rect 9956 6802 10008 6808
rect 9968 6662 9996 6802
rect 10244 6798 10272 7346
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 10244 6186 10272 6734
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10140 6112 10192 6118
rect 9968 6060 10140 6066
rect 9968 6054 10192 6060
rect 10230 6080 10286 6089
rect 9968 6038 10180 6054
rect 9968 5710 9996 6038
rect 10230 6015 10286 6024
rect 10244 5914 10272 6015
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10060 5234 10088 5714
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10244 5370 10272 5646
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10140 5228 10192 5234
rect 10244 5216 10272 5306
rect 10192 5188 10272 5216
rect 10140 5170 10192 5176
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 4729 9996 5102
rect 9954 4720 10010 4729
rect 9954 4655 10010 4664
rect 10152 4554 10180 5170
rect 10336 5114 10364 9590
rect 10428 7478 10456 12838
rect 10784 12786 10836 12792
rect 10600 12776 10652 12782
rect 10598 12744 10600 12753
rect 10652 12744 10654 12753
rect 10598 12679 10654 12688
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 10044 10548 12038
rect 10612 10198 10640 12679
rect 10796 12306 10824 12786
rect 10888 12345 10916 13398
rect 10980 12714 11008 13790
rect 11072 13705 11100 14010
rect 11164 13802 11192 14470
rect 11348 14414 11376 14878
rect 11624 14804 11652 16487
rect 11716 14929 11744 16612
rect 11796 16594 11848 16600
rect 11808 15473 11836 16594
rect 11992 16250 12020 17750
rect 12176 17746 12204 18838
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12268 17882 12296 18090
rect 12346 17912 12402 17921
rect 12256 17876 12308 17882
rect 12346 17847 12402 17856
rect 12256 17818 12308 17824
rect 12360 17814 12388 17847
rect 12348 17808 12400 17814
rect 12254 17776 12310 17785
rect 12164 17740 12216 17746
rect 12348 17750 12400 17756
rect 12254 17711 12310 17720
rect 12164 17682 12216 17688
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11992 15638 12020 16186
rect 12084 15706 12112 17614
rect 12176 16130 12204 17682
rect 12268 17678 12296 17711
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12268 16561 12296 17614
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12530 17232 12586 17241
rect 12530 17167 12586 17176
rect 12544 17066 12572 17167
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12254 16552 12310 16561
rect 12254 16487 12310 16496
rect 12176 16102 12388 16130
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12072 15496 12124 15502
rect 11794 15464 11850 15473
rect 12072 15438 12124 15444
rect 11794 15399 11850 15408
rect 12084 15065 12112 15438
rect 12070 15056 12126 15065
rect 12070 14991 12126 15000
rect 11702 14920 11758 14929
rect 11702 14855 11758 14864
rect 11888 14816 11940 14822
rect 11624 14776 11836 14804
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11242 13968 11298 13977
rect 11624 13938 11652 14418
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11242 13903 11298 13912
rect 11612 13932 11664 13938
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11058 13696 11114 13705
rect 11256 13682 11284 13903
rect 11612 13874 11664 13880
rect 11716 13870 11744 14350
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11058 13631 11114 13640
rect 11164 13654 11284 13682
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11072 12986 11100 13330
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11164 12866 11192 13654
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11072 12838 11192 12866
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10874 12336 10930 12345
rect 10784 12300 10836 12306
rect 10874 12271 10930 12280
rect 10784 12242 10836 12248
rect 10690 11792 10746 11801
rect 10796 11762 10824 12242
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10690 11727 10746 11736
rect 10784 11756 10836 11762
rect 10704 11694 10732 11727
rect 10784 11698 10836 11704
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 10266 10732 11494
rect 10796 10810 10824 11698
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10888 10606 10916 12038
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10980 10130 11008 12650
rect 11072 12646 11100 12838
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11072 10690 11100 12582
rect 11164 12102 11192 12582
rect 11532 12238 11560 12854
rect 11624 12442 11652 13262
rect 11716 12442 11744 13670
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11150 11792 11206 11801
rect 11624 11762 11652 12378
rect 11704 12300 11756 12306
rect 11808 12288 11836 14776
rect 11888 14758 11940 14764
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11900 14006 11928 14758
rect 11992 14657 12020 14758
rect 11978 14648 12034 14657
rect 11978 14583 12034 14592
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11756 12260 11836 12288
rect 11704 12242 11756 12248
rect 11150 11727 11206 11736
rect 11612 11756 11664 11762
rect 11164 10810 11192 11727
rect 11612 11698 11664 11704
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11624 11218 11652 11290
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11072 10662 11192 10690
rect 11164 10606 11192 10662
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 11072 10062 11100 10474
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10266 11192 10406
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11716 10198 11744 12242
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11808 10538 11836 11834
rect 11992 11257 12020 14282
rect 12084 13977 12112 14991
rect 12070 13968 12126 13977
rect 12070 13903 12126 13912
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 10784 10056 10836 10062
rect 10520 10016 10640 10044
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10520 8809 10548 9386
rect 10612 8922 10640 10016
rect 10784 9998 10836 10004
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10612 8894 10732 8922
rect 10506 8800 10562 8809
rect 10506 8735 10562 8744
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10520 8362 10548 8570
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10598 8256 10654 8265
rect 10598 8191 10654 8200
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10520 7342 10548 7958
rect 10508 7336 10560 7342
rect 10506 7304 10508 7313
rect 10560 7304 10562 7313
rect 10612 7274 10640 8191
rect 10704 7954 10732 8894
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7585 10732 7686
rect 10690 7576 10746 7585
rect 10690 7511 10746 7520
rect 10506 7239 10562 7248
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10796 7154 10824 9998
rect 10968 9648 11020 9654
rect 10966 9616 10968 9625
rect 11020 9616 11022 9625
rect 10966 9551 11022 9560
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 9042 10916 9318
rect 11072 9178 11100 9998
rect 11164 9704 11192 10066
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11164 9676 11560 9704
rect 11336 9580 11388 9586
rect 11164 9540 11336 9568
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10244 5086 10364 5114
rect 10428 7126 10824 7154
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9968 1426 9996 4150
rect 10060 2650 10088 4422
rect 10152 4078 10180 4490
rect 10244 4214 10272 5086
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10336 4826 10364 4966
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10140 4072 10192 4078
rect 10428 4026 10456 7126
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10520 6662 10548 6870
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 6254 10548 6598
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10520 4826 10548 5510
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10612 4622 10640 6122
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10704 5574 10732 5850
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10690 4856 10746 4865
rect 10690 4791 10746 4800
rect 10704 4690 10732 4791
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10140 4014 10192 4020
rect 10244 3998 10456 4026
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3058 10180 3878
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9956 1420 10008 1426
rect 9956 1362 10008 1368
rect 10244 800 10272 3998
rect 10612 3913 10640 4558
rect 10692 3936 10744 3942
rect 10598 3904 10654 3913
rect 10692 3878 10744 3884
rect 10598 3839 10654 3848
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10336 3194 10364 3538
rect 10598 3224 10654 3233
rect 10324 3188 10376 3194
rect 10598 3159 10654 3168
rect 10324 3130 10376 3136
rect 10336 2446 10364 3130
rect 10416 2848 10468 2854
rect 10612 2825 10640 3159
rect 10704 2922 10732 3878
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10416 2790 10468 2796
rect 10598 2816 10654 2825
rect 10428 2650 10456 2790
rect 10796 2802 10824 5782
rect 10888 5710 10916 8774
rect 10980 7954 11008 9046
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8673 11100 8910
rect 11058 8664 11114 8673
rect 11058 8599 11060 8608
rect 11112 8599 11114 8608
rect 11060 8570 11112 8576
rect 11072 8539 11100 8570
rect 11164 8498 11192 9540
rect 11336 9522 11388 9528
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11440 9450 11468 9522
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11532 9194 11560 9676
rect 11624 9466 11652 10066
rect 11808 9926 11836 10474
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11900 9518 11928 10474
rect 11992 10266 12020 10950
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9586 12020 9862
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 9512 11940 9518
rect 11624 9438 11836 9466
rect 11888 9454 11940 9460
rect 11702 9208 11758 9217
rect 11532 9166 11652 9194
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8514 11652 9166
rect 11702 9143 11704 9152
rect 11756 9143 11758 9152
rect 11704 9114 11756 9120
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 8634 11744 8910
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11152 8492 11204 8498
rect 11624 8486 11744 8514
rect 11152 8434 11204 8440
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 8090 11652 8230
rect 11612 8084 11664 8090
rect 11072 8044 11284 8072
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 11072 7834 11100 8044
rect 10980 7806 11100 7834
rect 11256 7818 11284 8044
rect 11612 8026 11664 8032
rect 11244 7812 11296 7818
rect 10980 6934 11008 7806
rect 11244 7754 11296 7760
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7002 11100 7686
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11164 7002 11192 7210
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10888 4146 10916 5510
rect 10980 5166 11008 6734
rect 11072 6497 11100 6802
rect 11058 6488 11114 6497
rect 11058 6423 11114 6432
rect 11164 6322 11192 6938
rect 11348 6798 11376 7210
rect 11532 6934 11560 7210
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11716 6361 11744 8486
rect 11702 6352 11758 6361
rect 11152 6316 11204 6322
rect 11702 6287 11758 6296
rect 11152 6258 11204 6264
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5953 11560 6054
rect 11242 5944 11298 5953
rect 11242 5879 11298 5888
rect 11518 5944 11574 5953
rect 11518 5879 11574 5888
rect 11256 5710 11284 5879
rect 11716 5846 11744 6122
rect 11808 5914 11836 9438
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11886 9208 11942 9217
rect 11886 9143 11942 9152
rect 11900 7154 11928 9143
rect 11992 8673 12020 9386
rect 11978 8664 12034 8673
rect 11978 8599 12034 8608
rect 12084 7478 12112 13806
rect 12176 13802 12204 15506
rect 12268 14482 12296 15982
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12268 13870 12296 14418
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12162 13696 12218 13705
rect 12162 13631 12218 13640
rect 12176 12764 12204 13631
rect 12268 12918 12296 13806
rect 12256 12912 12308 12918
rect 12360 12889 12388 16102
rect 12452 15570 12480 16934
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12544 15994 12572 16594
rect 12636 16114 12664 17478
rect 12820 17082 12848 19178
rect 13004 18714 13032 19246
rect 13096 19224 13124 22000
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13280 19378 13308 19858
rect 13464 19394 13492 22000
rect 13832 20058 13860 22000
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13268 19372 13320 19378
rect 13464 19366 13584 19394
rect 13268 19314 13320 19320
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13176 19236 13228 19242
rect 13096 19196 13176 19224
rect 13176 19178 13228 19184
rect 13464 18970 13492 19246
rect 13556 19242 13584 19366
rect 13832 19366 14044 19394
rect 13832 19310 13860 19366
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13924 18902 13952 19246
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13004 18686 13216 18714
rect 13188 18426 13216 18686
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 13004 18154 13032 18294
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 12898 18048 12954 18057
rect 12898 17983 12954 17992
rect 12912 17202 12940 17983
rect 13464 17678 13492 18566
rect 13740 17746 13768 18566
rect 13832 18290 13860 18770
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13452 17672 13504 17678
rect 13280 17632 13452 17660
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 13004 17105 13032 17274
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12728 17054 12848 17082
rect 12990 17096 13046 17105
rect 12728 16833 12756 17054
rect 12990 17031 13046 17040
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12714 16824 12770 16833
rect 12912 16794 12940 16934
rect 12714 16759 12770 16768
rect 12900 16788 12952 16794
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12544 15966 12664 15994
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12986 12480 13126
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12256 12854 12308 12860
rect 12346 12880 12402 12889
rect 12346 12815 12402 12824
rect 12176 12736 12296 12764
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12176 11665 12204 12310
rect 12162 11656 12218 11665
rect 12162 11591 12218 11600
rect 12162 11248 12218 11257
rect 12162 11183 12218 11192
rect 12176 10044 12204 11183
rect 12268 10996 12296 12736
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11694 12388 12038
rect 12348 11688 12400 11694
rect 12400 11648 12480 11676
rect 12348 11630 12400 11636
rect 12452 11150 12480 11648
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12268 10968 12388 10996
rect 12176 10016 12296 10044
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12176 9110 12204 9522
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12162 8800 12218 8809
rect 12162 8735 12218 8744
rect 12176 8566 12204 8735
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11900 7126 12020 7154
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11072 5098 11100 5646
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11072 4622 11100 5034
rect 11532 5001 11560 5034
rect 11518 4992 11574 5001
rect 11518 4927 11574 4936
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 11072 3720 11100 4422
rect 11164 4214 11192 4626
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11624 4146 11652 4558
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11716 4078 11744 5510
rect 11900 5352 11928 6967
rect 11992 6225 12020 7126
rect 11978 6216 12034 6225
rect 11978 6151 12034 6160
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5794 12020 6054
rect 12084 5914 12112 7414
rect 12176 7206 12204 8502
rect 12268 7954 12296 10016
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12360 7750 12388 10968
rect 12438 10976 12494 10985
rect 12438 10911 12494 10920
rect 12452 10606 12480 10911
rect 12544 10792 12572 15846
rect 12636 14929 12664 15966
rect 12622 14920 12678 14929
rect 12622 14855 12678 14864
rect 12636 12646 12664 14855
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12728 11393 12756 16759
rect 12900 16730 12952 16736
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12820 15609 12848 15642
rect 12900 15632 12952 15638
rect 12806 15600 12862 15609
rect 12900 15574 12952 15580
rect 12806 15535 12862 15544
rect 12912 15450 12940 15574
rect 12820 15422 12940 15450
rect 12820 13977 12848 15422
rect 12806 13968 12862 13977
rect 12806 13903 12862 13912
rect 12820 13462 12848 13903
rect 12898 13832 12954 13841
rect 13096 13802 13124 17138
rect 13280 17134 13308 17632
rect 13452 17614 13504 17620
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13280 16250 13308 16526
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13372 15994 13400 16118
rect 13280 15966 13400 15994
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14074 13216 14758
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12898 13767 12954 13776
rect 13084 13796 13136 13802
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12808 13184 12860 13190
rect 12912 13161 12940 13767
rect 13084 13738 13136 13744
rect 13096 13326 13124 13738
rect 13280 13530 13308 15966
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15706 13400 15846
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13556 15178 13584 16730
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 15706 13676 16390
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13648 15337 13676 15438
rect 13740 15434 13768 17682
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13832 16250 13860 16594
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 14016 16153 14044 19366
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14108 16182 14136 19178
rect 14200 19174 14228 22000
rect 14660 20346 14688 22000
rect 14568 20318 14688 20346
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14292 16998 14320 18770
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14292 16454 14320 16662
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14096 16176 14148 16182
rect 14002 16144 14058 16153
rect 14096 16118 14148 16124
rect 14002 16079 14058 16088
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14016 15638 14044 15982
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13634 15328 13690 15337
rect 13634 15263 13690 15272
rect 13556 15150 13768 15178
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13648 14550 13676 14894
rect 13740 14822 13768 15150
rect 13832 15116 14044 15144
rect 13832 14822 13860 15116
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13924 14618 13952 14962
rect 14016 14618 14044 15116
rect 14200 15026 14228 16050
rect 14384 15994 14412 19246
rect 14568 19174 14596 20318
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15028 19174 15056 22000
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15212 19378 15240 20198
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 15120 18902 15148 19246
rect 15396 19174 15424 22000
rect 15764 20058 15792 22000
rect 16132 20058 16160 22000
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15108 18896 15160 18902
rect 15108 18838 15160 18844
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14554 17640 14610 17649
rect 14554 17575 14556 17584
rect 14608 17575 14610 17584
rect 14556 17546 14608 17552
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14476 17066 14504 17478
rect 14568 17066 14872 17082
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14568 17060 14884 17066
rect 14568 17054 14832 17060
rect 14476 16114 14504 17002
rect 14568 16998 14596 17054
rect 14832 17002 14884 17008
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14568 16590 14596 16934
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14660 16250 14688 16594
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14280 15972 14332 15978
rect 14384 15966 14596 15994
rect 14280 15914 14332 15920
rect 14292 15042 14320 15914
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15706 14412 15846
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14568 15570 14596 15966
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14188 15020 14240 15026
rect 14292 15014 14412 15042
rect 14188 14962 14240 14968
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13832 13870 13860 14418
rect 13924 14006 13952 14554
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13464 13530 13492 13670
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13280 13326 13308 13466
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13372 13172 13400 13330
rect 12808 13126 12860 13132
rect 12898 13152 12954 13161
rect 12714 11384 12770 11393
rect 12714 11319 12770 11328
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12544 10764 12664 10792
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12636 10418 12664 10764
rect 12728 10742 12756 11154
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12820 10606 12848 13126
rect 12898 13087 12954 13096
rect 13188 13144 13400 13172
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11694 13032 12038
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 10674 12940 11494
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12636 10390 12848 10418
rect 12820 10130 12848 10390
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12544 9761 12572 9930
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12452 8634 12480 9454
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 7886 12480 8570
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12348 7744 12400 7750
rect 12346 7712 12348 7721
rect 12400 7712 12402 7721
rect 12346 7647 12402 7656
rect 12360 7621 12388 7647
rect 12452 7546 12480 7822
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12360 7313 12388 7482
rect 12452 7342 12480 7482
rect 12440 7336 12492 7342
rect 12346 7304 12402 7313
rect 12440 7278 12492 7284
rect 12636 7256 12664 9998
rect 12820 9722 12848 10066
rect 13096 10062 13124 10542
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 13082 9616 13138 9625
rect 13082 9551 13138 9560
rect 13096 9330 13124 9551
rect 12912 9302 13124 9330
rect 12912 9058 12940 9302
rect 12820 9030 12940 9058
rect 12820 8974 12848 9030
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12808 8832 12860 8838
rect 12806 8800 12808 8809
rect 12860 8800 12862 8809
rect 12806 8735 12862 8744
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12346 7239 12402 7248
rect 12544 7228 12664 7256
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12348 7200 12400 7206
rect 12544 7154 12572 7228
rect 12348 7142 12400 7148
rect 12360 7018 12388 7142
rect 12268 6990 12388 7018
rect 12452 7126 12572 7154
rect 12268 6322 12296 6990
rect 12452 6662 12480 7126
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12622 6896 12678 6905
rect 12622 6831 12678 6840
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12440 6452 12492 6458
rect 12544 6440 12572 6598
rect 12492 6412 12572 6440
rect 12440 6394 12492 6400
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12254 6080 12310 6089
rect 12254 6015 12310 6024
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 12268 5846 12296 6015
rect 12256 5840 12308 5846
rect 11992 5766 12204 5794
rect 12256 5782 12308 5788
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5574 12020 5646
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12070 5536 12126 5545
rect 12070 5471 12126 5480
rect 12084 5352 12112 5471
rect 11900 5324 12112 5352
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11808 4214 11836 4490
rect 11900 4282 11928 5170
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 10980 3692 11100 3720
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10888 2990 10916 3334
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10980 2922 11008 3692
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10796 2774 11008 2802
rect 10598 2751 10654 2760
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10600 1420 10652 1426
rect 10600 1362 10652 1368
rect 10612 800 10640 1362
rect 10980 800 11008 2774
rect 11072 2582 11100 3538
rect 11164 2854 11192 3878
rect 11702 3768 11758 3777
rect 11808 3738 11836 3878
rect 11702 3703 11758 3712
rect 11796 3732 11848 3738
rect 11716 3670 11744 3703
rect 11796 3674 11848 3680
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11624 1170 11652 2246
rect 11348 1142 11652 1170
rect 11348 800 11376 1142
rect 11716 898 11744 3334
rect 11808 2990 11836 3334
rect 11992 3097 12020 4626
rect 12084 3738 12112 5324
rect 12176 4282 12204 5766
rect 12346 4992 12402 5001
rect 12346 4927 12402 4936
rect 12360 4826 12388 4927
rect 12636 4826 12664 6831
rect 12728 6254 12756 6938
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12820 5302 12848 8230
rect 12912 7834 12940 8910
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 8498 13032 8774
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8022 13032 8434
rect 13096 8022 13124 9302
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 12912 7806 13124 7834
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6186 12940 7142
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 13004 6905 13032 6938
rect 12990 6896 13046 6905
rect 12990 6831 13046 6840
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 13096 6066 13124 7806
rect 13004 6038 13124 6066
rect 13004 5370 13032 6038
rect 13082 5400 13138 5409
rect 12992 5364 13044 5370
rect 13082 5335 13138 5344
rect 12992 5306 13044 5312
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12176 3534 12204 4014
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12544 3738 12572 3878
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12728 3670 12756 4422
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 11978 3088 12034 3097
rect 12452 3058 12480 3402
rect 11978 3023 12034 3032
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 11796 2984 11848 2990
rect 13004 2961 13032 5306
rect 13096 4690 13124 5335
rect 13188 5216 13216 13144
rect 13464 12889 13492 13330
rect 13740 13326 13768 13738
rect 13832 13734 13860 13806
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13450 12880 13506 12889
rect 13450 12815 13506 12824
rect 13648 12458 13676 13262
rect 13740 12850 13768 13262
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13832 12730 13860 13330
rect 14016 13190 14044 14418
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13556 12430 13676 12458
rect 13740 12702 13860 12730
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13280 10674 13308 11630
rect 13372 11354 13400 12378
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13280 9450 13308 9998
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13280 8498 13308 9386
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13266 7168 13322 7177
rect 13266 7103 13322 7112
rect 13280 6866 13308 7103
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13268 5228 13320 5234
rect 13188 5188 13268 5216
rect 13268 5170 13320 5176
rect 13280 5030 13308 5170
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13084 4684 13136 4690
rect 13136 4644 13216 4672
rect 13084 4626 13136 4632
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13096 3194 13124 3470
rect 13188 3466 13216 4644
rect 13280 3641 13308 4966
rect 13266 3632 13322 3641
rect 13266 3567 13322 3576
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 11796 2926 11848 2932
rect 12990 2952 13046 2961
rect 11888 2916 11940 2922
rect 13280 2922 13308 3470
rect 12990 2887 13046 2896
rect 13268 2916 13320 2922
rect 11888 2858 11940 2864
rect 13268 2858 13320 2864
rect 11900 2514 11928 2858
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12912 2446 12940 2586
rect 13096 2514 13124 2790
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 13372 2446 13400 10746
rect 13452 9036 13504 9042
rect 13556 9024 13584 12430
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10674 13676 10950
rect 13740 10713 13768 12702
rect 14016 12442 14044 13126
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 11286 13860 11494
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13726 10704 13782 10713
rect 13636 10668 13688 10674
rect 13726 10639 13782 10648
rect 13636 10610 13688 10616
rect 13648 10062 13676 10610
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13636 10056 13688 10062
rect 13740 10033 13768 10066
rect 13832 10062 13860 11222
rect 13924 10470 13952 12242
rect 14108 12186 14136 13466
rect 14200 13410 14228 14554
rect 14292 13530 14320 14826
rect 14384 13569 14412 15014
rect 14370 13560 14426 13569
rect 14280 13524 14332 13530
rect 14370 13495 14426 13504
rect 14280 13466 14332 13472
rect 14200 13382 14320 13410
rect 14292 12889 14320 13382
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14384 12918 14412 13262
rect 14372 12912 14424 12918
rect 14278 12880 14334 12889
rect 14372 12854 14424 12860
rect 14278 12815 14334 12824
rect 14016 12158 14136 12186
rect 13912 10464 13964 10470
rect 14016 10441 14044 12158
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11098 14136 12038
rect 14108 11070 14228 11098
rect 14094 10704 14150 10713
rect 14094 10639 14150 10648
rect 13912 10406 13964 10412
rect 14002 10432 14058 10441
rect 13820 10056 13872 10062
rect 13636 9998 13688 10004
rect 13726 10024 13782 10033
rect 13648 9625 13676 9998
rect 13820 9998 13872 10004
rect 13726 9959 13782 9968
rect 13634 9616 13690 9625
rect 13634 9551 13690 9560
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 9110 13860 9318
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13556 8996 13676 9024
rect 13452 8978 13504 8984
rect 13464 8650 13492 8978
rect 13464 8622 13584 8650
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13464 7342 13492 8502
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 4078 13492 7142
rect 13556 5114 13584 8622
rect 13648 7886 13676 8996
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13740 8430 13768 8774
rect 13832 8673 13860 8774
rect 13818 8664 13874 8673
rect 13818 8599 13874 8608
rect 13924 8430 13952 10406
rect 14002 10367 14058 10376
rect 14108 10266 14136 10639
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14094 10024 14150 10033
rect 14016 9586 14044 9998
rect 14094 9959 14096 9968
rect 14148 9959 14150 9968
rect 14096 9930 14148 9936
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14016 8974 14044 9522
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14094 8664 14150 8673
rect 14094 8599 14150 8608
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7410 13676 7686
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13648 6934 13676 7346
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13740 5778 13768 7958
rect 13832 7342 13860 8230
rect 14108 8090 14136 8599
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13820 7336 13872 7342
rect 13912 7336 13964 7342
rect 13820 7278 13872 7284
rect 13910 7304 13912 7313
rect 13964 7304 13966 7313
rect 13910 7239 13966 7248
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 6089 13860 6666
rect 13924 6390 13952 7142
rect 14016 6390 14044 7890
rect 14108 7041 14136 8026
rect 14094 7032 14150 7041
rect 14094 6967 14150 6976
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14200 6882 14228 11070
rect 14292 10606 14320 12815
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 11354 14412 12242
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14384 10130 14412 11086
rect 14476 10713 14504 15438
rect 15028 15094 15056 18770
rect 15856 17338 15884 19858
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15948 18630 15976 19246
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 15212 16658 15240 16934
rect 16132 16726 16160 16934
rect 16120 16720 16172 16726
rect 15290 16688 15346 16697
rect 15200 16652 15252 16658
rect 16120 16662 16172 16668
rect 15290 16623 15346 16632
rect 15200 16594 15252 16600
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15120 15706 15148 15846
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15212 15502 15240 16594
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15212 15026 15240 15438
rect 15304 15065 15332 16623
rect 15290 15056 15346 15065
rect 15200 15020 15252 15026
rect 15290 14991 15346 15000
rect 15200 14962 15252 14968
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 12102 14596 14758
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 15212 13938 15240 14962
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15106 13832 15162 13841
rect 15106 13767 15162 13776
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14660 13002 14688 13330
rect 15028 13326 15056 13670
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14660 12986 14780 13002
rect 14660 12980 14792 12986
rect 14660 12974 14740 12980
rect 14740 12922 14792 12928
rect 15120 12918 15148 13767
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15120 12442 15148 12582
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15212 12322 15240 13874
rect 15304 12986 15332 14991
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15948 14618 15976 14758
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15580 13258 15608 14418
rect 16040 14414 16068 14758
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15660 13864 15712 13870
rect 16028 13864 16080 13870
rect 15712 13824 15884 13852
rect 15660 13806 15712 13812
rect 15658 13424 15714 13433
rect 15856 13394 15884 13824
rect 16026 13832 16028 13841
rect 16080 13832 16082 13841
rect 16026 13767 16082 13776
rect 15658 13359 15660 13368
rect 15712 13359 15714 13368
rect 15844 13388 15896 13394
rect 15660 13330 15712 13336
rect 15844 13330 15896 13336
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15120 12294 15240 12322
rect 15580 12306 15608 12786
rect 15384 12300 15436 12306
rect 15120 12238 15148 12294
rect 15384 12242 15436 12248
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 15120 11694 15148 12174
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15212 11354 15240 12106
rect 15396 11898 15424 12242
rect 15672 12186 15700 13330
rect 16132 12986 16160 14418
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16224 13530 16252 14350
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16316 13138 16344 19790
rect 16500 19394 16528 22000
rect 16500 19366 16620 19394
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16500 18902 16528 19246
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16592 16794 16620 19366
rect 16868 19174 16896 22000
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16684 16522 16712 17070
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15706 16436 15846
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16500 15570 16528 16050
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16408 14074 16436 14894
rect 16500 14822 16528 15506
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16408 13258 16436 14010
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16316 13110 16436 13138
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 15488 12158 15700 12186
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15304 11218 15332 11562
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14462 10704 14518 10713
rect 14462 10639 14518 10648
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14476 9976 14504 10639
rect 14292 9948 14504 9976
rect 14292 8294 14320 9948
rect 14462 9888 14518 9897
rect 14462 9823 14518 9832
rect 14370 9616 14426 9625
rect 14370 9551 14426 9560
rect 14384 9353 14412 9551
rect 14476 9450 14504 9823
rect 14464 9444 14516 9450
rect 14568 9432 14596 11154
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15028 10810 15056 11086
rect 15304 11082 15332 11154
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15106 10568 15162 10577
rect 15106 10503 15108 10512
rect 15160 10503 15162 10512
rect 15108 10474 15160 10480
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14738 10160 14794 10169
rect 14738 10095 14740 10104
rect 14792 10095 14794 10104
rect 14740 10066 14792 10072
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14936 9489 14964 9522
rect 14464 9386 14516 9392
rect 14559 9404 14596 9432
rect 14922 9480 14978 9489
rect 14922 9415 14978 9424
rect 14370 9344 14426 9353
rect 14559 9330 14587 9404
rect 15028 9364 15056 10406
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 9518 15148 9862
rect 15212 9722 15240 9930
rect 15290 9752 15346 9761
rect 15200 9716 15252 9722
rect 15290 9687 15346 9696
rect 15200 9658 15252 9664
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15200 9376 15252 9382
rect 15028 9336 15148 9364
rect 14559 9302 14596 9330
rect 14370 9279 14426 9288
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14384 8634 14412 9046
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14384 8090 14412 8366
rect 14476 8362 14504 8774
rect 14568 8362 14596 9302
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15028 9042 15056 9114
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14740 8560 14792 8566
rect 14844 8548 14872 8910
rect 15120 8673 15148 9336
rect 15200 9318 15252 9324
rect 15212 9178 15240 9318
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15198 9072 15254 9081
rect 15198 9007 15200 9016
rect 15252 9007 15254 9016
rect 15200 8978 15252 8984
rect 15106 8664 15162 8673
rect 15106 8599 15162 8608
rect 14792 8520 14872 8548
rect 14740 8502 14792 8508
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 15016 8288 15068 8294
rect 14462 8256 14518 8265
rect 15016 8230 15068 8236
rect 14462 8191 14518 8200
rect 14476 8090 14504 8191
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14292 7290 14320 7482
rect 14556 7404 14608 7410
rect 15028 7392 15056 8230
rect 15120 7954 15148 8434
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15028 7364 15148 7392
rect 14556 7346 14608 7352
rect 14292 7262 14504 7290
rect 14292 6984 14320 7262
rect 14476 7206 14504 7262
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14462 7032 14518 7041
rect 14292 6956 14412 6984
rect 14462 6967 14518 6976
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13912 6112 13964 6118
rect 13818 6080 13874 6089
rect 13912 6054 13964 6060
rect 13818 6015 13874 6024
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13924 5409 13952 6054
rect 13910 5400 13966 5409
rect 14108 5370 14136 6870
rect 14200 6854 14320 6882
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14200 5914 14228 6734
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 13910 5335 13966 5344
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13818 5128 13874 5137
rect 13556 5086 13676 5114
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4146 13584 4966
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13556 2990 13584 3606
rect 13648 3058 13676 5086
rect 13818 5063 13874 5072
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13740 4214 13768 4422
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13740 3670 13768 4150
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13464 2446 13492 2518
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 13636 2372 13688 2378
rect 13636 2314 13688 2320
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 11716 870 11836 898
rect 11808 800 11836 870
rect 12176 800 12204 2246
rect 12544 800 12572 2314
rect 13268 1488 13320 1494
rect 13268 1430 13320 1436
rect 12900 1420 12952 1426
rect 12900 1362 12952 1368
rect 12912 800 12940 1362
rect 13280 800 13308 1430
rect 13648 800 13676 2314
rect 13740 1494 13768 3062
rect 13832 2514 13860 5063
rect 13924 5030 13952 5170
rect 14016 5030 14044 5306
rect 14200 5234 14228 5646
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14094 4992 14150 5001
rect 14094 4927 14150 4936
rect 14108 4690 14136 4927
rect 14292 4865 14320 6854
rect 14384 6118 14412 6956
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14278 4856 14334 4865
rect 14384 4826 14412 5510
rect 14278 4791 14334 4800
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13924 4214 13952 4626
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 13912 4072 13964 4078
rect 13910 4040 13912 4049
rect 13964 4040 13966 4049
rect 13910 3975 13966 3984
rect 14278 3496 14334 3505
rect 14278 3431 14334 3440
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13728 1488 13780 1494
rect 13728 1430 13780 1436
rect 14016 800 14044 2586
rect 14292 2514 14320 3431
rect 14476 2514 14504 6967
rect 14568 6662 14596 7346
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14660 6474 14688 6870
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14568 6446 14688 6474
rect 14568 3738 14596 6446
rect 14936 6100 14964 6734
rect 15028 6730 15056 7210
rect 15120 6934 15148 7364
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15016 6112 15068 6118
rect 14936 6072 15016 6100
rect 15016 6054 15068 6060
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15028 5710 15056 6054
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14830 4448 14886 4457
rect 14830 4383 14886 4392
rect 14844 4146 14872 4383
rect 15028 4146 15056 5646
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 4865 15148 5578
rect 15212 5370 15240 5714
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15106 4856 15162 4865
rect 15106 4791 15162 4800
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15304 3777 15332 9687
rect 15396 8294 15424 10406
rect 15488 10010 15516 12158
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15672 10810 15700 11154
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 10130 15608 10610
rect 15764 10266 15792 12922
rect 15936 12912 15988 12918
rect 15934 12880 15936 12889
rect 15988 12880 15990 12889
rect 15934 12815 15990 12824
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15488 9982 15608 10010
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15488 9178 15516 9522
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15474 9072 15530 9081
rect 15474 9007 15530 9016
rect 15488 8906 15516 9007
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 8090 15424 8230
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15396 6458 15424 7210
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15396 5817 15424 5850
rect 15382 5808 15438 5817
rect 15382 5743 15438 5752
rect 15290 3768 15346 3777
rect 14556 3732 14608 3738
rect 15290 3703 15346 3712
rect 14556 3674 14608 3680
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14108 1426 14136 2246
rect 14096 1420 14148 1426
rect 14096 1362 14148 1368
rect 14384 800 14412 2246
rect 14752 800 14780 2518
rect 15488 2514 15516 7482
rect 15580 5386 15608 9982
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15672 8906 15700 9862
rect 15842 9480 15898 9489
rect 15842 9415 15898 9424
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15764 8945 15792 9114
rect 15750 8936 15806 8945
rect 15660 8900 15712 8906
rect 15750 8871 15806 8880
rect 15660 8842 15712 8848
rect 15672 7750 15700 8842
rect 15856 8566 15884 9415
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 6322 15700 7686
rect 15764 7206 15792 8230
rect 15842 7440 15898 7449
rect 15842 7375 15898 7384
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15856 7002 15884 7375
rect 15948 7274 15976 12718
rect 16040 11898 16068 12786
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16040 11694 16068 11834
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16132 11354 16160 12582
rect 16408 12442 16436 13110
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 16040 7041 16068 10134
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16026 7032 16082 7041
rect 15844 6996 15896 7002
rect 16026 6967 16082 6976
rect 15844 6938 15896 6944
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15672 5642 15700 6258
rect 15764 6225 15792 6734
rect 15750 6216 15806 6225
rect 15750 6151 15806 6160
rect 15856 5778 15884 6938
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15948 5710 15976 6054
rect 16040 5778 16068 6734
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15580 5358 15792 5386
rect 15660 5160 15712 5166
rect 15658 5128 15660 5137
rect 15712 5128 15714 5137
rect 15658 5063 15714 5072
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4185 15608 4966
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4593 15700 4626
rect 15658 4584 15714 4593
rect 15658 4519 15714 4528
rect 15566 4176 15622 4185
rect 15566 4111 15622 4120
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15580 3058 15608 3878
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 15120 800 15148 2314
rect 15672 1442 15700 2790
rect 15764 2514 15792 5358
rect 15948 5234 15976 5646
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16040 4622 16068 5714
rect 16132 5302 16160 9386
rect 16120 5296 16172 5302
rect 16118 5264 16120 5273
rect 16172 5264 16174 5273
rect 16118 5199 16174 5208
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15842 4176 15898 4185
rect 15842 4111 15898 4120
rect 15936 4140 15988 4146
rect 15856 3670 15884 4111
rect 15936 4082 15988 4088
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15948 3058 15976 4082
rect 16132 3670 16160 5102
rect 16224 4690 16252 12378
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16316 11354 16344 12174
rect 16408 11898 16436 12242
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16500 11778 16528 14554
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16592 14074 16620 14350
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 12442 16620 13262
rect 16684 12850 16712 15030
rect 16776 13297 16804 18770
rect 16960 18698 16988 19246
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 17144 18329 17172 19178
rect 17328 18970 17356 22000
rect 17696 19394 17724 22000
rect 18064 19802 18092 22000
rect 18432 20754 18460 22000
rect 18432 20726 18736 20754
rect 18602 20632 18658 20641
rect 18602 20567 18658 20576
rect 17604 19366 17724 19394
rect 17972 19774 18092 19802
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17604 18426 17632 19366
rect 17684 19304 17736 19310
rect 17682 19272 17684 19281
rect 17736 19272 17738 19281
rect 17682 19207 17738 19216
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17130 18320 17186 18329
rect 17130 18255 17186 18264
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17512 17241 17540 18158
rect 17498 17232 17554 17241
rect 17498 17167 17554 17176
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15162 16896 15846
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 13802 16988 14350
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 16960 13530 16988 13738
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16762 13288 16818 13297
rect 16762 13223 16818 13232
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16500 11750 16620 11778
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16396 11144 16448 11150
rect 16592 11098 16620 11750
rect 16396 11086 16448 11092
rect 16408 10538 16436 11086
rect 16500 11070 16620 11098
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16408 10266 16436 10474
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16316 4729 16344 10202
rect 16396 9376 16448 9382
rect 16394 9344 16396 9353
rect 16448 9344 16450 9353
rect 16394 9279 16450 9288
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16408 7750 16436 8434
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7342 16436 7686
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16302 4720 16358 4729
rect 16212 4684 16264 4690
rect 16408 4690 16436 6870
rect 16302 4655 16358 4664
rect 16396 4684 16448 4690
rect 16212 4626 16264 4632
rect 16396 4626 16448 4632
rect 16224 3942 16252 4626
rect 16500 4078 16528 11070
rect 16684 10810 16712 12650
rect 16776 12238 16804 13223
rect 16960 12850 16988 13330
rect 17040 13184 17092 13190
rect 17038 13152 17040 13161
rect 17092 13152 17094 13161
rect 17038 13087 17094 13096
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16854 12744 16910 12753
rect 16854 12679 16856 12688
rect 16908 12679 16910 12688
rect 16856 12650 16908 12656
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16960 12170 16988 12786
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16776 11257 16804 11766
rect 17052 11286 17080 13087
rect 17040 11280 17092 11286
rect 16762 11248 16818 11257
rect 17040 11222 17092 11228
rect 16762 11183 16818 11192
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16776 10470 16804 11183
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10606 16988 11086
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16764 10464 16816 10470
rect 16670 10432 16726 10441
rect 16764 10406 16816 10412
rect 16670 10367 16726 10376
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8401 16620 9318
rect 16684 9110 16712 10367
rect 16868 9761 16896 10542
rect 16854 9752 16910 9761
rect 16854 9687 16910 9696
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16776 9110 16804 9522
rect 16868 9194 16896 9687
rect 16946 9616 17002 9625
rect 16946 9551 17002 9560
rect 16960 9382 16988 9551
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16868 9166 16988 9194
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16762 8800 16818 8809
rect 16762 8735 16818 8744
rect 16776 8401 16804 8735
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16578 8392 16634 8401
rect 16578 8327 16634 8336
rect 16762 8392 16818 8401
rect 16762 8327 16818 8336
rect 16762 7984 16818 7993
rect 16672 7948 16724 7954
rect 16868 7954 16896 8570
rect 16762 7919 16818 7928
rect 16856 7948 16908 7954
rect 16672 7890 16724 7896
rect 16684 7732 16712 7890
rect 16776 7834 16804 7919
rect 16856 7890 16908 7896
rect 16776 7806 16896 7834
rect 16764 7744 16816 7750
rect 16684 7704 16764 7732
rect 16764 7686 16816 7692
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16684 5642 16712 6122
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16408 3466 16436 3878
rect 16500 3670 16528 4014
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16592 3534 16620 5170
rect 16684 4622 16712 5578
rect 16868 5030 16896 7806
rect 16960 5166 16988 9166
rect 17144 8634 17172 16050
rect 17236 12345 17264 16594
rect 17512 14958 17540 17167
rect 17972 16250 18000 19774
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18340 18834 18368 19246
rect 18616 19242 18644 20567
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18708 18986 18736 20726
rect 18800 19310 18828 22000
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18708 18958 18828 18986
rect 18694 18864 18750 18873
rect 18328 18828 18380 18834
rect 18694 18799 18750 18808
rect 18328 18770 18380 18776
rect 18708 18766 18736 18799
rect 18144 18760 18196 18766
rect 18142 18728 18144 18737
rect 18696 18760 18748 18766
rect 18196 18728 18198 18737
rect 18696 18702 18748 18708
rect 18142 18663 18198 18672
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 18604 15972 18656 15978
rect 18604 15914 18656 15920
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17604 14550 17632 15370
rect 17682 15192 17738 15201
rect 17682 15127 17738 15136
rect 17696 14550 17724 15127
rect 17972 14958 18000 15846
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18418 14920 18474 14929
rect 18418 14855 18474 14864
rect 18432 14822 18460 14855
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 18524 14482 18552 15642
rect 18616 15162 18644 15914
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18708 14822 18736 17750
rect 18800 15502 18828 18958
rect 18984 18766 19012 22607
rect 19062 22264 19118 22273
rect 19062 22199 19118 22208
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19076 18698 19104 22199
rect 19154 22000 19210 22800
rect 19522 22000 19578 22800
rect 19890 22000 19946 22800
rect 20350 22000 20406 22800
rect 20718 22000 20774 22800
rect 21086 22000 21142 22800
rect 21454 22000 21510 22800
rect 21822 22000 21878 22800
rect 22190 22000 22246 22800
rect 22558 22000 22614 22800
rect 19168 19854 19196 22000
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19352 19922 19380 20198
rect 19536 19922 19564 22000
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19168 18970 19196 19790
rect 19352 19174 19380 19858
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19352 18816 19380 19110
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19432 18828 19484 18834
rect 19352 18788 19432 18816
rect 19432 18770 19484 18776
rect 19064 18692 19116 18698
rect 19064 18634 19116 18640
rect 19444 17202 19472 18770
rect 19536 18222 19564 18906
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 19444 16538 19472 17002
rect 19536 16658 19564 18158
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19444 16510 19564 16538
rect 19536 16182 19564 16510
rect 19524 16176 19576 16182
rect 19524 16118 19576 16124
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18880 15088 18932 15094
rect 18878 15056 18880 15065
rect 18932 15056 18934 15065
rect 18788 15020 18840 15026
rect 18878 14991 18934 15000
rect 18788 14962 18840 14968
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 17406 14376 17462 14385
rect 17406 14311 17462 14320
rect 17420 13802 17448 14311
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 13938 17908 14214
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 17408 13796 17460 13802
rect 17408 13738 17460 13744
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17328 12730 17356 13670
rect 17328 12702 17448 12730
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17222 12336 17278 12345
rect 17222 12271 17278 12280
rect 17236 9382 17264 12271
rect 17328 12102 17356 12582
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17420 11558 17448 12702
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17316 11144 17368 11150
rect 17314 11112 17316 11121
rect 17368 11112 17370 11121
rect 17314 11047 17370 11056
rect 17314 10976 17370 10985
rect 17314 10911 17370 10920
rect 17328 10742 17356 10911
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 17512 10656 17540 13670
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17604 12306 17632 13398
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17420 10628 17540 10656
rect 17420 9897 17448 10628
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17512 10062 17540 10474
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17406 9888 17462 9897
rect 17406 9823 17462 9832
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17328 9081 17356 9454
rect 17314 9072 17370 9081
rect 17314 9007 17370 9016
rect 17132 8628 17184 8634
rect 17420 8616 17448 9823
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17132 8570 17184 8576
rect 17236 8588 17448 8616
rect 17236 8514 17264 8588
rect 17144 8486 17264 8514
rect 17408 8492 17460 8498
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17052 7478 17080 8298
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17052 6458 17080 6598
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16776 4162 16804 4966
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16684 4134 16804 4162
rect 16684 4078 16712 4134
rect 16868 4078 16896 4558
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16960 4026 16988 4626
rect 17052 4146 17080 4694
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16960 3998 17080 4026
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3738 16896 3878
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 16028 2984 16080 2990
rect 15856 2932 16028 2938
rect 15856 2926 16080 2932
rect 15856 2922 16068 2926
rect 15844 2916 16068 2922
rect 15896 2910 16068 2916
rect 15844 2858 15896 2864
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15488 1414 15700 1442
rect 15844 1420 15896 1426
rect 15488 800 15516 1414
rect 15844 1362 15896 1368
rect 15856 800 15884 1362
rect 16316 898 16344 3334
rect 16592 2922 16620 3470
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16500 2650 16528 2790
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16776 2582 16804 2926
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 16868 2514 16896 3470
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16224 870 16344 898
rect 16224 800 16252 870
rect 16592 800 16620 2314
rect 16960 800 16988 3062
rect 17052 2514 17080 3998
rect 17144 3534 17172 8486
rect 17408 8434 17460 8440
rect 17420 8378 17448 8434
rect 17236 8350 17448 8378
rect 17236 7206 17264 8350
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 8090 17448 8230
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17314 7712 17370 7721
rect 17314 7647 17370 7656
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 6254 17264 7142
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17328 5681 17356 7647
rect 17314 5672 17370 5681
rect 17314 5607 17370 5616
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17236 3194 17264 3606
rect 17328 3534 17356 4082
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17328 3194 17356 3470
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17420 2990 17448 5238
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17512 2825 17540 9658
rect 17604 5234 17632 11494
rect 17696 11354 17724 12718
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17788 10962 17816 12650
rect 17880 12374 17908 13874
rect 18328 13864 18380 13870
rect 18326 13832 18328 13841
rect 18380 13832 18382 13841
rect 18326 13767 18382 13776
rect 18432 13530 18460 13874
rect 18524 13818 18552 13942
rect 18524 13790 18644 13818
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17972 12850 18000 13330
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12986 18552 13670
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 18616 12646 18644 13790
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18708 12986 18736 13738
rect 18800 13190 18828 14962
rect 18878 13968 18934 13977
rect 18878 13903 18934 13912
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17880 11762 17908 12310
rect 17972 11898 18000 12582
rect 18708 12442 18736 12786
rect 18788 12708 18840 12714
rect 18788 12650 18840 12656
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 11082 17908 11698
rect 18432 11626 18460 11766
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18524 11257 18552 11494
rect 18510 11248 18566 11257
rect 18510 11183 18566 11192
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17788 10934 17908 10962
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17774 9616 17830 9625
rect 17696 8650 17724 9590
rect 17774 9551 17830 9560
rect 17788 8974 17816 9551
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17696 8622 17816 8650
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17696 8022 17724 8502
rect 17788 8430 17816 8622
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17880 7857 17908 10934
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18248 10577 18276 10678
rect 18234 10568 18290 10577
rect 18234 10503 18290 10512
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17972 9178 18000 10134
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17972 8498 18000 9114
rect 18524 9042 18552 11086
rect 18616 9178 18644 12038
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18708 10538 18736 11698
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18708 10266 18736 10474
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18800 9518 18828 12650
rect 18892 12646 18920 13903
rect 18880 12640 18932 12646
rect 18984 12628 19012 15506
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19076 13530 19104 13874
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19168 12714 19196 15574
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19260 14482 19288 15302
rect 19352 14550 19380 15914
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 18984 12600 19104 12628
rect 18880 12582 18932 12588
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18892 9654 18920 11086
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18786 9344 18842 9353
rect 18708 9302 18786 9330
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18512 8832 18564 8838
rect 18604 8832 18656 8838
rect 18512 8774 18564 8780
rect 18602 8800 18604 8809
rect 18656 8800 18658 8809
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18524 8430 18552 8774
rect 18602 8735 18658 8744
rect 18602 8664 18658 8673
rect 18602 8599 18604 8608
rect 18656 8599 18658 8608
rect 18604 8570 18656 8576
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 17866 7848 17922 7857
rect 17866 7783 17922 7792
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7410 17724 7686
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 18524 7342 18552 7890
rect 18616 7886 18644 8434
rect 18708 8022 18736 9302
rect 18786 9279 18842 9288
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18892 8514 18920 9114
rect 18800 8486 18920 8514
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18694 7848 18750 7857
rect 18694 7783 18750 7792
rect 18602 7712 18658 7721
rect 18602 7647 18658 7656
rect 18616 7546 18644 7647
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18156 6934 18184 7142
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6186 17908 6802
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 17972 5914 18000 6870
rect 18420 6860 18472 6866
rect 18524 6848 18552 7278
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18472 6820 18552 6848
rect 18420 6802 18472 6808
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17684 5160 17736 5166
rect 17590 5128 17646 5137
rect 17684 5102 17736 5108
rect 17590 5063 17646 5072
rect 17498 2816 17554 2825
rect 17498 2751 17554 2760
rect 17604 2514 17632 5063
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17512 1426 17540 2246
rect 17500 1420 17552 1426
rect 17500 1362 17552 1368
rect 17604 1170 17632 2246
rect 17420 1142 17632 1170
rect 17420 800 17448 1142
rect 4158 232 4214 241
rect 4158 167 4214 176
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17696 241 17724 5102
rect 17880 4978 17908 5850
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17972 5545 18000 5646
rect 17958 5536 18014 5545
rect 17958 5471 18014 5480
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 18512 5228 18564 5234
rect 17972 5098 18000 5199
rect 18512 5170 18564 5176
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 17880 4950 18000 4978
rect 17972 4049 18000 4950
rect 18064 4826 18092 5034
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18432 4826 18460 4966
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18524 4622 18552 5170
rect 18616 5137 18644 7142
rect 18602 5128 18658 5137
rect 18602 5063 18658 5072
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17958 4040 18014 4049
rect 18524 4010 18552 4558
rect 17958 3975 18014 3984
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 17972 3194 18000 3538
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18420 2984 18472 2990
rect 18418 2952 18420 2961
rect 18472 2952 18474 2961
rect 17960 2916 18012 2922
rect 18418 2887 18474 2896
rect 17960 2858 18012 2864
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17788 800 17816 2518
rect 17972 1442 18000 2858
rect 18524 2650 18552 3538
rect 18616 3398 18644 4966
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18708 2990 18736 7783
rect 18800 5914 18828 8486
rect 18984 7818 19012 11630
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18800 5030 18828 5850
rect 18892 5370 18920 7210
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18694 2816 18750 2825
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18616 2553 18644 2790
rect 18694 2751 18750 2760
rect 18602 2544 18658 2553
rect 18708 2514 18736 2751
rect 18800 2650 18828 4762
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18892 3942 18920 4626
rect 18972 4616 19024 4622
rect 18970 4584 18972 4593
rect 19024 4584 19026 4593
rect 18970 4519 19026 4528
rect 18970 4448 19026 4457
rect 18970 4383 19026 4392
rect 18984 4282 19012 4383
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18984 3534 19012 4014
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 19076 3380 19104 12600
rect 19260 12306 19288 13330
rect 19352 12986 19380 13670
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19444 12866 19472 15982
rect 19536 13734 19564 16118
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19352 12838 19472 12866
rect 19352 12646 19380 12838
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19444 12442 19472 12650
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19248 12300 19300 12306
rect 19300 12260 19380 12288
rect 19248 12242 19300 12248
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 19168 11234 19196 11766
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 11354 19288 11494
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19168 11206 19288 11234
rect 19352 11218 19380 12260
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19168 10198 19196 11086
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19260 9450 19288 11206
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19444 9654 19472 11222
rect 19522 11112 19578 11121
rect 19522 11047 19578 11056
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 8090 19196 8774
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19154 7984 19210 7993
rect 19154 7919 19210 7928
rect 19168 7002 19196 7919
rect 19260 7206 19288 8978
rect 19352 8974 19380 9522
rect 19432 9104 19484 9110
rect 19536 9081 19564 11047
rect 19628 11014 19656 19178
rect 19812 18834 19840 19858
rect 19904 19310 19932 22000
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19812 17746 19840 18770
rect 19890 18728 19946 18737
rect 19890 18663 19946 18672
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19904 17338 19932 18663
rect 20364 18630 20392 22000
rect 20534 21448 20590 21457
rect 20534 21383 20590 21392
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20456 19310 20484 19858
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18442 20392 18566
rect 20272 18414 20392 18442
rect 20272 18290 20300 18414
rect 20456 18306 20484 19246
rect 20548 18902 20576 21383
rect 20732 21162 20760 22000
rect 20810 21856 20866 21865
rect 20810 21791 20866 21800
rect 20640 21134 20760 21162
rect 20640 20262 20668 21134
rect 20718 21040 20774 21049
rect 20718 20975 20774 20984
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20732 19310 20760 20975
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20364 18278 20484 18306
rect 20824 18290 20852 21791
rect 21100 18970 21128 22000
rect 21468 19990 21496 22000
rect 21456 19984 21508 19990
rect 21456 19926 21508 19932
rect 21836 19854 21864 22000
rect 22204 20058 22232 22000
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 22572 18358 22600 22000
rect 22560 18352 22612 18358
rect 21086 18320 21142 18329
rect 20812 18284 20864 18290
rect 20364 18222 20392 18278
rect 22560 18294 22612 18300
rect 21086 18255 21142 18264
rect 20812 18226 20864 18232
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19706 15464 19762 15473
rect 19706 15399 19762 15408
rect 19720 15162 19748 15399
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19708 14816 19760 14822
rect 19706 14784 19708 14793
rect 19760 14784 19762 14793
rect 19706 14719 19762 14728
rect 19812 13954 19840 17070
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19904 14550 19932 15438
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 14074 19932 14350
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19996 13977 20024 18090
rect 20258 17912 20314 17921
rect 21100 17882 21128 18255
rect 20258 17847 20314 17856
rect 21088 17876 21140 17882
rect 20272 17338 20300 17847
rect 21088 17818 21140 17824
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20628 17128 20680 17134
rect 20350 17096 20406 17105
rect 20628 17070 20680 17076
rect 20350 17031 20406 17040
rect 20364 16250 20392 17031
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20640 16114 20668 17070
rect 20916 16658 20944 17546
rect 21178 17504 21234 17513
rect 21178 17439 21234 17448
rect 21192 17338 21220 17439
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21100 16697 21128 16730
rect 21086 16688 21142 16697
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20904 16652 20956 16658
rect 21086 16623 21142 16632
rect 20904 16594 20956 16600
rect 20718 16280 20774 16289
rect 20718 16215 20720 16224
rect 20772 16215 20774 16224
rect 20720 16186 20772 16192
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20088 14550 20116 15506
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 19720 13926 19840 13954
rect 19982 13968 20038 13977
rect 19720 11898 19748 13926
rect 19982 13903 20038 13912
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19996 12986 20024 13738
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19892 12912 19944 12918
rect 20088 12866 20116 13466
rect 19944 12860 20116 12866
rect 19892 12854 20116 12860
rect 19904 12838 20116 12854
rect 20088 12782 20116 12838
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19720 10470 19748 11698
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19812 9518 19840 12378
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 19904 10810 19932 11222
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 20180 10606 20208 15982
rect 20628 15904 20680 15910
rect 20258 15872 20314 15881
rect 20628 15846 20680 15852
rect 20258 15807 20314 15816
rect 20272 15706 20300 15807
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20272 12753 20300 14826
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20364 13977 20392 14758
rect 20456 14385 20484 15302
rect 20640 15201 20668 15846
rect 20626 15192 20682 15201
rect 20626 15127 20682 15136
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20442 14376 20498 14385
rect 20442 14311 20498 14320
rect 20350 13968 20406 13977
rect 20350 13903 20406 13912
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 12782 20392 13670
rect 20456 13190 20484 13874
rect 20444 13184 20496 13190
rect 20548 13161 20576 15030
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 13938 20760 14894
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20628 13864 20680 13870
rect 20626 13832 20628 13841
rect 20680 13832 20682 13841
rect 20626 13767 20682 13776
rect 20628 13184 20680 13190
rect 20444 13126 20496 13132
rect 20534 13152 20590 13161
rect 20352 12776 20404 12782
rect 20258 12744 20314 12753
rect 20352 12718 20404 12724
rect 20258 12679 20314 12688
rect 20456 12374 20484 13126
rect 20628 13126 20680 13132
rect 20534 13087 20590 13096
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 11286 20392 11698
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 19800 9512 19852 9518
rect 19628 9460 19800 9466
rect 19628 9454 19852 9460
rect 19628 9438 19840 9454
rect 19432 9046 19484 9052
rect 19522 9072 19578 9081
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19168 5166 19196 6394
rect 19260 6186 19288 6598
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19260 5710 19288 6122
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 19260 5234 19288 5646
rect 19352 5370 19380 8366
rect 19444 8022 19472 9046
rect 19522 9007 19578 9016
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19444 7478 19472 7958
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19536 7206 19564 9007
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6458 19472 6802
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19432 5840 19484 5846
rect 19536 5828 19564 6734
rect 19628 6254 19656 9438
rect 19904 9382 19932 10542
rect 20364 10266 20392 10542
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20350 10160 20406 10169
rect 19984 10124 20036 10130
rect 20350 10095 20406 10104
rect 19984 10066 20036 10072
rect 19996 9722 20024 10066
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19812 8498 19840 9318
rect 19904 8537 19932 9318
rect 19996 8974 20024 9386
rect 20088 9178 20116 9998
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19890 8528 19946 8537
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19800 8492 19852 8498
rect 19890 8463 19946 8472
rect 19800 8434 19852 8440
rect 19720 7342 19748 8434
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19904 7546 19932 8298
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19720 7002 19748 7278
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5846 19656 6054
rect 19484 5800 19564 5828
rect 19616 5840 19668 5846
rect 19432 5782 19484 5788
rect 19616 5782 19668 5788
rect 19720 5692 19748 6802
rect 19444 5664 19748 5692
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5250 19472 5664
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19352 5222 19472 5250
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 19246 5128 19302 5137
rect 19246 5063 19302 5072
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 18892 3352 19104 3380
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18602 2479 18658 2488
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1414 18184 1442
rect 18156 800 18184 1414
rect 18524 800 18552 2314
rect 18708 1737 18736 2450
rect 18694 1728 18750 1737
rect 18694 1663 18750 1672
rect 18800 921 18828 2586
rect 18786 912 18842 921
rect 18786 847 18842 856
rect 18892 800 18920 3352
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18984 2446 19012 2994
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 17682 232 17738 241
rect 17682 167 17738 176
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19168 513 19196 4966
rect 19260 2553 19288 5063
rect 19246 2544 19302 2553
rect 19352 2514 19380 5222
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19444 4729 19472 4966
rect 19430 4720 19486 4729
rect 19430 4655 19486 4664
rect 19536 3670 19564 5238
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 19628 4282 19656 4626
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19628 3618 19656 4218
rect 19628 3590 19748 3618
rect 19720 3534 19748 3590
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19812 2514 19840 7142
rect 19996 4826 20024 8910
rect 20180 8498 20208 9318
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20180 7750 20208 8434
rect 20272 8090 20300 8842
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 7002 20300 7142
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20074 6352 20130 6361
rect 20180 6322 20208 6802
rect 20074 6287 20130 6296
rect 20168 6316 20220 6322
rect 20088 5914 20116 6287
rect 20168 6258 20220 6264
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20088 5166 20116 5510
rect 20076 5160 20128 5166
rect 20076 5102 20128 5108
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 19246 2479 19302 2488
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 20180 2145 20208 6122
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20272 2961 20300 5646
rect 20258 2952 20314 2961
rect 20258 2887 20314 2896
rect 20166 2136 20222 2145
rect 20166 2071 20222 2080
rect 20364 800 20392 10095
rect 20456 8673 20484 10406
rect 20548 9382 20576 12038
rect 20640 11937 20668 13126
rect 20626 11928 20682 11937
rect 20626 11863 20682 11872
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10742 20760 10950
rect 20824 10742 20852 16594
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20916 13530 20944 15982
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21100 13569 21128 15302
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21086 13560 21142 13569
rect 20904 13524 20956 13530
rect 21086 13495 21142 13504
rect 20904 13466 20956 13472
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20916 11762 20944 13330
rect 21192 12345 21220 14214
rect 21178 12336 21234 12345
rect 20996 12300 21048 12306
rect 21178 12271 21234 12280
rect 20996 12242 21048 12248
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20812 10736 20864 10742
rect 20812 10678 20864 10684
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20442 8664 20498 8673
rect 20442 8599 20498 8608
rect 20548 8362 20576 9046
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20640 8430 20668 8978
rect 20824 8634 20852 10542
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20456 6458 20484 7346
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20456 5234 20484 6394
rect 20548 5846 20576 8298
rect 20640 6254 20668 8366
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20548 3466 20576 5102
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20640 1329 20668 6190
rect 20824 5658 20852 6258
rect 20732 5642 20852 5658
rect 20720 5636 20852 5642
rect 20772 5630 20852 5636
rect 20720 5578 20772 5584
rect 20732 4826 20760 5578
rect 20916 5234 20944 11154
rect 21008 10674 21036 12242
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21192 11665 21220 12038
rect 21178 11656 21234 11665
rect 21178 11591 21234 11600
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21100 11257 21128 11290
rect 21086 11248 21142 11257
rect 21086 11183 21142 11192
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 21284 4690 21312 17002
rect 21376 9654 21404 17614
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 20626 1320 20682 1329
rect 20626 1255 20682 1264
rect 21560 950 21588 9522
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 20720 944 20772 950
rect 20720 886 20772 892
rect 21548 944 21600 950
rect 21548 886 21600 892
rect 20732 800 20760 886
rect 22204 800 22232 4626
rect 22572 800 22600 10678
rect 19154 504 19210 513
rect 19154 439 19210 448
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
<< via2 >>
rect 18970 22616 19026 22672
rect 2962 20576 3018 20632
rect 2962 19216 3018 19272
rect 1674 18672 1730 18728
rect 1306 18128 1362 18184
rect 2410 18400 2466 18456
rect 1950 18300 1952 18320
rect 1952 18300 2004 18320
rect 2004 18300 2006 18320
rect 1950 18264 2006 18300
rect 1950 17448 2006 17504
rect 1582 17040 1638 17096
rect 1582 16632 1638 16688
rect 1398 16496 1454 16552
rect 1950 16224 2006 16280
rect 1582 15408 1638 15464
rect 1950 14320 2006 14376
rect 1766 13912 1822 13968
rect 1582 12824 1638 12880
rect 1766 13096 1822 13152
rect 1674 12688 1730 12744
rect 1582 12280 1638 12336
rect 1674 11872 1730 11928
rect 1398 11056 1454 11112
rect 2870 18400 2926 18456
rect 3238 18964 3294 19000
rect 3238 18944 3240 18964
rect 3240 18944 3292 18964
rect 3292 18944 3294 18964
rect 3422 18536 3478 18592
rect 2870 15816 2926 15872
rect 2226 15408 2282 15464
rect 2318 14764 2320 14784
rect 2320 14764 2372 14784
rect 2372 14764 2374 14784
rect 2318 14728 2374 14764
rect 2778 15156 2834 15192
rect 3330 17212 3332 17232
rect 3332 17212 3384 17232
rect 3384 17212 3386 17232
rect 3330 17176 3386 17212
rect 2778 15136 2780 15156
rect 2780 15136 2832 15156
rect 2832 15136 2834 15156
rect 2778 13504 2834 13560
rect 2410 13368 2466 13424
rect 1306 8744 1362 8800
rect 3054 11600 3110 11656
rect 2870 11192 2926 11248
rect 2778 9424 2834 9480
rect 3698 20984 3754 21040
rect 4066 20204 4068 20224
rect 4068 20204 4120 20224
rect 4120 20204 4122 20224
rect 4066 20168 4122 20204
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 3698 18264 3754 18320
rect 3698 18148 3754 18184
rect 3698 18128 3700 18148
rect 3700 18128 3752 18148
rect 3752 18128 3754 18148
rect 3606 17992 3662 18048
rect 3606 17856 3662 17912
rect 3974 19352 4030 19408
rect 3974 18808 4030 18864
rect 3974 18536 4030 18592
rect 4066 17756 4068 17776
rect 4068 17756 4120 17776
rect 4120 17756 4122 17776
rect 4066 17720 4122 17756
rect 3790 15036 3792 15056
rect 3792 15036 3844 15056
rect 3844 15036 3846 15056
rect 3790 15000 3846 15036
rect 2686 7112 2742 7168
rect 4802 19760 4858 19816
rect 4710 19080 4766 19136
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4342 17992 4398 18048
rect 4710 17992 4766 18048
rect 4526 17620 4528 17640
rect 4528 17620 4580 17640
rect 4580 17620 4582 17640
rect 4526 17584 4582 17620
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3422 10512 3478 10568
rect 2686 5480 2742 5536
rect 2318 2488 2374 2544
rect 1766 856 1822 912
rect 2962 2916 3018 2952
rect 2962 2896 2964 2916
rect 2964 2896 3016 2916
rect 3016 2896 3018 2916
rect 2778 2488 2834 2544
rect 2502 1672 2558 1728
rect 3422 8336 3478 8392
rect 3422 7404 3478 7440
rect 3422 7384 3424 7404
rect 3424 7384 3476 7404
rect 3476 7384 3478 7404
rect 4894 17176 4950 17232
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4894 15852 4896 15872
rect 4896 15852 4948 15872
rect 4948 15852 4950 15872
rect 4894 15816 4950 15852
rect 4802 15136 4858 15192
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 5354 17584 5410 17640
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 3790 10804 3846 10840
rect 3790 10784 3792 10804
rect 3792 10784 3844 10804
rect 3844 10784 3846 10804
rect 3790 10648 3846 10704
rect 4618 11600 4674 11656
rect 4066 10784 4122 10840
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4434 10548 4436 10568
rect 4436 10548 4488 10568
rect 4488 10548 4490 10568
rect 4434 10512 4490 10548
rect 4066 9968 4122 10024
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 3514 5208 3570 5264
rect 3790 7148 3792 7168
rect 3792 7148 3844 7168
rect 3844 7148 3846 7168
rect 3790 7112 3846 7148
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4618 8336 4674 8392
rect 4066 7692 4068 7712
rect 4068 7692 4120 7712
rect 4120 7692 4122 7712
rect 4066 7656 4122 7692
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4066 7248 4122 7304
rect 3330 3032 3386 3088
rect 3238 2080 3294 2136
rect 3330 1264 3386 1320
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4066 6432 4122 6488
rect 4066 6024 4122 6080
rect 3974 5616 4030 5672
rect 4618 6024 4674 6080
rect 4986 11600 5042 11656
rect 4986 9832 5042 9888
rect 5998 18964 6054 19000
rect 5998 18944 6000 18964
rect 6000 18944 6052 18964
rect 6052 18944 6054 18964
rect 5998 17584 6054 17640
rect 5354 15136 5410 15192
rect 5814 15408 5870 15464
rect 5630 14456 5686 14512
rect 5262 10648 5318 10704
rect 5170 10240 5226 10296
rect 5078 9424 5134 9480
rect 5078 8336 5134 8392
rect 5078 6568 5134 6624
rect 4986 5888 5042 5944
rect 4250 5480 4306 5536
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4250 5208 4306 5264
rect 4066 4800 4122 4856
rect 4066 4392 4122 4448
rect 4066 3304 4122 3360
rect 3790 448 3846 504
rect 6366 16360 6422 16416
rect 5630 10104 5686 10160
rect 5538 7384 5594 7440
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4526 4120 4582 4176
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 5354 4800 5410 4856
rect 4986 3712 5042 3768
rect 4894 2508 4950 2544
rect 4894 2488 4896 2508
rect 4896 2488 4948 2508
rect 4948 2488 4950 2508
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4618 1944 4674 2000
rect 5814 7384 5870 7440
rect 5998 6432 6054 6488
rect 5446 3848 5502 3904
rect 5814 4528 5870 4584
rect 5906 4256 5962 4312
rect 5814 4120 5870 4176
rect 5630 3712 5686 3768
rect 6642 17040 6698 17096
rect 6182 12416 6238 12472
rect 6182 8744 6238 8800
rect 6274 8336 6330 8392
rect 6274 7520 6330 7576
rect 6182 5788 6184 5808
rect 6184 5788 6236 5808
rect 6236 5788 6238 5808
rect 6182 5752 6238 5788
rect 6550 12280 6606 12336
rect 6458 8744 6514 8800
rect 6458 8472 6514 8528
rect 6734 14320 6790 14376
rect 6918 13252 6974 13288
rect 6918 13232 6920 13252
rect 6920 13232 6972 13252
rect 6972 13232 6974 13252
rect 7286 14728 7342 14784
rect 7010 12552 7066 12608
rect 6734 11872 6790 11928
rect 6826 11212 6882 11248
rect 6826 11192 6828 11212
rect 6828 11192 6880 11212
rect 6880 11192 6882 11212
rect 7102 11736 7158 11792
rect 7102 9152 7158 9208
rect 6550 7248 6606 7304
rect 6826 8780 6828 8800
rect 6828 8780 6880 8800
rect 6880 8780 6882 8800
rect 6826 8744 6882 8780
rect 6550 5072 6606 5128
rect 6734 6332 6736 6352
rect 6736 6332 6788 6352
rect 6788 6332 6790 6352
rect 6734 6296 6790 6332
rect 6734 6160 6790 6216
rect 6734 4664 6790 4720
rect 7010 3848 7066 3904
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8482 17856 8538 17912
rect 8574 17584 8630 17640
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 8758 17040 8814 17096
rect 8758 16632 8814 16688
rect 8758 16360 8814 16416
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7930 15408 7986 15464
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 8482 15408 8538 15464
rect 8390 14728 8446 14784
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7654 12144 7710 12200
rect 7654 12008 7710 12064
rect 7470 10004 7472 10024
rect 7472 10004 7524 10024
rect 7524 10004 7526 10024
rect 7470 9968 7526 10004
rect 7470 9832 7526 9888
rect 7470 8880 7526 8936
rect 7194 5888 7250 5944
rect 7102 3032 7158 3088
rect 7286 4800 7342 4856
rect 7562 7948 7618 7984
rect 7562 7928 7564 7948
rect 7564 7928 7616 7948
rect 7616 7928 7618 7948
rect 8482 14592 8538 14648
rect 8114 13096 8170 13152
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 8390 12688 8446 12744
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8298 10512 8354 10568
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8206 9968 8262 10024
rect 8298 9560 8354 9616
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 8114 8336 8170 8392
rect 8298 8608 8354 8664
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7562 6840 7618 6896
rect 7930 7656 7986 7712
rect 8298 8336 8354 8392
rect 8482 12416 8538 12472
rect 8850 15272 8906 15328
rect 8666 12688 8722 12744
rect 9126 18128 9182 18184
rect 9126 16532 9128 16552
rect 9128 16532 9180 16552
rect 9180 16532 9182 16552
rect 9126 16496 9182 16532
rect 9402 15136 9458 15192
rect 9310 13232 9366 13288
rect 9218 13096 9274 13152
rect 9310 12552 9366 12608
rect 8574 10784 8630 10840
rect 8666 10548 8668 10568
rect 8668 10548 8720 10568
rect 8720 10548 8722 10568
rect 8666 10512 8722 10548
rect 8666 10376 8722 10432
rect 8574 9968 8630 10024
rect 8574 9152 8630 9208
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 8206 6976 8262 7032
rect 7930 6740 7932 6760
rect 7932 6740 7984 6760
rect 7984 6740 7986 6760
rect 7930 6704 7986 6740
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7746 5616 7802 5672
rect 7470 5228 7526 5264
rect 7470 5208 7472 5228
rect 7472 5208 7524 5228
rect 7524 5208 7526 5228
rect 7654 5208 7710 5264
rect 6826 2488 6882 2544
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 9218 10920 9274 10976
rect 8942 9444 8998 9480
rect 8942 9424 8944 9444
rect 8944 9424 8996 9444
rect 8996 9424 8998 9444
rect 8942 7268 8998 7304
rect 8942 7248 8944 7268
rect 8944 7248 8996 7268
rect 8996 7248 8998 7268
rect 8850 6840 8906 6896
rect 8298 4936 8354 4992
rect 7654 4120 7710 4176
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 8206 3304 8262 3360
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8574 5208 8630 5264
rect 8482 4664 8538 4720
rect 8666 4276 8722 4312
rect 8942 4528 8998 4584
rect 8666 4256 8668 4276
rect 8668 4256 8720 4276
rect 8720 4256 8722 4276
rect 8666 4120 8722 4176
rect 8666 3848 8722 3904
rect 8574 3460 8630 3496
rect 8574 3440 8576 3460
rect 8576 3440 8628 3460
rect 8628 3440 8630 3460
rect 8574 3304 8630 3360
rect 8574 2760 8630 2816
rect 8850 3712 8906 3768
rect 9218 9288 9274 9344
rect 9678 17856 9734 17912
rect 9586 15272 9642 15328
rect 9494 11228 9496 11248
rect 9496 11228 9548 11248
rect 9548 11228 9550 11248
rect 9494 11192 9550 11228
rect 9402 10512 9458 10568
rect 9402 8064 9458 8120
rect 9126 5752 9182 5808
rect 9678 12280 9734 12336
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 9954 14612 10010 14648
rect 9954 14592 9956 14612
rect 9956 14592 10008 14612
rect 10008 14592 10010 14612
rect 9770 11192 9826 11248
rect 9770 8608 9826 8664
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11702 17992 11758 18048
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11426 17040 11482 17096
rect 11334 16788 11390 16824
rect 11334 16768 11336 16788
rect 11336 16768 11388 16788
rect 11388 16768 11390 16788
rect 11610 16496 11666 16552
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 10966 16088 11022 16144
rect 10230 13812 10232 13832
rect 10232 13812 10284 13832
rect 10284 13812 10286 13832
rect 10230 13776 10286 13812
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11150 14764 11152 14784
rect 11152 14764 11204 14784
rect 11204 14764 11206 14784
rect 11150 14728 11206 14764
rect 10230 13368 10286 13424
rect 10414 13368 10470 13424
rect 10230 12008 10286 12064
rect 10138 10376 10194 10432
rect 10046 7928 10102 7984
rect 10690 13232 10746 13288
rect 10230 8200 10286 8256
rect 9770 7520 9826 7576
rect 9678 5888 9734 5944
rect 9402 3032 9458 3088
rect 9586 3712 9642 3768
rect 10138 6876 10140 6896
rect 10140 6876 10192 6896
rect 10192 6876 10194 6896
rect 10138 6840 10194 6876
rect 10230 6024 10286 6080
rect 9954 4664 10010 4720
rect 10598 12724 10600 12744
rect 10600 12724 10652 12744
rect 10652 12724 10654 12744
rect 10598 12688 10654 12724
rect 12346 17856 12402 17912
rect 12254 17720 12310 17776
rect 12530 17176 12586 17232
rect 12254 16496 12310 16552
rect 11794 15408 11850 15464
rect 12070 15000 12126 15056
rect 11702 14864 11758 14920
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11242 13912 11298 13968
rect 11058 13640 11114 13696
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 10874 12280 10930 12336
rect 10690 11736 10746 11792
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11150 11736 11206 11792
rect 11978 14592 12034 14648
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 12070 13912 12126 13968
rect 11978 11192 12034 11248
rect 10506 8744 10562 8800
rect 10598 8200 10654 8256
rect 10506 7284 10508 7304
rect 10508 7284 10560 7304
rect 10560 7284 10562 7304
rect 10506 7248 10562 7284
rect 10690 7520 10746 7576
rect 10966 9596 10968 9616
rect 10968 9596 11020 9616
rect 11020 9596 11022 9616
rect 10966 9560 11022 9596
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 10690 4800 10746 4856
rect 10598 3848 10654 3904
rect 10598 3168 10654 3224
rect 10598 2760 10654 2816
rect 11058 8628 11114 8664
rect 11058 8608 11060 8628
rect 11060 8608 11112 8628
rect 11112 8608 11114 8628
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11702 9172 11758 9208
rect 11702 9152 11704 9172
rect 11704 9152 11756 9172
rect 11756 9152 11758 9172
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11058 6432 11114 6488
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11702 6296 11758 6352
rect 11242 5888 11298 5944
rect 11518 5888 11574 5944
rect 11886 9152 11942 9208
rect 11978 8608 12034 8664
rect 12162 13640 12218 13696
rect 12898 17992 12954 18048
rect 12990 17040 13046 17096
rect 12714 16768 12770 16824
rect 12346 12824 12402 12880
rect 12162 11600 12218 11656
rect 12162 11192 12218 11248
rect 12162 8744 12218 8800
rect 11886 6976 11942 7032
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11518 4936 11574 4992
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11978 6160 12034 6216
rect 12438 10920 12494 10976
rect 12622 14864 12678 14920
rect 12806 15544 12862 15600
rect 12806 13912 12862 13968
rect 12898 13776 12954 13832
rect 14002 16088 14058 16144
rect 13634 15272 13690 15328
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14554 17604 14610 17640
rect 14554 17584 14556 17604
rect 14556 17584 14608 17604
rect 14608 17584 14610 17604
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 12714 11328 12770 11384
rect 12898 13096 12954 13152
rect 12530 9696 12586 9752
rect 12346 7692 12348 7712
rect 12348 7692 12400 7712
rect 12400 7692 12402 7712
rect 12346 7656 12402 7692
rect 12346 7248 12402 7304
rect 13082 9560 13138 9616
rect 12806 8780 12808 8800
rect 12808 8780 12860 8800
rect 12860 8780 12862 8800
rect 12806 8744 12862 8780
rect 12622 6840 12678 6896
rect 12254 6024 12310 6080
rect 12070 5480 12126 5536
rect 11702 3712 11758 3768
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12346 4936 12402 4992
rect 12990 6840 13046 6896
rect 13082 5344 13138 5400
rect 11978 3032 12034 3088
rect 13450 12824 13506 12880
rect 13266 7112 13322 7168
rect 13266 3576 13322 3632
rect 12990 2896 13046 2952
rect 13726 10648 13782 10704
rect 14370 13504 14426 13560
rect 14278 12824 14334 12880
rect 14094 10648 14150 10704
rect 13726 9968 13782 10024
rect 13634 9560 13690 9616
rect 13818 8608 13874 8664
rect 14002 10376 14058 10432
rect 14094 9988 14150 10024
rect 14094 9968 14096 9988
rect 14096 9968 14148 9988
rect 14148 9968 14150 9988
rect 14094 8608 14150 8664
rect 13910 7284 13912 7304
rect 13912 7284 13964 7304
rect 13964 7284 13966 7304
rect 13910 7248 13966 7284
rect 14094 6976 14150 7032
rect 15290 16632 15346 16688
rect 15290 15000 15346 15056
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 15106 13776 15162 13832
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 15658 13388 15714 13424
rect 16026 13812 16028 13832
rect 16028 13812 16080 13832
rect 16080 13812 16082 13832
rect 16026 13776 16082 13812
rect 15658 13368 15660 13388
rect 15660 13368 15712 13388
rect 15712 13368 15714 13388
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14462 10648 14518 10704
rect 14462 9832 14518 9888
rect 14370 9560 14426 9616
rect 15106 10532 15162 10568
rect 15106 10512 15108 10532
rect 15108 10512 15160 10532
rect 15160 10512 15162 10532
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14738 10124 14794 10160
rect 14738 10104 14740 10124
rect 14740 10104 14792 10124
rect 14792 10104 14794 10124
rect 14922 9424 14978 9480
rect 14370 9288 14426 9344
rect 15290 9696 15346 9752
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 15198 9036 15254 9072
rect 15198 9016 15200 9036
rect 15200 9016 15252 9036
rect 15252 9016 15254 9036
rect 15106 8608 15162 8664
rect 14462 8200 14518 8256
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14462 6976 14518 7032
rect 13818 6024 13874 6080
rect 13910 5344 13966 5400
rect 13818 5072 13874 5128
rect 14094 4936 14150 4992
rect 14278 4800 14334 4856
rect 13910 4020 13912 4040
rect 13912 4020 13964 4040
rect 13964 4020 13966 4040
rect 13910 3984 13966 4020
rect 14278 3440 14334 3496
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14830 4392 14886 4448
rect 15106 4800 15162 4856
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 15934 12860 15936 12880
rect 15936 12860 15988 12880
rect 15988 12860 15990 12880
rect 15934 12824 15990 12860
rect 15474 9016 15530 9072
rect 15382 5752 15438 5808
rect 15290 3712 15346 3768
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15842 9424 15898 9480
rect 15750 8880 15806 8936
rect 15842 7384 15898 7440
rect 16026 6976 16082 7032
rect 15750 6160 15806 6216
rect 15658 5108 15660 5128
rect 15660 5108 15712 5128
rect 15712 5108 15714 5128
rect 15658 5072 15714 5108
rect 15658 4528 15714 4584
rect 15566 4120 15622 4176
rect 16118 5244 16120 5264
rect 16120 5244 16172 5264
rect 16172 5244 16174 5264
rect 16118 5208 16174 5244
rect 15842 4120 15898 4176
rect 18602 20576 18658 20632
rect 17682 19252 17684 19272
rect 17684 19252 17736 19272
rect 17736 19252 17738 19272
rect 17682 19216 17738 19252
rect 17130 18264 17186 18320
rect 17498 17176 17554 17232
rect 16762 13232 16818 13288
rect 16394 9324 16396 9344
rect 16396 9324 16448 9344
rect 16448 9324 16450 9344
rect 16394 9288 16450 9324
rect 16302 4664 16358 4720
rect 17038 13132 17040 13152
rect 17040 13132 17092 13152
rect 17092 13132 17094 13152
rect 17038 13096 17094 13132
rect 16854 12708 16910 12744
rect 16854 12688 16856 12708
rect 16856 12688 16908 12708
rect 16908 12688 16910 12708
rect 16762 11192 16818 11248
rect 16670 10376 16726 10432
rect 16854 9696 16910 9752
rect 16946 9560 17002 9616
rect 16762 8744 16818 8800
rect 16578 8336 16634 8392
rect 16762 8336 16818 8392
rect 16762 7928 16818 7984
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18694 18808 18750 18864
rect 18142 18708 18144 18728
rect 18144 18708 18196 18728
rect 18196 18708 18198 18728
rect 18142 18672 18198 18708
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 17682 15136 17738 15192
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18418 14864 18474 14920
rect 19062 22208 19118 22264
rect 18878 15036 18880 15056
rect 18880 15036 18932 15056
rect 18932 15036 18934 15056
rect 18878 15000 18934 15036
rect 17406 14320 17462 14376
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 17222 12280 17278 12336
rect 17314 11092 17316 11112
rect 17316 11092 17368 11112
rect 17368 11092 17370 11112
rect 17314 11056 17370 11092
rect 17314 10920 17370 10976
rect 17406 9832 17462 9888
rect 17314 9016 17370 9072
rect 17314 7656 17370 7712
rect 17314 5616 17370 5672
rect 18326 13812 18328 13832
rect 18328 13812 18380 13832
rect 18380 13812 18382 13832
rect 18326 13776 18382 13812
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18878 13912 18934 13968
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18510 11192 18566 11248
rect 17774 9560 17830 9616
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18234 10512 18290 10568
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18602 8780 18604 8800
rect 18604 8780 18656 8800
rect 18656 8780 18658 8800
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18602 8744 18658 8780
rect 18602 8628 18658 8664
rect 18602 8608 18604 8628
rect 18604 8608 18656 8628
rect 18656 8608 18658 8628
rect 17866 7792 17922 7848
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18786 9288 18842 9344
rect 18694 7792 18750 7848
rect 18602 7656 18658 7712
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17590 5072 17646 5128
rect 17498 2760 17554 2816
rect 4158 176 4214 232
rect 17958 5480 18014 5536
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 17958 5208 18014 5264
rect 18602 5072 18658 5128
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17958 3984 18014 4040
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18418 2932 18420 2952
rect 18420 2932 18472 2952
rect 18472 2932 18474 2952
rect 18418 2896 18474 2932
rect 18694 2760 18750 2816
rect 18602 2488 18658 2544
rect 18970 4564 18972 4584
rect 18972 4564 19024 4584
rect 19024 4564 19026 4584
rect 18970 4528 19026 4564
rect 18970 4392 19026 4448
rect 19522 11056 19578 11112
rect 19154 7928 19210 7984
rect 19890 18672 19946 18728
rect 20534 21392 20590 21448
rect 20810 21800 20866 21856
rect 20718 20984 20774 21040
rect 21086 18264 21142 18320
rect 19706 15408 19762 15464
rect 19706 14764 19708 14784
rect 19708 14764 19760 14784
rect 19760 14764 19762 14784
rect 19706 14728 19762 14764
rect 20258 17856 20314 17912
rect 20350 17040 20406 17096
rect 21178 17448 21234 17504
rect 21086 16632 21142 16688
rect 20718 16244 20774 16280
rect 20718 16224 20720 16244
rect 20720 16224 20772 16244
rect 20772 16224 20774 16244
rect 19982 13912 20038 13968
rect 20258 15816 20314 15872
rect 20626 15136 20682 15192
rect 20442 14320 20498 14376
rect 20350 13912 20406 13968
rect 20626 13812 20628 13832
rect 20628 13812 20680 13832
rect 20680 13812 20682 13832
rect 20626 13776 20682 13812
rect 20258 12688 20314 12744
rect 20534 13096 20590 13152
rect 19522 9016 19578 9072
rect 20350 10104 20406 10160
rect 19890 8472 19946 8528
rect 19246 5072 19302 5128
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18694 1672 18750 1728
rect 18786 856 18842 912
rect 17682 176 17738 232
rect 19246 2488 19302 2544
rect 19430 4664 19486 4720
rect 20074 6296 20130 6352
rect 20258 2896 20314 2952
rect 20166 2080 20222 2136
rect 20626 11872 20682 11928
rect 21086 13504 21142 13560
rect 21178 12280 21234 12336
rect 20442 8608 20498 8664
rect 21178 11600 21234 11656
rect 21086 11192 21142 11248
rect 20626 1264 20682 1320
rect 19154 448 19210 504
<< metal3 >>
rect 0 22584 800 22704
rect 18965 22674 19031 22677
rect 22000 22674 22800 22704
rect 18965 22672 22800 22674
rect 18965 22616 18970 22672
rect 19026 22616 22800 22672
rect 18965 22614 22800 22616
rect 18965 22611 19031 22614
rect 22000 22584 22800 22614
rect 0 22176 800 22296
rect 19057 22266 19123 22269
rect 22000 22266 22800 22296
rect 19057 22264 22800 22266
rect 19057 22208 19062 22264
rect 19118 22208 22800 22264
rect 19057 22206 22800 22208
rect 19057 22203 19123 22206
rect 22000 22176 22800 22206
rect 0 21768 800 21888
rect 20805 21858 20871 21861
rect 22000 21858 22800 21888
rect 20805 21856 22800 21858
rect 20805 21800 20810 21856
rect 20866 21800 22800 21856
rect 20805 21798 22800 21800
rect 20805 21795 20871 21798
rect 22000 21768 22800 21798
rect 0 21360 800 21480
rect 20529 21450 20595 21453
rect 22000 21450 22800 21480
rect 20529 21448 22800 21450
rect 20529 21392 20534 21448
rect 20590 21392 22800 21448
rect 20529 21390 22800 21392
rect 20529 21387 20595 21390
rect 22000 21360 22800 21390
rect 0 21042 800 21072
rect 3693 21042 3759 21045
rect 0 21040 3759 21042
rect 0 20984 3698 21040
rect 3754 20984 3759 21040
rect 0 20982 3759 20984
rect 0 20952 800 20982
rect 3693 20979 3759 20982
rect 20713 21042 20779 21045
rect 22000 21042 22800 21072
rect 20713 21040 22800 21042
rect 20713 20984 20718 21040
rect 20774 20984 22800 21040
rect 20713 20982 22800 20984
rect 20713 20979 20779 20982
rect 22000 20952 22800 20982
rect 0 20634 800 20664
rect 2957 20634 3023 20637
rect 0 20632 3023 20634
rect 0 20576 2962 20632
rect 3018 20576 3023 20632
rect 0 20574 3023 20576
rect 0 20544 800 20574
rect 2957 20571 3023 20574
rect 18597 20634 18663 20637
rect 22000 20634 22800 20664
rect 18597 20632 22800 20634
rect 18597 20576 18602 20632
rect 18658 20576 22800 20632
rect 18597 20574 22800 20576
rect 18597 20571 18663 20574
rect 22000 20544 22800 20574
rect 0 20226 800 20256
rect 4061 20226 4127 20229
rect 0 20224 4127 20226
rect 0 20168 4066 20224
rect 4122 20168 4127 20224
rect 0 20166 4127 20168
rect 0 20136 800 20166
rect 4061 20163 4127 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22000 20136 22800 20256
rect 14672 20095 14992 20096
rect 0 19818 800 19848
rect 4797 19818 4863 19821
rect 0 19816 4863 19818
rect 0 19760 4802 19816
rect 4858 19760 4863 19816
rect 0 19758 4863 19760
rect 0 19728 800 19758
rect 4797 19755 4863 19758
rect 22000 19728 22800 19848
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19410 800 19440
rect 3969 19410 4035 19413
rect 0 19408 4035 19410
rect 0 19352 3974 19408
rect 4030 19352 4035 19408
rect 0 19350 4035 19352
rect 0 19320 800 19350
rect 3969 19347 4035 19350
rect 22000 19320 22800 19440
rect 2957 19274 3023 19277
rect 17677 19274 17743 19277
rect 2957 19272 17743 19274
rect 2957 19216 2962 19272
rect 3018 19216 17682 19272
rect 17738 19216 17743 19272
rect 2957 19214 17743 19216
rect 2957 19211 3023 19214
rect 17677 19211 17743 19214
rect 0 19138 800 19168
rect 4705 19138 4771 19141
rect 5022 19138 5028 19140
rect 0 19078 3112 19138
rect 0 19048 800 19078
rect 0 18730 800 18760
rect 1669 18730 1735 18733
rect 0 18728 1735 18730
rect 0 18672 1674 18728
rect 1730 18672 1735 18728
rect 0 18670 1735 18672
rect 3052 18730 3112 19078
rect 4705 19136 5028 19138
rect 4705 19080 4710 19136
rect 4766 19080 5028 19136
rect 4705 19078 5028 19080
rect 4705 19075 4771 19078
rect 5022 19076 5028 19078
rect 5092 19076 5098 19140
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 22000 19048 22800 19168
rect 14672 19007 14992 19008
rect 3233 19002 3299 19005
rect 5993 19002 6059 19005
rect 3233 19000 6059 19002
rect 3233 18944 3238 19000
rect 3294 18944 5998 19000
rect 6054 18944 6059 19000
rect 3233 18942 6059 18944
rect 3233 18939 3299 18942
rect 5993 18939 6059 18942
rect 3969 18866 4035 18869
rect 18689 18866 18755 18869
rect 3969 18864 18755 18866
rect 3969 18808 3974 18864
rect 4030 18808 18694 18864
rect 18750 18808 18755 18864
rect 3969 18806 18755 18808
rect 3969 18803 4035 18806
rect 18689 18803 18755 18806
rect 18137 18730 18203 18733
rect 3052 18728 18203 18730
rect 3052 18672 18142 18728
rect 18198 18672 18203 18728
rect 3052 18670 18203 18672
rect 0 18640 800 18670
rect 1669 18667 1735 18670
rect 18137 18667 18203 18670
rect 19885 18730 19951 18733
rect 22000 18730 22800 18760
rect 19885 18728 22800 18730
rect 19885 18672 19890 18728
rect 19946 18672 22800 18728
rect 19885 18670 22800 18672
rect 19885 18667 19951 18670
rect 22000 18640 22800 18670
rect 3417 18594 3483 18597
rect 3969 18594 4035 18597
rect 3417 18592 4035 18594
rect 3417 18536 3422 18592
rect 3478 18536 3974 18592
rect 4030 18536 4035 18592
rect 3417 18534 4035 18536
rect 3417 18531 3483 18534
rect 3969 18531 4035 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 2405 18458 2471 18461
rect 2865 18458 2931 18461
rect 2405 18456 2931 18458
rect 2405 18400 2410 18456
rect 2466 18400 2870 18456
rect 2926 18400 2931 18456
rect 2405 18398 2931 18400
rect 2405 18395 2471 18398
rect 2865 18395 2931 18398
rect 0 18322 800 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 800 18262
rect 1945 18259 2011 18262
rect 3693 18322 3759 18325
rect 17125 18322 17191 18325
rect 3693 18320 17191 18322
rect 3693 18264 3698 18320
rect 3754 18264 17130 18320
rect 17186 18264 17191 18320
rect 3693 18262 17191 18264
rect 3693 18259 3759 18262
rect 17125 18259 17191 18262
rect 21081 18322 21147 18325
rect 22000 18322 22800 18352
rect 21081 18320 22800 18322
rect 21081 18264 21086 18320
rect 21142 18264 22800 18320
rect 21081 18262 22800 18264
rect 21081 18259 21147 18262
rect 22000 18232 22800 18262
rect 1301 18186 1367 18189
rect 3693 18186 3759 18189
rect 9121 18186 9187 18189
rect 1301 18184 3759 18186
rect 1301 18128 1306 18184
rect 1362 18128 3698 18184
rect 3754 18128 3759 18184
rect 1301 18126 3759 18128
rect 1301 18123 1367 18126
rect 3693 18123 3759 18126
rect 7652 18184 9187 18186
rect 7652 18128 9126 18184
rect 9182 18128 9187 18184
rect 7652 18126 9187 18128
rect 3601 18050 3667 18053
rect 4337 18050 4403 18053
rect 3601 18048 4403 18050
rect 3601 17992 3606 18048
rect 3662 17992 4342 18048
rect 4398 17992 4403 18048
rect 3601 17990 4403 17992
rect 3601 17987 3667 17990
rect 4337 17987 4403 17990
rect 4705 18050 4771 18053
rect 7652 18050 7712 18126
rect 9121 18123 9187 18126
rect 4705 18048 7712 18050
rect 4705 17992 4710 18048
rect 4766 17992 7712 18048
rect 4705 17990 7712 17992
rect 11697 18050 11763 18053
rect 12893 18050 12959 18053
rect 11697 18048 12959 18050
rect 11697 17992 11702 18048
rect 11758 17992 12898 18048
rect 12954 17992 12959 18048
rect 11697 17990 12959 17992
rect 4705 17987 4771 17990
rect 11697 17987 11763 17990
rect 12893 17987 12959 17990
rect 7808 17984 8128 17985
rect 0 17914 800 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 3601 17914 3667 17917
rect 0 17912 3667 17914
rect 0 17856 3606 17912
rect 3662 17856 3667 17912
rect 0 17854 3667 17856
rect 0 17824 800 17854
rect 3601 17851 3667 17854
rect 8477 17916 8543 17917
rect 8477 17912 8524 17916
rect 8588 17914 8594 17916
rect 9673 17914 9739 17917
rect 12341 17914 12407 17917
rect 8477 17856 8482 17912
rect 8477 17852 8524 17856
rect 8588 17854 8634 17914
rect 9673 17912 12407 17914
rect 9673 17856 9678 17912
rect 9734 17856 12346 17912
rect 12402 17856 12407 17912
rect 9673 17854 12407 17856
rect 8588 17852 8594 17854
rect 8477 17851 8543 17852
rect 9673 17851 9739 17854
rect 12341 17851 12407 17854
rect 20253 17914 20319 17917
rect 22000 17914 22800 17944
rect 20253 17912 22800 17914
rect 20253 17856 20258 17912
rect 20314 17856 22800 17912
rect 20253 17854 22800 17856
rect 20253 17851 20319 17854
rect 22000 17824 22800 17854
rect 4061 17778 4127 17781
rect 12249 17778 12315 17781
rect 4061 17776 12315 17778
rect 4061 17720 4066 17776
rect 4122 17720 12254 17776
rect 12310 17720 12315 17776
rect 4061 17718 12315 17720
rect 4061 17715 4127 17718
rect 12249 17715 12315 17718
rect 4521 17642 4587 17645
rect 5349 17642 5415 17645
rect 4521 17640 5415 17642
rect 4521 17584 4526 17640
rect 4582 17584 5354 17640
rect 5410 17584 5415 17640
rect 4521 17582 5415 17584
rect 4521 17579 4587 17582
rect 5349 17579 5415 17582
rect 5993 17642 6059 17645
rect 8334 17642 8340 17644
rect 5993 17640 8340 17642
rect 5993 17584 5998 17640
rect 6054 17584 8340 17640
rect 5993 17582 8340 17584
rect 5993 17579 6059 17582
rect 8334 17580 8340 17582
rect 8404 17580 8410 17644
rect 8569 17642 8635 17645
rect 9070 17642 9076 17644
rect 8569 17640 9076 17642
rect 8569 17584 8574 17640
rect 8630 17584 9076 17640
rect 8569 17582 9076 17584
rect 8569 17579 8635 17582
rect 9070 17580 9076 17582
rect 9140 17642 9146 17644
rect 14549 17642 14615 17645
rect 9140 17640 14615 17642
rect 9140 17584 14554 17640
rect 14610 17584 14615 17640
rect 9140 17582 14615 17584
rect 9140 17580 9146 17582
rect 14549 17579 14615 17582
rect 0 17506 800 17536
rect 1945 17506 2011 17509
rect 0 17504 2011 17506
rect 0 17448 1950 17504
rect 2006 17448 2011 17504
rect 0 17446 2011 17448
rect 0 17416 800 17446
rect 1945 17443 2011 17446
rect 21173 17506 21239 17509
rect 22000 17506 22800 17536
rect 21173 17504 22800 17506
rect 21173 17448 21178 17504
rect 21234 17448 22800 17504
rect 21173 17446 22800 17448
rect 21173 17443 21239 17446
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 22000 17416 22800 17446
rect 18104 17375 18424 17376
rect 3325 17234 3391 17237
rect 4889 17234 4955 17237
rect 3325 17232 4955 17234
rect 3325 17176 3330 17232
rect 3386 17176 4894 17232
rect 4950 17176 4955 17232
rect 3325 17174 4955 17176
rect 3325 17171 3391 17174
rect 4889 17171 4955 17174
rect 9806 17172 9812 17236
rect 9876 17234 9882 17236
rect 12525 17234 12591 17237
rect 17493 17234 17559 17237
rect 9876 17232 17559 17234
rect 9876 17176 12530 17232
rect 12586 17176 17498 17232
rect 17554 17176 17559 17232
rect 9876 17174 17559 17176
rect 9876 17172 9882 17174
rect 12525 17171 12591 17174
rect 17493 17171 17559 17174
rect 0 17098 800 17128
rect 1577 17098 1643 17101
rect 0 17096 1643 17098
rect 0 17040 1582 17096
rect 1638 17040 1643 17096
rect 0 17038 1643 17040
rect 0 17008 800 17038
rect 1577 17035 1643 17038
rect 6637 17098 6703 17101
rect 8753 17100 8819 17101
rect 7598 17098 7604 17100
rect 6637 17096 7604 17098
rect 6637 17040 6642 17096
rect 6698 17040 7604 17096
rect 6637 17038 7604 17040
rect 6637 17035 6703 17038
rect 7598 17036 7604 17038
rect 7668 17036 7674 17100
rect 8702 17098 8708 17100
rect 8662 17038 8708 17098
rect 8772 17096 8819 17100
rect 8814 17040 8819 17096
rect 8702 17036 8708 17038
rect 8772 17036 8819 17040
rect 8753 17035 8819 17036
rect 11421 17098 11487 17101
rect 12985 17098 13051 17101
rect 11421 17096 13051 17098
rect 11421 17040 11426 17096
rect 11482 17040 12990 17096
rect 13046 17040 13051 17096
rect 11421 17038 13051 17040
rect 11421 17035 11487 17038
rect 12985 17035 13051 17038
rect 20345 17098 20411 17101
rect 22000 17098 22800 17128
rect 20345 17096 22800 17098
rect 20345 17040 20350 17096
rect 20406 17040 22800 17096
rect 20345 17038 22800 17040
rect 20345 17035 20411 17038
rect 22000 17008 22800 17038
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 11329 16826 11395 16829
rect 12709 16826 12775 16829
rect 11329 16824 12775 16826
rect 11329 16768 11334 16824
rect 11390 16768 12714 16824
rect 12770 16768 12775 16824
rect 11329 16766 12775 16768
rect 11329 16763 11395 16766
rect 12709 16763 12775 16766
rect 0 16690 800 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 800 16630
rect 1577 16627 1643 16630
rect 8753 16690 8819 16693
rect 15285 16690 15351 16693
rect 8753 16688 15351 16690
rect 8753 16632 8758 16688
rect 8814 16632 15290 16688
rect 15346 16632 15351 16688
rect 8753 16630 15351 16632
rect 8753 16627 8819 16630
rect 15285 16627 15351 16630
rect 21081 16690 21147 16693
rect 22000 16690 22800 16720
rect 21081 16688 22800 16690
rect 21081 16632 21086 16688
rect 21142 16632 22800 16688
rect 21081 16630 22800 16632
rect 21081 16627 21147 16630
rect 22000 16600 22800 16630
rect 1393 16554 1459 16557
rect 8886 16554 8892 16556
rect 1393 16552 8892 16554
rect 1393 16496 1398 16552
rect 1454 16496 8892 16552
rect 1393 16494 8892 16496
rect 1393 16491 1459 16494
rect 8886 16492 8892 16494
rect 8956 16554 8962 16556
rect 9121 16554 9187 16557
rect 8956 16552 9187 16554
rect 8956 16496 9126 16552
rect 9182 16496 9187 16552
rect 8956 16494 9187 16496
rect 8956 16492 8962 16494
rect 9121 16491 9187 16494
rect 11605 16554 11671 16557
rect 12249 16554 12315 16557
rect 11605 16552 12315 16554
rect 11605 16496 11610 16552
rect 11666 16496 12254 16552
rect 12310 16496 12315 16552
rect 11605 16494 12315 16496
rect 11605 16491 11671 16494
rect 12249 16491 12315 16494
rect 6361 16418 6427 16421
rect 8753 16418 8819 16421
rect 6361 16416 8819 16418
rect 6361 16360 6366 16416
rect 6422 16360 8758 16416
rect 8814 16360 8819 16416
rect 6361 16358 8819 16360
rect 6361 16355 6427 16358
rect 8753 16355 8819 16358
rect 4376 16352 4696 16353
rect 0 16282 800 16312
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 1945 16282 2011 16285
rect 0 16280 2011 16282
rect 0 16224 1950 16280
rect 2006 16224 2011 16280
rect 0 16222 2011 16224
rect 0 16192 800 16222
rect 1945 16219 2011 16222
rect 20713 16282 20779 16285
rect 22000 16282 22800 16312
rect 20713 16280 22800 16282
rect 20713 16224 20718 16280
rect 20774 16224 22800 16280
rect 20713 16222 22800 16224
rect 20713 16219 20779 16222
rect 22000 16192 22800 16222
rect 10961 16146 11027 16149
rect 13997 16146 14063 16149
rect 10961 16144 14063 16146
rect 10961 16088 10966 16144
rect 11022 16088 14002 16144
rect 14058 16088 14063 16144
rect 10961 16086 14063 16088
rect 10961 16083 11027 16086
rect 13997 16083 14063 16086
rect 0 15874 800 15904
rect 2865 15874 2931 15877
rect 0 15872 2931 15874
rect 0 15816 2870 15872
rect 2926 15816 2931 15872
rect 0 15814 2931 15816
rect 0 15784 800 15814
rect 2865 15811 2931 15814
rect 4889 15874 4955 15877
rect 5206 15874 5212 15876
rect 4889 15872 5212 15874
rect 4889 15816 4894 15872
rect 4950 15816 5212 15872
rect 4889 15814 5212 15816
rect 4889 15811 4955 15814
rect 5206 15812 5212 15814
rect 5276 15812 5282 15876
rect 20253 15874 20319 15877
rect 22000 15874 22800 15904
rect 20253 15872 22800 15874
rect 20253 15816 20258 15872
rect 20314 15816 22800 15872
rect 20253 15814 22800 15816
rect 20253 15811 20319 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 22000 15784 22800 15814
rect 14672 15743 14992 15744
rect 12801 15602 12867 15605
rect 12934 15602 12940 15604
rect 12801 15600 12940 15602
rect 12801 15544 12806 15600
rect 12862 15544 12940 15600
rect 12801 15542 12940 15544
rect 12801 15539 12867 15542
rect 12934 15540 12940 15542
rect 13004 15540 13010 15604
rect 0 15466 800 15496
rect 1577 15466 1643 15469
rect 0 15464 1643 15466
rect 0 15408 1582 15464
rect 1638 15408 1643 15464
rect 0 15406 1643 15408
rect 0 15376 800 15406
rect 1577 15403 1643 15406
rect 2221 15466 2287 15469
rect 5809 15466 5875 15469
rect 7925 15466 7991 15469
rect 2221 15464 7991 15466
rect 2221 15408 2226 15464
rect 2282 15408 5814 15464
rect 5870 15408 7930 15464
rect 7986 15408 7991 15464
rect 2221 15406 7991 15408
rect 2221 15403 2287 15406
rect 5809 15403 5875 15406
rect 7925 15403 7991 15406
rect 8477 15466 8543 15469
rect 11789 15468 11855 15469
rect 8477 15464 11714 15466
rect 8477 15408 8482 15464
rect 8538 15408 11714 15464
rect 8477 15406 11714 15408
rect 8477 15403 8543 15406
rect 8845 15330 8911 15333
rect 9581 15330 9647 15333
rect 8845 15328 9647 15330
rect 8845 15272 8850 15328
rect 8906 15272 9586 15328
rect 9642 15272 9647 15328
rect 8845 15270 9647 15272
rect 8845 15267 8911 15270
rect 9581 15267 9647 15270
rect 4376 15264 4696 15265
rect 0 15194 800 15224
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 2773 15194 2839 15197
rect 0 15192 2839 15194
rect 0 15136 2778 15192
rect 2834 15136 2839 15192
rect 0 15134 2839 15136
rect 0 15104 800 15134
rect 2773 15131 2839 15134
rect 4797 15196 4863 15197
rect 4797 15192 4844 15196
rect 4908 15194 4914 15196
rect 5349 15194 5415 15197
rect 9397 15194 9463 15197
rect 4797 15136 4802 15192
rect 4797 15132 4844 15136
rect 4908 15134 4954 15194
rect 5349 15192 9463 15194
rect 5349 15136 5354 15192
rect 5410 15136 9402 15192
rect 9458 15136 9463 15192
rect 5349 15134 9463 15136
rect 11654 15194 11714 15406
rect 11789 15464 11836 15468
rect 11900 15466 11906 15468
rect 19701 15466 19767 15469
rect 22000 15466 22800 15496
rect 11789 15408 11794 15464
rect 11789 15404 11836 15408
rect 11900 15406 11946 15466
rect 19701 15464 22800 15466
rect 19701 15408 19706 15464
rect 19762 15408 22800 15464
rect 19701 15406 22800 15408
rect 11900 15404 11906 15406
rect 11789 15403 11855 15404
rect 19701 15403 19767 15406
rect 22000 15376 22800 15406
rect 13629 15332 13695 15333
rect 13629 15328 13676 15332
rect 13740 15330 13746 15332
rect 13629 15272 13634 15328
rect 13629 15268 13676 15272
rect 13740 15270 13786 15330
rect 13740 15268 13746 15270
rect 13629 15267 13695 15268
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 15142 15194 15148 15196
rect 11654 15134 15148 15194
rect 4908 15132 4914 15134
rect 4797 15131 4863 15132
rect 5349 15131 5415 15134
rect 9397 15131 9463 15134
rect 15142 15132 15148 15134
rect 15212 15194 15218 15196
rect 17677 15194 17743 15197
rect 15212 15192 17743 15194
rect 15212 15136 17682 15192
rect 17738 15136 17743 15192
rect 15212 15134 17743 15136
rect 15212 15132 15218 15134
rect 17677 15131 17743 15134
rect 20621 15194 20687 15197
rect 22000 15194 22800 15224
rect 20621 15192 22800 15194
rect 20621 15136 20626 15192
rect 20682 15136 22800 15192
rect 20621 15134 22800 15136
rect 20621 15131 20687 15134
rect 22000 15104 22800 15134
rect 3785 15058 3851 15061
rect 12065 15058 12131 15061
rect 3785 15056 12131 15058
rect 3785 15000 3790 15056
rect 3846 15000 12070 15056
rect 12126 15000 12131 15056
rect 3785 14998 12131 15000
rect 3785 14995 3851 14998
rect 12065 14995 12131 14998
rect 15285 15058 15351 15061
rect 18873 15058 18939 15061
rect 15285 15056 18939 15058
rect 15285 15000 15290 15056
rect 15346 15000 18878 15056
rect 18934 15000 18939 15056
rect 15285 14998 18939 15000
rect 15285 14995 15351 14998
rect 18873 14995 18939 14998
rect 11697 14922 11763 14925
rect 7652 14920 11763 14922
rect 7652 14864 11702 14920
rect 11758 14864 11763 14920
rect 7652 14862 11763 14864
rect 0 14786 800 14816
rect 2313 14786 2379 14789
rect 0 14784 2379 14786
rect 0 14728 2318 14784
rect 2374 14728 2379 14784
rect 0 14726 2379 14728
rect 0 14696 800 14726
rect 2313 14723 2379 14726
rect 7046 14724 7052 14788
rect 7116 14786 7122 14788
rect 7281 14786 7347 14789
rect 7652 14786 7712 14862
rect 11697 14859 11763 14862
rect 12617 14922 12683 14925
rect 18413 14922 18479 14925
rect 12617 14920 18479 14922
rect 12617 14864 12622 14920
rect 12678 14864 18418 14920
rect 18474 14864 18479 14920
rect 12617 14862 18479 14864
rect 12617 14859 12683 14862
rect 18413 14859 18479 14862
rect 8385 14788 8451 14789
rect 7116 14784 7712 14786
rect 7116 14728 7286 14784
rect 7342 14728 7712 14784
rect 7116 14726 7712 14728
rect 7116 14724 7122 14726
rect 7281 14723 7347 14726
rect 8334 14724 8340 14788
rect 8404 14786 8451 14788
rect 11145 14786 11211 14789
rect 12014 14786 12020 14788
rect 8404 14784 8496 14786
rect 8446 14728 8496 14784
rect 8404 14726 8496 14728
rect 9814 14784 12020 14786
rect 9814 14728 11150 14784
rect 11206 14728 12020 14784
rect 9814 14726 12020 14728
rect 8404 14724 8451 14726
rect 8385 14723 8451 14724
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 8477 14650 8543 14653
rect 9622 14650 9628 14652
rect 8477 14648 9628 14650
rect 8477 14592 8482 14648
rect 8538 14592 9628 14648
rect 8477 14590 9628 14592
rect 8477 14587 8543 14590
rect 9622 14588 9628 14590
rect 9692 14588 9698 14652
rect 5625 14514 5691 14517
rect 9814 14514 9874 14726
rect 11145 14723 11211 14726
rect 12014 14724 12020 14726
rect 12084 14724 12090 14788
rect 19701 14786 19767 14789
rect 22000 14786 22800 14816
rect 19701 14784 22800 14786
rect 19701 14728 19706 14784
rect 19762 14728 22800 14784
rect 19701 14726 22800 14728
rect 19701 14723 19767 14726
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 22000 14696 22800 14726
rect 14672 14655 14992 14656
rect 9949 14650 10015 14653
rect 11973 14650 12039 14653
rect 9949 14648 12039 14650
rect 9949 14592 9954 14648
rect 10010 14592 11978 14648
rect 12034 14592 12039 14648
rect 9949 14590 12039 14592
rect 9949 14587 10015 14590
rect 11973 14587 12039 14590
rect 5625 14512 9874 14514
rect 5625 14456 5630 14512
rect 5686 14456 9874 14512
rect 5625 14454 9874 14456
rect 5625 14451 5691 14454
rect 0 14378 800 14408
rect 1945 14378 2011 14381
rect 0 14376 2011 14378
rect 0 14320 1950 14376
rect 2006 14320 2011 14376
rect 0 14318 2011 14320
rect 0 14288 800 14318
rect 1945 14315 2011 14318
rect 6729 14378 6795 14381
rect 17401 14378 17467 14381
rect 6729 14376 17467 14378
rect 6729 14320 6734 14376
rect 6790 14320 17406 14376
rect 17462 14320 17467 14376
rect 6729 14318 17467 14320
rect 6729 14315 6795 14318
rect 17401 14315 17467 14318
rect 20437 14378 20503 14381
rect 22000 14378 22800 14408
rect 20437 14376 22800 14378
rect 20437 14320 20442 14376
rect 20498 14320 22800 14376
rect 20437 14318 22800 14320
rect 20437 14315 20503 14318
rect 22000 14288 22800 14318
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 0 13970 800 14000
rect 1761 13970 1827 13973
rect 0 13968 1827 13970
rect 0 13912 1766 13968
rect 1822 13912 1827 13968
rect 0 13910 1827 13912
rect 0 13880 800 13910
rect 1761 13907 1827 13910
rect 11237 13970 11303 13973
rect 12065 13970 12131 13973
rect 11237 13968 12131 13970
rect 11237 13912 11242 13968
rect 11298 13912 12070 13968
rect 12126 13912 12131 13968
rect 11237 13910 12131 13912
rect 11237 13907 11303 13910
rect 12065 13907 12131 13910
rect 12801 13970 12867 13973
rect 18873 13970 18939 13973
rect 12801 13968 18939 13970
rect 12801 13912 12806 13968
rect 12862 13912 18878 13968
rect 18934 13912 18939 13968
rect 12801 13910 18939 13912
rect 12801 13907 12867 13910
rect 18873 13907 18939 13910
rect 19977 13970 20043 13973
rect 20110 13970 20116 13972
rect 19977 13968 20116 13970
rect 19977 13912 19982 13968
rect 20038 13912 20116 13968
rect 19977 13910 20116 13912
rect 19977 13907 20043 13910
rect 20110 13908 20116 13910
rect 20180 13908 20186 13972
rect 20345 13970 20411 13973
rect 22000 13970 22800 14000
rect 20345 13968 22800 13970
rect 20345 13912 20350 13968
rect 20406 13912 22800 13968
rect 20345 13910 22800 13912
rect 20345 13907 20411 13910
rect 22000 13880 22800 13910
rect 10225 13834 10291 13837
rect 10358 13834 10364 13836
rect 10225 13832 10364 13834
rect 10225 13776 10230 13832
rect 10286 13776 10364 13832
rect 10225 13774 10364 13776
rect 10225 13771 10291 13774
rect 10358 13772 10364 13774
rect 10428 13834 10434 13836
rect 12893 13834 12959 13837
rect 10428 13832 12959 13834
rect 10428 13776 12898 13832
rect 12954 13776 12959 13832
rect 10428 13774 12959 13776
rect 10428 13772 10434 13774
rect 12893 13771 12959 13774
rect 15101 13834 15167 13837
rect 16021 13834 16087 13837
rect 15101 13832 16087 13834
rect 15101 13776 15106 13832
rect 15162 13776 16026 13832
rect 16082 13776 16087 13832
rect 15101 13774 16087 13776
rect 15101 13771 15167 13774
rect 16021 13771 16087 13774
rect 18321 13834 18387 13837
rect 20621 13834 20687 13837
rect 18321 13832 20687 13834
rect 18321 13776 18326 13832
rect 18382 13776 20626 13832
rect 20682 13776 20687 13832
rect 18321 13774 20687 13776
rect 18321 13771 18387 13774
rect 20621 13771 20687 13774
rect 11053 13698 11119 13701
rect 12157 13698 12223 13701
rect 11053 13696 12223 13698
rect 11053 13640 11058 13696
rect 11114 13640 12162 13696
rect 12218 13640 12223 13696
rect 11053 13638 12223 13640
rect 11053 13635 11119 13638
rect 12157 13635 12223 13638
rect 7808 13632 8128 13633
rect 0 13562 800 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 2773 13562 2839 13565
rect 0 13560 2839 13562
rect 0 13504 2778 13560
rect 2834 13504 2839 13560
rect 0 13502 2839 13504
rect 0 13472 800 13502
rect 2773 13499 2839 13502
rect 11646 13500 11652 13564
rect 11716 13562 11722 13564
rect 14365 13562 14431 13565
rect 11716 13560 14431 13562
rect 11716 13504 14370 13560
rect 14426 13504 14431 13560
rect 11716 13502 14431 13504
rect 11716 13500 11722 13502
rect 14365 13499 14431 13502
rect 21081 13562 21147 13565
rect 22000 13562 22800 13592
rect 21081 13560 22800 13562
rect 21081 13504 21086 13560
rect 21142 13504 22800 13560
rect 21081 13502 22800 13504
rect 21081 13499 21147 13502
rect 22000 13472 22800 13502
rect 2405 13426 2471 13429
rect 10225 13426 10291 13429
rect 2405 13424 10291 13426
rect 2405 13368 2410 13424
rect 2466 13368 10230 13424
rect 10286 13368 10291 13424
rect 2405 13366 10291 13368
rect 2405 13363 2471 13366
rect 10225 13363 10291 13366
rect 10409 13426 10475 13429
rect 15653 13426 15719 13429
rect 10409 13424 15719 13426
rect 10409 13368 10414 13424
rect 10470 13368 15658 13424
rect 15714 13368 15719 13424
rect 10409 13366 15719 13368
rect 10409 13363 10475 13366
rect 15653 13363 15719 13366
rect 6913 13290 6979 13293
rect 9305 13290 9371 13293
rect 6913 13288 9371 13290
rect 6913 13232 6918 13288
rect 6974 13232 9310 13288
rect 9366 13232 9371 13288
rect 6913 13230 9371 13232
rect 6913 13227 6979 13230
rect 9305 13227 9371 13230
rect 10685 13290 10751 13293
rect 16757 13290 16823 13293
rect 10685 13288 16823 13290
rect 10685 13232 10690 13288
rect 10746 13232 16762 13288
rect 16818 13232 16823 13288
rect 10685 13230 16823 13232
rect 10685 13227 10751 13230
rect 16757 13227 16823 13230
rect 0 13154 800 13184
rect 1761 13154 1827 13157
rect 0 13152 1827 13154
rect 0 13096 1766 13152
rect 1822 13096 1827 13152
rect 0 13094 1827 13096
rect 0 13064 800 13094
rect 1761 13091 1827 13094
rect 8109 13154 8175 13157
rect 9213 13154 9279 13157
rect 8109 13152 9279 13154
rect 8109 13096 8114 13152
rect 8170 13096 9218 13152
rect 9274 13096 9279 13152
rect 8109 13094 9279 13096
rect 8109 13091 8175 13094
rect 9213 13091 9279 13094
rect 12893 13154 12959 13157
rect 17033 13154 17099 13157
rect 12893 13152 17099 13154
rect 12893 13096 12898 13152
rect 12954 13096 17038 13152
rect 17094 13096 17099 13152
rect 12893 13094 17099 13096
rect 12893 13091 12959 13094
rect 17033 13091 17099 13094
rect 20529 13154 20595 13157
rect 22000 13154 22800 13184
rect 20529 13152 22800 13154
rect 20529 13096 20534 13152
rect 20590 13096 22800 13152
rect 20529 13094 22800 13096
rect 20529 13091 20595 13094
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 22000 13064 22800 13094
rect 18104 13023 18424 13024
rect 1577 12882 1643 12885
rect 12341 12882 12407 12885
rect 13445 12882 13511 12885
rect 1577 12880 8448 12882
rect 1577 12824 1582 12880
rect 1638 12824 8448 12880
rect 1577 12822 8448 12824
rect 1577 12819 1643 12822
rect 0 12746 800 12776
rect 8388 12749 8448 12822
rect 9124 12880 13511 12882
rect 9124 12824 12346 12880
rect 12402 12824 13450 12880
rect 13506 12824 13511 12880
rect 9124 12822 13511 12824
rect 1669 12746 1735 12749
rect 0 12744 1735 12746
rect 0 12688 1674 12744
rect 1730 12688 1735 12744
rect 0 12686 1735 12688
rect 0 12656 800 12686
rect 1669 12683 1735 12686
rect 8385 12746 8451 12749
rect 8661 12746 8727 12749
rect 8385 12744 8727 12746
rect 8385 12688 8390 12744
rect 8446 12688 8666 12744
rect 8722 12688 8727 12744
rect 8385 12686 8727 12688
rect 8385 12683 8451 12686
rect 8661 12683 8727 12686
rect 6862 12548 6868 12612
rect 6932 12610 6938 12612
rect 7005 12610 7071 12613
rect 9124 12610 9184 12822
rect 12341 12819 12407 12822
rect 13445 12819 13511 12822
rect 14273 12882 14339 12885
rect 15929 12882 15995 12885
rect 14273 12880 15995 12882
rect 14273 12824 14278 12880
rect 14334 12824 15934 12880
rect 15990 12824 15995 12880
rect 14273 12822 15995 12824
rect 14273 12819 14339 12822
rect 15929 12819 15995 12822
rect 10593 12746 10659 12749
rect 16849 12746 16915 12749
rect 10593 12744 16915 12746
rect 10593 12688 10598 12744
rect 10654 12688 16854 12744
rect 16910 12688 16915 12744
rect 10593 12686 16915 12688
rect 10593 12683 10659 12686
rect 16849 12683 16915 12686
rect 20253 12746 20319 12749
rect 22000 12746 22800 12776
rect 20253 12744 22800 12746
rect 20253 12688 20258 12744
rect 20314 12688 22800 12744
rect 20253 12686 22800 12688
rect 20253 12683 20319 12686
rect 22000 12656 22800 12686
rect 6932 12608 7071 12610
rect 6932 12552 7010 12608
rect 7066 12552 7071 12608
rect 6932 12550 7071 12552
rect 6932 12548 6938 12550
rect 7005 12547 7071 12550
rect 8480 12550 9184 12610
rect 9305 12610 9371 12613
rect 10174 12610 10180 12612
rect 9305 12608 10180 12610
rect 9305 12552 9310 12608
rect 9366 12552 10180 12608
rect 9305 12550 10180 12552
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 8480 12477 8540 12550
rect 9305 12547 9371 12550
rect 10174 12548 10180 12550
rect 10244 12548 10250 12612
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 6177 12474 6243 12477
rect 6177 12472 6608 12474
rect 6177 12416 6182 12472
rect 6238 12416 6608 12472
rect 6177 12414 6608 12416
rect 6177 12411 6243 12414
rect 0 12338 800 12368
rect 6548 12341 6608 12414
rect 8477 12472 8543 12477
rect 8477 12416 8482 12472
rect 8538 12416 8543 12472
rect 8477 12411 8543 12416
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 6545 12336 6611 12341
rect 6545 12280 6550 12336
rect 6606 12280 6611 12336
rect 6545 12275 6611 12280
rect 9673 12338 9739 12341
rect 10869 12338 10935 12341
rect 9673 12336 10935 12338
rect 9673 12280 9678 12336
rect 9734 12280 10874 12336
rect 10930 12280 10935 12336
rect 9673 12278 10935 12280
rect 9673 12275 9739 12278
rect 10869 12275 10935 12278
rect 12198 12276 12204 12340
rect 12268 12338 12274 12340
rect 17217 12338 17283 12341
rect 12268 12336 17283 12338
rect 12268 12280 17222 12336
rect 17278 12280 17283 12336
rect 12268 12278 17283 12280
rect 12268 12276 12274 12278
rect 7414 12140 7420 12204
rect 7484 12202 7490 12204
rect 7649 12202 7715 12205
rect 12206 12202 12266 12276
rect 17217 12275 17283 12278
rect 21173 12338 21239 12341
rect 22000 12338 22800 12368
rect 21173 12336 22800 12338
rect 21173 12280 21178 12336
rect 21234 12280 22800 12336
rect 21173 12278 22800 12280
rect 21173 12275 21239 12278
rect 22000 12248 22800 12278
rect 7484 12200 7715 12202
rect 7484 12144 7654 12200
rect 7710 12144 7715 12200
rect 7484 12142 7715 12144
rect 7484 12140 7490 12142
rect 7649 12139 7715 12142
rect 10734 12142 12266 12202
rect 6862 12004 6868 12068
rect 6932 12066 6938 12068
rect 7649 12066 7715 12069
rect 10225 12068 10291 12069
rect 6932 12064 7715 12066
rect 6932 12008 7654 12064
rect 7710 12008 7715 12064
rect 6932 12006 7715 12008
rect 6932 12004 6938 12006
rect 7649 12003 7715 12006
rect 10174 12004 10180 12068
rect 10244 12066 10291 12068
rect 10244 12064 10336 12066
rect 10286 12008 10336 12064
rect 10244 12006 10336 12008
rect 10244 12004 10291 12006
rect 10225 12003 10291 12004
rect 4376 12000 4696 12001
rect 0 11930 800 11960
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 1669 11930 1735 11933
rect 0 11928 1735 11930
rect 0 11872 1674 11928
rect 1730 11872 1735 11928
rect 0 11870 1735 11872
rect 0 11840 800 11870
rect 1669 11867 1735 11870
rect 6729 11930 6795 11933
rect 10734 11930 10794 12142
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 6729 11928 10794 11930
rect 6729 11872 6734 11928
rect 6790 11872 10794 11928
rect 6729 11870 10794 11872
rect 20621 11930 20687 11933
rect 22000 11930 22800 11960
rect 20621 11928 22800 11930
rect 20621 11872 20626 11928
rect 20682 11872 22800 11928
rect 20621 11870 22800 11872
rect 6729 11867 6795 11870
rect 20621 11867 20687 11870
rect 22000 11840 22800 11870
rect 5022 11732 5028 11796
rect 5092 11794 5098 11796
rect 7097 11794 7163 11797
rect 5092 11792 7163 11794
rect 5092 11736 7102 11792
rect 7158 11736 7163 11792
rect 5092 11734 7163 11736
rect 5092 11732 5098 11734
rect 7097 11731 7163 11734
rect 10685 11794 10751 11797
rect 11145 11794 11211 11797
rect 10685 11792 11211 11794
rect 10685 11736 10690 11792
rect 10746 11736 11150 11792
rect 11206 11736 11211 11792
rect 10685 11734 11211 11736
rect 10685 11731 10751 11734
rect 11145 11731 11211 11734
rect 0 11658 800 11688
rect 3049 11658 3115 11661
rect 0 11656 3115 11658
rect 0 11600 3054 11656
rect 3110 11600 3115 11656
rect 0 11598 3115 11600
rect 0 11568 800 11598
rect 3049 11595 3115 11598
rect 4613 11658 4679 11661
rect 4981 11660 5047 11661
rect 4838 11658 4844 11660
rect 4613 11656 4844 11658
rect 4613 11600 4618 11656
rect 4674 11600 4844 11656
rect 4613 11598 4844 11600
rect 4613 11595 4679 11598
rect 4838 11596 4844 11598
rect 4908 11596 4914 11660
rect 4981 11656 5028 11660
rect 5092 11658 5098 11660
rect 12157 11658 12223 11661
rect 5092 11656 12223 11658
rect 4981 11600 4986 11656
rect 5092 11600 12162 11656
rect 12218 11600 12223 11656
rect 4981 11596 5028 11600
rect 5092 11598 12223 11600
rect 5092 11596 5098 11598
rect 4981 11595 5047 11596
rect 12157 11595 12223 11598
rect 21173 11658 21239 11661
rect 22000 11658 22800 11688
rect 21173 11656 22800 11658
rect 21173 11600 21178 11656
rect 21234 11600 22800 11656
rect 21173 11598 22800 11600
rect 21173 11595 21239 11598
rect 22000 11568 22800 11598
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 12382 11324 12388 11388
rect 12452 11386 12458 11388
rect 12709 11386 12775 11389
rect 12452 11384 12775 11386
rect 12452 11328 12714 11384
rect 12770 11328 12775 11384
rect 12452 11326 12775 11328
rect 12452 11324 12458 11326
rect 12709 11323 12775 11326
rect 0 11250 800 11280
rect 2865 11250 2931 11253
rect 0 11248 2931 11250
rect 0 11192 2870 11248
rect 2926 11192 2931 11248
rect 0 11190 2931 11192
rect 0 11160 800 11190
rect 2865 11187 2931 11190
rect 6821 11250 6887 11253
rect 9489 11250 9555 11253
rect 9765 11252 9831 11253
rect 9765 11250 9812 11252
rect 6821 11248 9555 11250
rect 6821 11192 6826 11248
rect 6882 11192 9494 11248
rect 9550 11192 9555 11248
rect 6821 11190 9555 11192
rect 9720 11248 9812 11250
rect 9720 11192 9770 11248
rect 9720 11190 9812 11192
rect 6821 11187 6887 11190
rect 9489 11187 9555 11190
rect 9765 11188 9812 11190
rect 9876 11188 9882 11252
rect 11973 11250 12039 11253
rect 12157 11250 12223 11253
rect 16757 11250 16823 11253
rect 18505 11250 18571 11253
rect 11973 11248 16823 11250
rect 11973 11192 11978 11248
rect 12034 11192 12162 11248
rect 12218 11192 16762 11248
rect 16818 11192 16823 11248
rect 11973 11190 16823 11192
rect 9765 11187 9831 11188
rect 11973 11187 12039 11190
rect 12157 11187 12223 11190
rect 16757 11187 16823 11190
rect 18462 11248 18571 11250
rect 18462 11192 18510 11248
rect 18566 11192 18571 11248
rect 18462 11187 18571 11192
rect 21081 11250 21147 11253
rect 22000 11250 22800 11280
rect 21081 11248 22800 11250
rect 21081 11192 21086 11248
rect 21142 11192 22800 11248
rect 21081 11190 22800 11192
rect 21081 11187 21147 11190
rect 1393 11114 1459 11117
rect 1393 11112 7666 11114
rect 1393 11056 1398 11112
rect 1454 11056 7666 11112
rect 1393 11054 7666 11056
rect 1393 11051 1459 11054
rect 7606 10978 7666 11054
rect 9438 11052 9444 11116
rect 9508 11114 9514 11116
rect 17309 11114 17375 11117
rect 9508 11112 17375 11114
rect 9508 11056 17314 11112
rect 17370 11056 17375 11112
rect 9508 11054 17375 11056
rect 18462 11114 18522 11187
rect 22000 11160 22800 11190
rect 19517 11114 19583 11117
rect 18462 11112 19583 11114
rect 18462 11056 19522 11112
rect 19578 11056 19583 11112
rect 18462 11054 19583 11056
rect 9508 11052 9514 11054
rect 17309 11051 17375 11054
rect 19517 11051 19583 11054
rect 9213 10978 9279 10981
rect 7606 10976 9279 10978
rect 7606 10920 9218 10976
rect 9274 10920 9279 10976
rect 7606 10918 9279 10920
rect 9213 10915 9279 10918
rect 12433 10978 12499 10981
rect 17309 10978 17375 10981
rect 12433 10976 17375 10978
rect 12433 10920 12438 10976
rect 12494 10920 17314 10976
rect 17370 10920 17375 10976
rect 12433 10918 17375 10920
rect 12433 10915 12499 10918
rect 17309 10915 17375 10918
rect 4376 10912 4696 10913
rect 0 10842 800 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3785 10842 3851 10845
rect 4061 10842 4127 10845
rect 0 10840 3851 10842
rect 0 10784 3790 10840
rect 3846 10784 3851 10840
rect 0 10782 3851 10784
rect 0 10752 800 10782
rect 3785 10779 3851 10782
rect 3926 10840 4127 10842
rect 3926 10784 4066 10840
rect 4122 10784 4127 10840
rect 3926 10782 4127 10784
rect 3785 10706 3851 10709
rect 3926 10706 3986 10782
rect 4061 10779 4127 10782
rect 7598 10780 7604 10844
rect 7668 10842 7674 10844
rect 8569 10842 8635 10845
rect 22000 10842 22800 10872
rect 7668 10840 8635 10842
rect 7668 10784 8574 10840
rect 8630 10784 8635 10840
rect 7668 10782 8635 10784
rect 7668 10780 7674 10782
rect 8569 10779 8635 10782
rect 18600 10782 22800 10842
rect 3785 10704 3986 10706
rect 3785 10648 3790 10704
rect 3846 10648 3986 10704
rect 3785 10646 3986 10648
rect 5257 10706 5323 10709
rect 8518 10706 8524 10708
rect 5257 10704 8524 10706
rect 5257 10648 5262 10704
rect 5318 10648 8524 10704
rect 5257 10646 8524 10648
rect 3785 10643 3851 10646
rect 5257 10643 5323 10646
rect 8518 10644 8524 10646
rect 8588 10644 8594 10708
rect 13721 10706 13787 10709
rect 14089 10706 14155 10709
rect 13721 10704 14155 10706
rect 13721 10648 13726 10704
rect 13782 10648 14094 10704
rect 14150 10648 14155 10704
rect 13721 10646 14155 10648
rect 13721 10643 13787 10646
rect 14089 10643 14155 10646
rect 14457 10706 14523 10709
rect 18600 10706 18660 10782
rect 22000 10752 22800 10782
rect 14457 10704 18660 10706
rect 14457 10648 14462 10704
rect 14518 10648 18660 10704
rect 14457 10646 18660 10648
rect 14457 10643 14523 10646
rect 3417 10570 3483 10573
rect 4429 10570 4495 10573
rect 8293 10570 8359 10573
rect 3417 10568 4495 10570
rect 3417 10512 3422 10568
rect 3478 10512 4434 10568
rect 4490 10512 4495 10568
rect 3417 10510 4495 10512
rect 3417 10507 3483 10510
rect 4429 10507 4495 10510
rect 4846 10568 8359 10570
rect 4846 10512 8298 10568
rect 8354 10512 8359 10568
rect 4846 10510 8359 10512
rect 0 10434 800 10464
rect 4846 10434 4906 10510
rect 8293 10507 8359 10510
rect 8661 10570 8727 10573
rect 9397 10570 9463 10573
rect 15101 10570 15167 10573
rect 8661 10568 15167 10570
rect 8661 10512 8666 10568
rect 8722 10512 9402 10568
rect 9458 10512 15106 10568
rect 15162 10512 15167 10568
rect 8661 10510 15167 10512
rect 8661 10507 8727 10510
rect 9397 10507 9463 10510
rect 15101 10507 15167 10510
rect 18229 10570 18295 10573
rect 18638 10570 18644 10572
rect 18229 10568 18644 10570
rect 18229 10512 18234 10568
rect 18290 10512 18644 10568
rect 18229 10510 18644 10512
rect 18229 10507 18295 10510
rect 18638 10508 18644 10510
rect 18708 10508 18714 10572
rect 0 10374 4906 10434
rect 8661 10434 8727 10437
rect 8886 10434 8892 10436
rect 8661 10432 8892 10434
rect 8661 10376 8666 10432
rect 8722 10376 8892 10432
rect 8661 10374 8892 10376
rect 0 10344 800 10374
rect 8661 10371 8727 10374
rect 8886 10372 8892 10374
rect 8956 10372 8962 10436
rect 10133 10434 10199 10437
rect 13997 10436 14063 10437
rect 10358 10434 10364 10436
rect 10133 10432 10364 10434
rect 10133 10376 10138 10432
rect 10194 10376 10364 10432
rect 10133 10374 10364 10376
rect 10133 10371 10199 10374
rect 10358 10372 10364 10374
rect 10428 10372 10434 10436
rect 13997 10434 14044 10436
rect 13952 10432 14044 10434
rect 13952 10376 14002 10432
rect 13952 10374 14044 10376
rect 13997 10372 14044 10374
rect 14108 10372 14114 10436
rect 16665 10434 16731 10437
rect 22000 10434 22800 10464
rect 16665 10432 22800 10434
rect 16665 10376 16670 10432
rect 16726 10376 22800 10432
rect 16665 10374 22800 10376
rect 13997 10371 14063 10372
rect 16665 10371 16731 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22000 10344 22800 10374
rect 14672 10303 14992 10304
rect 5165 10300 5231 10301
rect 5165 10296 5212 10300
rect 5276 10298 5282 10300
rect 5165 10240 5170 10296
rect 5165 10236 5212 10240
rect 5276 10238 5322 10298
rect 5276 10236 5282 10238
rect 5165 10235 5231 10236
rect 5625 10162 5691 10165
rect 14733 10162 14799 10165
rect 5625 10160 14799 10162
rect 5625 10104 5630 10160
rect 5686 10104 14738 10160
rect 14794 10104 14799 10160
rect 5625 10102 14799 10104
rect 5625 10099 5691 10102
rect 14733 10099 14799 10102
rect 20110 10100 20116 10164
rect 20180 10162 20186 10164
rect 20345 10162 20411 10165
rect 20180 10160 20411 10162
rect 20180 10104 20350 10160
rect 20406 10104 20411 10160
rect 20180 10102 20411 10104
rect 20180 10100 20186 10102
rect 20345 10099 20411 10102
rect 0 10026 800 10056
rect 4061 10026 4127 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 800 9966
rect 4061 9963 4127 9966
rect 7465 10026 7531 10029
rect 8201 10026 8267 10029
rect 7465 10024 8267 10026
rect 7465 9968 7470 10024
rect 7526 9968 8206 10024
rect 8262 9968 8267 10024
rect 7465 9966 8267 9968
rect 7465 9963 7531 9966
rect 8201 9963 8267 9966
rect 8569 10026 8635 10029
rect 13721 10028 13787 10029
rect 8569 10024 11714 10026
rect 8569 9968 8574 10024
rect 8630 9968 11714 10024
rect 8569 9966 11714 9968
rect 8569 9963 8635 9966
rect 4981 9890 5047 9893
rect 7465 9890 7531 9893
rect 4981 9888 7531 9890
rect 4981 9832 4986 9888
rect 5042 9832 7470 9888
rect 7526 9832 7531 9888
rect 4981 9830 7531 9832
rect 11654 9890 11714 9966
rect 13670 9964 13676 10028
rect 13740 10026 13787 10028
rect 14089 10026 14155 10029
rect 22000 10026 22800 10056
rect 13740 10024 13832 10026
rect 13782 9968 13832 10024
rect 13740 9966 13832 9968
rect 14089 10024 22800 10026
rect 14089 9968 14094 10024
rect 14150 9968 22800 10024
rect 14089 9966 22800 9968
rect 13740 9964 13787 9966
rect 13721 9963 13787 9964
rect 14089 9963 14155 9966
rect 22000 9936 22800 9966
rect 14457 9890 14523 9893
rect 17401 9890 17467 9893
rect 11654 9888 17467 9890
rect 11654 9832 14462 9888
rect 14518 9832 17406 9888
rect 17462 9832 17467 9888
rect 11654 9830 17467 9832
rect 4981 9827 5047 9830
rect 7465 9827 7531 9830
rect 14457 9827 14523 9830
rect 17401 9827 17467 9830
rect 17542 9830 17970 9890
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 12525 9754 12591 9757
rect 15285 9754 15351 9757
rect 12525 9752 15351 9754
rect 12525 9696 12530 9752
rect 12586 9696 15290 9752
rect 15346 9696 15351 9752
rect 12525 9694 15351 9696
rect 12525 9691 12591 9694
rect 15285 9691 15351 9694
rect 16849 9754 16915 9757
rect 17542 9754 17602 9830
rect 17910 9754 17970 9830
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 16849 9752 17602 9754
rect 16849 9696 16854 9752
rect 16910 9696 17602 9752
rect 16849 9694 17602 9696
rect 17772 9694 17970 9754
rect 16849 9691 16915 9694
rect 0 9618 800 9648
rect 17772 9621 17832 9694
rect 8293 9618 8359 9621
rect 0 9616 8359 9618
rect 0 9560 8298 9616
rect 8354 9560 8359 9616
rect 0 9558 8359 9560
rect 0 9528 800 9558
rect 8293 9555 8359 9558
rect 10961 9618 11027 9621
rect 11646 9618 11652 9620
rect 10961 9616 11652 9618
rect 10961 9560 10966 9616
rect 11022 9560 11652 9616
rect 10961 9558 11652 9560
rect 10961 9555 11027 9558
rect 11646 9556 11652 9558
rect 11716 9556 11722 9620
rect 12934 9556 12940 9620
rect 13004 9618 13010 9620
rect 13077 9618 13143 9621
rect 13004 9616 13143 9618
rect 13004 9560 13082 9616
rect 13138 9560 13143 9616
rect 13004 9558 13143 9560
rect 13004 9556 13010 9558
rect 13077 9555 13143 9558
rect 13629 9618 13695 9621
rect 14365 9618 14431 9621
rect 16941 9618 17007 9621
rect 13629 9616 13922 9618
rect 13629 9560 13634 9616
rect 13690 9560 13922 9616
rect 13629 9558 13922 9560
rect 13629 9555 13695 9558
rect 2773 9482 2839 9485
rect 1350 9480 2839 9482
rect 1350 9424 2778 9480
rect 2834 9424 2839 9480
rect 1350 9422 2839 9424
rect 0 9210 800 9240
rect 1350 9210 1410 9422
rect 2773 9419 2839 9422
rect 5073 9482 5139 9485
rect 8937 9482 9003 9485
rect 13670 9482 13676 9484
rect 5073 9480 8402 9482
rect 5073 9424 5078 9480
rect 5134 9424 8402 9480
rect 5073 9422 8402 9424
rect 5073 9419 5139 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 0 9150 1410 9210
rect 7097 9210 7163 9213
rect 7230 9210 7236 9212
rect 7097 9208 7236 9210
rect 7097 9152 7102 9208
rect 7158 9152 7236 9208
rect 7097 9150 7236 9152
rect 0 9120 800 9150
rect 7097 9147 7163 9150
rect 7230 9148 7236 9150
rect 7300 9148 7306 9212
rect 8342 9074 8402 9422
rect 8937 9480 13676 9482
rect 8937 9424 8942 9480
rect 8998 9424 13676 9480
rect 8937 9422 13676 9424
rect 8937 9419 9003 9422
rect 13670 9420 13676 9422
rect 13740 9420 13746 9484
rect 13862 9482 13922 9558
rect 14365 9616 17007 9618
rect 14365 9560 14370 9616
rect 14426 9560 16946 9616
rect 17002 9560 17007 9616
rect 14365 9558 17007 9560
rect 14365 9555 14431 9558
rect 16941 9555 17007 9558
rect 17769 9616 17835 9621
rect 22000 9618 22800 9648
rect 17769 9560 17774 9616
rect 17830 9560 17835 9616
rect 17769 9555 17835 9560
rect 19934 9558 22800 9618
rect 14917 9482 14983 9485
rect 13862 9480 14983 9482
rect 13862 9424 14922 9480
rect 14978 9424 14983 9480
rect 13862 9422 14983 9424
rect 14917 9419 14983 9422
rect 15837 9482 15903 9485
rect 19934 9482 19994 9558
rect 22000 9528 22800 9558
rect 15837 9480 19994 9482
rect 15837 9424 15842 9480
rect 15898 9424 19994 9480
rect 15837 9422 19994 9424
rect 15837 9419 15903 9422
rect 9213 9346 9279 9349
rect 14365 9346 14431 9349
rect 9213 9344 14431 9346
rect 9213 9288 9218 9344
rect 9274 9288 14370 9344
rect 14426 9288 14431 9344
rect 9213 9286 14431 9288
rect 9213 9283 9279 9286
rect 14365 9283 14431 9286
rect 16389 9346 16455 9349
rect 18781 9346 18847 9349
rect 16389 9344 18847 9346
rect 16389 9288 16394 9344
rect 16450 9288 18786 9344
rect 18842 9288 18847 9344
rect 16389 9286 18847 9288
rect 16389 9283 16455 9286
rect 18781 9283 18847 9286
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 8569 9210 8635 9213
rect 8702 9210 8708 9212
rect 8569 9208 8708 9210
rect 8569 9152 8574 9208
rect 8630 9152 8708 9208
rect 8569 9150 8708 9152
rect 8569 9147 8635 9150
rect 8702 9148 8708 9150
rect 8772 9210 8778 9212
rect 11697 9210 11763 9213
rect 11881 9212 11947 9213
rect 8772 9208 11763 9210
rect 8772 9152 11702 9208
rect 11758 9152 11763 9208
rect 8772 9150 11763 9152
rect 8772 9148 8778 9150
rect 11697 9147 11763 9150
rect 11830 9148 11836 9212
rect 11900 9210 11947 9212
rect 22000 9210 22800 9240
rect 11900 9208 11992 9210
rect 11942 9152 11992 9208
rect 11900 9150 11992 9152
rect 15472 9150 22800 9210
rect 11900 9148 11947 9150
rect 11881 9147 11947 9148
rect 15472 9077 15532 9150
rect 22000 9120 22800 9150
rect 15193 9074 15259 9077
rect 8342 9072 15259 9074
rect 8342 9016 15198 9072
rect 15254 9016 15259 9072
rect 8342 9014 15259 9016
rect 15193 9011 15259 9014
rect 15469 9072 15535 9077
rect 15469 9016 15474 9072
rect 15530 9016 15535 9072
rect 15469 9011 15535 9016
rect 17309 9074 17375 9077
rect 19517 9074 19583 9077
rect 17309 9072 19583 9074
rect 17309 9016 17314 9072
rect 17370 9016 19522 9072
rect 19578 9016 19583 9072
rect 17309 9014 19583 9016
rect 17309 9011 17375 9014
rect 19517 9011 19583 9014
rect 7465 8938 7531 8941
rect 9622 8938 9628 8940
rect 7465 8936 9628 8938
rect 7465 8880 7470 8936
rect 7526 8880 9628 8936
rect 7465 8878 9628 8880
rect 7465 8875 7531 8878
rect 9622 8876 9628 8878
rect 9692 8938 9698 8940
rect 15745 8938 15811 8941
rect 9692 8936 15811 8938
rect 9692 8880 15750 8936
rect 15806 8880 15811 8936
rect 9692 8878 15811 8880
rect 9692 8876 9698 8878
rect 15745 8875 15811 8878
rect 0 8802 800 8832
rect 1301 8802 1367 8805
rect 6177 8802 6243 8805
rect 6453 8802 6519 8805
rect 6821 8802 6887 8805
rect 10501 8804 10567 8805
rect 9070 8802 9076 8804
rect 0 8800 4170 8802
rect 0 8744 1306 8800
rect 1362 8744 4170 8800
rect 0 8742 4170 8744
rect 0 8712 800 8742
rect 1301 8739 1367 8742
rect 4110 8530 4170 8742
rect 6177 8800 6746 8802
rect 6177 8744 6182 8800
rect 6238 8744 6458 8800
rect 6514 8744 6746 8800
rect 6177 8742 6746 8744
rect 6177 8739 6243 8742
rect 6453 8739 6519 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 6686 8666 6746 8742
rect 6821 8800 9076 8802
rect 6821 8744 6826 8800
rect 6882 8744 9076 8800
rect 6821 8742 9076 8744
rect 6821 8739 6887 8742
rect 9070 8740 9076 8742
rect 9140 8802 9146 8804
rect 10174 8802 10180 8804
rect 9140 8742 10180 8802
rect 9140 8740 9146 8742
rect 10174 8740 10180 8742
rect 10244 8740 10250 8804
rect 10501 8800 10548 8804
rect 10612 8802 10618 8804
rect 10501 8744 10506 8800
rect 10501 8740 10548 8744
rect 10612 8742 10658 8802
rect 10612 8740 10618 8742
rect 12014 8740 12020 8804
rect 12084 8802 12090 8804
rect 12157 8802 12223 8805
rect 12084 8800 12223 8802
rect 12084 8744 12162 8800
rect 12218 8744 12223 8800
rect 12084 8742 12223 8744
rect 12084 8740 12090 8742
rect 10501 8739 10567 8740
rect 12157 8739 12223 8742
rect 12801 8802 12867 8805
rect 16757 8802 16823 8805
rect 12801 8800 16823 8802
rect 12801 8744 12806 8800
rect 12862 8744 16762 8800
rect 16818 8744 16823 8800
rect 12801 8742 16823 8744
rect 12801 8739 12867 8742
rect 16757 8739 16823 8742
rect 18597 8802 18663 8805
rect 22000 8802 22800 8832
rect 18597 8800 22800 8802
rect 18597 8744 18602 8800
rect 18658 8744 22800 8800
rect 18597 8742 22800 8744
rect 18597 8739 18663 8742
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 22000 8712 22800 8742
rect 18104 8671 18424 8672
rect 8293 8666 8359 8669
rect 6686 8664 8359 8666
rect 6686 8608 8298 8664
rect 8354 8608 8359 8664
rect 6686 8606 8359 8608
rect 8293 8603 8359 8606
rect 9765 8666 9831 8669
rect 11053 8666 11119 8669
rect 9765 8664 11119 8666
rect 9765 8608 9770 8664
rect 9826 8608 11058 8664
rect 11114 8608 11119 8664
rect 9765 8606 11119 8608
rect 9765 8603 9831 8606
rect 11053 8603 11119 8606
rect 11973 8666 12039 8669
rect 13813 8666 13879 8669
rect 11973 8664 13879 8666
rect 11973 8608 11978 8664
rect 12034 8608 13818 8664
rect 13874 8608 13879 8664
rect 11973 8606 13879 8608
rect 11973 8603 12039 8606
rect 13813 8603 13879 8606
rect 14089 8666 14155 8669
rect 15101 8666 15167 8669
rect 14089 8664 15167 8666
rect 14089 8608 14094 8664
rect 14150 8608 15106 8664
rect 15162 8608 15167 8664
rect 14089 8606 15167 8608
rect 14089 8603 14155 8606
rect 15101 8603 15167 8606
rect 18597 8666 18663 8669
rect 20437 8666 20503 8669
rect 18597 8664 20503 8666
rect 18597 8608 18602 8664
rect 18658 8608 20442 8664
rect 20498 8608 20503 8664
rect 18597 8606 20503 8608
rect 18597 8603 18663 8606
rect 20437 8603 20503 8606
rect 6453 8530 6519 8533
rect 19885 8530 19951 8533
rect 4110 8528 19951 8530
rect 4110 8472 6458 8528
rect 6514 8472 19890 8528
rect 19946 8472 19951 8528
rect 4110 8470 19951 8472
rect 6453 8467 6519 8470
rect 19885 8467 19951 8470
rect 0 8394 800 8424
rect 3417 8394 3483 8397
rect 0 8392 3483 8394
rect 0 8336 3422 8392
rect 3478 8336 3483 8392
rect 0 8334 3483 8336
rect 0 8304 800 8334
rect 3417 8331 3483 8334
rect 4613 8394 4679 8397
rect 5073 8394 5139 8397
rect 4613 8392 5139 8394
rect 4613 8336 4618 8392
rect 4674 8336 5078 8392
rect 5134 8336 5139 8392
rect 4613 8334 5139 8336
rect 4613 8331 4679 8334
rect 5073 8331 5139 8334
rect 6269 8394 6335 8397
rect 8109 8394 8175 8397
rect 6269 8392 8175 8394
rect 6269 8336 6274 8392
rect 6330 8336 8114 8392
rect 8170 8336 8175 8392
rect 6269 8334 8175 8336
rect 6269 8331 6335 8334
rect 8109 8331 8175 8334
rect 8293 8394 8359 8397
rect 16573 8394 16639 8397
rect 8293 8392 16639 8394
rect 8293 8336 8298 8392
rect 8354 8336 16578 8392
rect 16634 8336 16639 8392
rect 8293 8334 16639 8336
rect 8293 8331 8359 8334
rect 16573 8331 16639 8334
rect 16757 8394 16823 8397
rect 22000 8394 22800 8424
rect 16757 8392 22800 8394
rect 16757 8336 16762 8392
rect 16818 8336 22800 8392
rect 16757 8334 22800 8336
rect 16757 8331 16823 8334
rect 22000 8304 22800 8334
rect 10225 8258 10291 8261
rect 10593 8258 10659 8261
rect 14457 8258 14523 8261
rect 10225 8256 14523 8258
rect 10225 8200 10230 8256
rect 10286 8200 10598 8256
rect 10654 8200 14462 8256
rect 14518 8200 14523 8256
rect 10225 8198 14523 8200
rect 10225 8195 10291 8198
rect 10593 8195 10659 8198
rect 14457 8195 14523 8198
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 9397 8122 9463 8125
rect 12198 8122 12204 8124
rect 9397 8120 12204 8122
rect 9397 8064 9402 8120
rect 9458 8064 12204 8120
rect 9397 8062 12204 8064
rect 9397 8059 9463 8062
rect 12198 8060 12204 8062
rect 12268 8060 12274 8124
rect 0 7986 800 8016
rect 7557 7986 7623 7989
rect 10041 7986 10107 7989
rect 16757 7986 16823 7989
rect 0 7926 4906 7986
rect 0 7896 800 7926
rect 4846 7850 4906 7926
rect 7557 7984 16823 7986
rect 7557 7928 7562 7984
rect 7618 7928 10046 7984
rect 10102 7928 16762 7984
rect 16818 7928 16823 7984
rect 7557 7926 16823 7928
rect 7557 7923 7623 7926
rect 10041 7923 10107 7926
rect 16757 7923 16823 7926
rect 19149 7986 19215 7989
rect 22000 7986 22800 8016
rect 19149 7984 22800 7986
rect 19149 7928 19154 7984
rect 19210 7928 22800 7984
rect 19149 7926 22800 7928
rect 19149 7923 19215 7926
rect 22000 7896 22800 7926
rect 15142 7850 15148 7852
rect 4846 7790 15148 7850
rect 15142 7788 15148 7790
rect 15212 7788 15218 7852
rect 17861 7850 17927 7853
rect 18689 7850 18755 7853
rect 17861 7848 18755 7850
rect 17861 7792 17866 7848
rect 17922 7792 18694 7848
rect 18750 7792 18755 7848
rect 17861 7790 18755 7792
rect 17861 7787 17927 7790
rect 18689 7787 18755 7790
rect 0 7714 800 7744
rect 4061 7714 4127 7717
rect 0 7712 4127 7714
rect 0 7656 4066 7712
rect 4122 7656 4127 7712
rect 0 7654 4127 7656
rect 0 7624 800 7654
rect 4061 7651 4127 7654
rect 7230 7652 7236 7716
rect 7300 7714 7306 7716
rect 7925 7714 7991 7717
rect 11094 7714 11100 7716
rect 7300 7712 11100 7714
rect 7300 7656 7930 7712
rect 7986 7656 11100 7712
rect 7300 7654 11100 7656
rect 7300 7652 7306 7654
rect 7925 7651 7991 7654
rect 11094 7652 11100 7654
rect 11164 7652 11170 7716
rect 12341 7714 12407 7717
rect 17309 7714 17375 7717
rect 12341 7712 17375 7714
rect 12341 7656 12346 7712
rect 12402 7656 17314 7712
rect 17370 7656 17375 7712
rect 12341 7654 17375 7656
rect 12341 7651 12407 7654
rect 17309 7651 17375 7654
rect 18597 7714 18663 7717
rect 22000 7714 22800 7744
rect 18597 7712 22800 7714
rect 18597 7656 18602 7712
rect 18658 7656 22800 7712
rect 18597 7654 22800 7656
rect 18597 7651 18663 7654
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 22000 7624 22800 7654
rect 18104 7583 18424 7584
rect 6269 7578 6335 7581
rect 9765 7578 9831 7581
rect 6269 7576 9831 7578
rect 6269 7520 6274 7576
rect 6330 7520 9770 7576
rect 9826 7520 9831 7576
rect 6269 7518 9831 7520
rect 6269 7515 6335 7518
rect 9765 7515 9831 7518
rect 10542 7516 10548 7580
rect 10612 7578 10618 7580
rect 10685 7578 10751 7581
rect 10612 7576 10751 7578
rect 10612 7520 10690 7576
rect 10746 7520 10751 7576
rect 10612 7518 10751 7520
rect 10612 7516 10618 7518
rect 10685 7515 10751 7518
rect 3417 7442 3483 7445
rect 5533 7442 5599 7445
rect 3417 7440 5599 7442
rect 3417 7384 3422 7440
rect 3478 7384 5538 7440
rect 5594 7384 5599 7440
rect 3417 7382 5599 7384
rect 3417 7379 3483 7382
rect 5533 7379 5599 7382
rect 5809 7442 5875 7445
rect 15837 7442 15903 7445
rect 5809 7440 15903 7442
rect 5809 7384 5814 7440
rect 5870 7384 15842 7440
rect 15898 7384 15903 7440
rect 5809 7382 15903 7384
rect 5809 7379 5875 7382
rect 15837 7379 15903 7382
rect 0 7306 800 7336
rect 4061 7306 4127 7309
rect 0 7304 4127 7306
rect 0 7248 4066 7304
rect 4122 7248 4127 7304
rect 0 7246 4127 7248
rect 0 7216 800 7246
rect 4061 7243 4127 7246
rect 6545 7306 6611 7309
rect 8937 7306 9003 7309
rect 9438 7306 9444 7308
rect 6545 7304 8402 7306
rect 6545 7248 6550 7304
rect 6606 7248 8402 7304
rect 6545 7246 8402 7248
rect 6545 7243 6611 7246
rect 2681 7170 2747 7173
rect 3785 7170 3851 7173
rect 2681 7168 3851 7170
rect 2681 7112 2686 7168
rect 2742 7112 3790 7168
rect 3846 7112 3851 7168
rect 2681 7110 3851 7112
rect 8342 7170 8402 7246
rect 8937 7304 9444 7306
rect 8937 7248 8942 7304
rect 8998 7248 9444 7304
rect 8937 7246 9444 7248
rect 8937 7243 9003 7246
rect 9438 7244 9444 7246
rect 9508 7244 9514 7308
rect 9806 7244 9812 7308
rect 9876 7306 9882 7308
rect 10501 7306 10567 7309
rect 9876 7304 10567 7306
rect 9876 7248 10506 7304
rect 10562 7248 10567 7304
rect 9876 7246 10567 7248
rect 9876 7244 9882 7246
rect 10501 7243 10567 7246
rect 12341 7306 12407 7309
rect 13905 7306 13971 7309
rect 12341 7304 13971 7306
rect 12341 7248 12346 7304
rect 12402 7248 13910 7304
rect 13966 7248 13971 7304
rect 12341 7246 13971 7248
rect 12341 7243 12407 7246
rect 13905 7243 13971 7246
rect 14038 7244 14044 7308
rect 14108 7306 14114 7308
rect 22000 7306 22800 7336
rect 14108 7246 22800 7306
rect 14108 7244 14114 7246
rect 13261 7170 13327 7173
rect 14046 7170 14106 7244
rect 22000 7216 22800 7246
rect 8342 7168 14106 7170
rect 8342 7112 13266 7168
rect 13322 7112 14106 7168
rect 8342 7110 14106 7112
rect 2681 7107 2747 7110
rect 3785 7107 3851 7110
rect 13261 7107 13327 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 8201 7034 8267 7037
rect 11881 7034 11947 7037
rect 8201 7032 11947 7034
rect 8201 6976 8206 7032
rect 8262 6976 11886 7032
rect 11942 6976 11947 7032
rect 8201 6974 11947 6976
rect 8201 6971 8267 6974
rect 11881 6971 11947 6974
rect 14089 7034 14155 7037
rect 14457 7034 14523 7037
rect 14089 7032 14523 7034
rect 14089 6976 14094 7032
rect 14150 6976 14462 7032
rect 14518 6976 14523 7032
rect 14089 6974 14523 6976
rect 14089 6971 14155 6974
rect 14457 6971 14523 6974
rect 16021 7034 16087 7037
rect 18822 7034 18828 7036
rect 16021 7032 18828 7034
rect 16021 6976 16026 7032
rect 16082 6976 18828 7032
rect 16021 6974 18828 6976
rect 16021 6971 16087 6974
rect 18822 6972 18828 6974
rect 18892 6972 18898 7036
rect 0 6898 800 6928
rect 7557 6898 7623 6901
rect 0 6896 7623 6898
rect 0 6840 7562 6896
rect 7618 6840 7623 6896
rect 0 6838 7623 6840
rect 0 6808 800 6838
rect 7557 6835 7623 6838
rect 8845 6898 8911 6901
rect 10133 6898 10199 6901
rect 12382 6898 12388 6900
rect 8845 6896 10199 6898
rect 8845 6840 8850 6896
rect 8906 6840 10138 6896
rect 10194 6840 10199 6896
rect 8845 6838 10199 6840
rect 8845 6835 8911 6838
rect 10133 6835 10199 6838
rect 10320 6838 12388 6898
rect 7925 6762 7991 6765
rect 10320 6762 10380 6838
rect 12382 6836 12388 6838
rect 12452 6836 12458 6900
rect 12617 6898 12683 6901
rect 12985 6898 13051 6901
rect 12617 6896 13051 6898
rect 12617 6840 12622 6896
rect 12678 6840 12990 6896
rect 13046 6840 13051 6896
rect 12617 6838 13051 6840
rect 12617 6835 12683 6838
rect 12985 6835 13051 6838
rect 13670 6836 13676 6900
rect 13740 6898 13746 6900
rect 22000 6898 22800 6928
rect 13740 6838 22800 6898
rect 13740 6836 13746 6838
rect 22000 6808 22800 6838
rect 12198 6762 12204 6764
rect 7925 6760 10380 6762
rect 7925 6704 7930 6760
rect 7986 6704 10380 6760
rect 7925 6702 10380 6704
rect 10550 6702 12204 6762
rect 7925 6699 7991 6702
rect 5073 6626 5139 6629
rect 10550 6626 10610 6702
rect 12198 6700 12204 6702
rect 12268 6700 12274 6764
rect 5073 6624 10610 6626
rect 5073 6568 5078 6624
rect 5134 6568 10610 6624
rect 5073 6566 10610 6568
rect 5073 6563 5139 6566
rect 4376 6560 4696 6561
rect 0 6490 800 6520
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 4061 6490 4127 6493
rect 0 6488 4127 6490
rect 0 6432 4066 6488
rect 4122 6432 4127 6488
rect 0 6430 4127 6432
rect 0 6400 800 6430
rect 4061 6427 4127 6430
rect 5993 6490 6059 6493
rect 7414 6490 7420 6492
rect 5993 6488 7420 6490
rect 5993 6432 5998 6488
rect 6054 6432 7420 6488
rect 5993 6430 7420 6432
rect 5993 6427 6059 6430
rect 7414 6428 7420 6430
rect 7484 6490 7490 6492
rect 11053 6490 11119 6493
rect 7484 6488 11119 6490
rect 7484 6432 11058 6488
rect 11114 6432 11119 6488
rect 7484 6430 11119 6432
rect 7484 6428 7490 6430
rect 11053 6427 11119 6430
rect 18638 6428 18644 6492
rect 18708 6490 18714 6492
rect 22000 6490 22800 6520
rect 18708 6430 22800 6490
rect 18708 6428 18714 6430
rect 22000 6400 22800 6430
rect 6729 6354 6795 6357
rect 11697 6354 11763 6357
rect 6729 6352 11763 6354
rect 6729 6296 6734 6352
rect 6790 6296 11702 6352
rect 11758 6296 11763 6352
rect 6729 6294 11763 6296
rect 6729 6291 6795 6294
rect 11697 6291 11763 6294
rect 12382 6292 12388 6356
rect 12452 6354 12458 6356
rect 20069 6354 20135 6357
rect 12452 6352 20135 6354
rect 12452 6296 20074 6352
rect 20130 6296 20135 6352
rect 12452 6294 20135 6296
rect 12452 6292 12458 6294
rect 20069 6291 20135 6294
rect 6729 6218 6795 6221
rect 11973 6218 12039 6221
rect 6729 6216 12039 6218
rect 6729 6160 6734 6216
rect 6790 6160 11978 6216
rect 12034 6160 12039 6216
rect 6729 6158 12039 6160
rect 6729 6155 6795 6158
rect 11973 6155 12039 6158
rect 12198 6156 12204 6220
rect 12268 6218 12274 6220
rect 15745 6218 15811 6221
rect 12268 6216 15811 6218
rect 12268 6160 15750 6216
rect 15806 6160 15811 6216
rect 12268 6158 15811 6160
rect 12268 6156 12274 6158
rect 15745 6155 15811 6158
rect 0 6082 800 6112
rect 4061 6082 4127 6085
rect 0 6080 4127 6082
rect 0 6024 4066 6080
rect 4122 6024 4127 6080
rect 0 6022 4127 6024
rect 0 5992 800 6022
rect 4061 6019 4127 6022
rect 4613 6082 4679 6085
rect 10225 6084 10291 6085
rect 4838 6082 4844 6084
rect 4613 6080 4844 6082
rect 4613 6024 4618 6080
rect 4674 6024 4844 6080
rect 4613 6022 4844 6024
rect 4613 6019 4679 6022
rect 4838 6020 4844 6022
rect 4908 6082 4914 6084
rect 7046 6082 7052 6084
rect 4908 6022 7052 6082
rect 4908 6020 4914 6022
rect 7046 6020 7052 6022
rect 7116 6020 7122 6084
rect 10174 6082 10180 6084
rect 10098 6022 10180 6082
rect 10244 6082 10291 6084
rect 12249 6082 12315 6085
rect 13813 6082 13879 6085
rect 22000 6082 22800 6112
rect 10244 6080 12315 6082
rect 10286 6024 12254 6080
rect 12310 6024 12315 6080
rect 10174 6020 10180 6022
rect 10244 6022 12315 6024
rect 10244 6020 10291 6022
rect 10225 6019 10291 6020
rect 12249 6019 12315 6022
rect 12574 6080 13879 6082
rect 12574 6024 13818 6080
rect 13874 6024 13879 6080
rect 12574 6022 13879 6024
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 4981 5946 5047 5949
rect 7189 5946 7255 5949
rect 4981 5944 7255 5946
rect 4981 5888 4986 5944
rect 5042 5888 7194 5944
rect 7250 5888 7255 5944
rect 4981 5886 7255 5888
rect 4981 5883 5047 5886
rect 7189 5883 7255 5886
rect 9673 5946 9739 5949
rect 11237 5946 11303 5949
rect 9673 5944 11303 5946
rect 9673 5888 9678 5944
rect 9734 5888 11242 5944
rect 11298 5888 11303 5944
rect 9673 5886 11303 5888
rect 9673 5883 9739 5886
rect 11237 5883 11303 5886
rect 11513 5946 11579 5949
rect 12574 5946 12634 6022
rect 13813 6019 13879 6022
rect 17174 6022 22800 6082
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 11513 5944 12634 5946
rect 11513 5888 11518 5944
rect 11574 5888 12634 5944
rect 11513 5886 12634 5888
rect 11513 5883 11579 5886
rect 6177 5810 6243 5813
rect 9121 5810 9187 5813
rect 15377 5810 15443 5813
rect 6177 5808 15443 5810
rect 6177 5752 6182 5808
rect 6238 5752 9126 5808
rect 9182 5752 15382 5808
rect 15438 5752 15443 5808
rect 6177 5750 15443 5752
rect 6177 5747 6243 5750
rect 9121 5747 9187 5750
rect 15377 5747 15443 5750
rect 0 5674 800 5704
rect 3969 5674 4035 5677
rect 0 5672 4035 5674
rect 0 5616 3974 5672
rect 4030 5616 4035 5672
rect 0 5614 4035 5616
rect 0 5584 800 5614
rect 3969 5611 4035 5614
rect 7741 5674 7807 5677
rect 17174 5674 17234 6022
rect 22000 5992 22800 6022
rect 7741 5672 17234 5674
rect 7741 5616 7746 5672
rect 7802 5616 17234 5672
rect 7741 5614 17234 5616
rect 17309 5674 17375 5677
rect 22000 5674 22800 5704
rect 17309 5672 22800 5674
rect 17309 5616 17314 5672
rect 17370 5616 22800 5672
rect 17309 5614 22800 5616
rect 7741 5611 7807 5614
rect 17309 5611 17375 5614
rect 22000 5584 22800 5614
rect 2681 5538 2747 5541
rect 4245 5538 4311 5541
rect 2681 5536 4311 5538
rect 2681 5480 2686 5536
rect 2742 5480 4250 5536
rect 4306 5480 4311 5536
rect 2681 5478 4311 5480
rect 2681 5475 2747 5478
rect 4245 5475 4311 5478
rect 12065 5538 12131 5541
rect 17953 5538 18019 5541
rect 12065 5536 18019 5538
rect 12065 5480 12070 5536
rect 12126 5480 17958 5536
rect 18014 5480 18019 5536
rect 12065 5478 18019 5480
rect 12065 5475 12131 5478
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 13077 5402 13143 5405
rect 13905 5402 13971 5405
rect 13077 5400 13971 5402
rect 13077 5344 13082 5400
rect 13138 5344 13910 5400
rect 13966 5344 13971 5400
rect 13077 5342 13971 5344
rect 13077 5339 13143 5342
rect 13905 5339 13971 5342
rect 0 5266 800 5296
rect 3509 5266 3575 5269
rect 0 5264 3575 5266
rect 0 5208 3514 5264
rect 3570 5208 3575 5264
rect 0 5206 3575 5208
rect 0 5176 800 5206
rect 3509 5203 3575 5206
rect 4245 5266 4311 5269
rect 5022 5266 5028 5268
rect 4245 5264 5028 5266
rect 4245 5208 4250 5264
rect 4306 5208 5028 5264
rect 4245 5206 5028 5208
rect 4245 5203 4311 5206
rect 5022 5204 5028 5206
rect 5092 5204 5098 5268
rect 7465 5266 7531 5269
rect 7649 5266 7715 5269
rect 8569 5268 8635 5269
rect 8518 5266 8524 5268
rect 7465 5264 7715 5266
rect 7465 5208 7470 5264
rect 7526 5208 7654 5264
rect 7710 5208 7715 5264
rect 7465 5206 7715 5208
rect 8442 5206 8524 5266
rect 8588 5266 8635 5268
rect 16113 5266 16179 5269
rect 8588 5264 16179 5266
rect 8630 5208 16118 5264
rect 16174 5208 16179 5264
rect 7465 5203 7531 5206
rect 7649 5203 7715 5206
rect 8518 5204 8524 5206
rect 8588 5206 16179 5208
rect 8588 5204 8635 5206
rect 8569 5203 8635 5204
rect 16113 5203 16179 5206
rect 17542 5133 17602 5478
rect 17953 5475 18019 5478
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 17953 5266 18019 5269
rect 22000 5266 22800 5296
rect 17953 5264 22800 5266
rect 17953 5208 17958 5264
rect 18014 5208 22800 5264
rect 17953 5206 22800 5208
rect 17953 5203 18019 5206
rect 22000 5176 22800 5206
rect 6545 5130 6611 5133
rect 13813 5130 13879 5133
rect 15653 5130 15719 5133
rect 6545 5128 15719 5130
rect 6545 5072 6550 5128
rect 6606 5072 13818 5128
rect 13874 5072 15658 5128
rect 15714 5072 15719 5128
rect 6545 5070 15719 5072
rect 17542 5128 17651 5133
rect 17542 5072 17590 5128
rect 17646 5072 17651 5128
rect 17542 5070 17651 5072
rect 6545 5067 6611 5070
rect 13813 5067 13879 5070
rect 15653 5067 15719 5070
rect 17585 5067 17651 5070
rect 18597 5130 18663 5133
rect 19241 5130 19307 5133
rect 18597 5128 19307 5130
rect 18597 5072 18602 5128
rect 18658 5072 19246 5128
rect 19302 5072 19307 5128
rect 18597 5070 19307 5072
rect 18597 5067 18663 5070
rect 19241 5067 19307 5070
rect 8293 4994 8359 4997
rect 11513 4994 11579 4997
rect 8293 4992 11579 4994
rect 8293 4936 8298 4992
rect 8354 4936 11518 4992
rect 11574 4936 11579 4992
rect 8293 4934 11579 4936
rect 8293 4931 8359 4934
rect 11513 4931 11579 4934
rect 12341 4994 12407 4997
rect 14089 4994 14155 4997
rect 12341 4992 14155 4994
rect 12341 4936 12346 4992
rect 12402 4936 14094 4992
rect 14150 4936 14155 4992
rect 12341 4934 14155 4936
rect 12341 4931 12407 4934
rect 14089 4931 14155 4934
rect 7808 4928 8128 4929
rect 0 4858 800 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 800 4798
rect 4061 4795 4127 4798
rect 5349 4858 5415 4861
rect 7281 4858 7347 4861
rect 5349 4856 7347 4858
rect 5349 4800 5354 4856
rect 5410 4800 7286 4856
rect 7342 4800 7347 4856
rect 5349 4798 7347 4800
rect 5349 4795 5415 4798
rect 7281 4795 7347 4798
rect 10685 4858 10751 4861
rect 14273 4858 14339 4861
rect 10685 4856 14339 4858
rect 10685 4800 10690 4856
rect 10746 4800 14278 4856
rect 14334 4800 14339 4856
rect 10685 4798 14339 4800
rect 10685 4795 10751 4798
rect 14273 4795 14339 4798
rect 15101 4858 15167 4861
rect 22000 4858 22800 4888
rect 15101 4856 22800 4858
rect 15101 4800 15106 4856
rect 15162 4800 22800 4856
rect 15101 4798 22800 4800
rect 15101 4795 15167 4798
rect 22000 4768 22800 4798
rect 6729 4722 6795 4725
rect 8477 4722 8543 4725
rect 6729 4720 8543 4722
rect 6729 4664 6734 4720
rect 6790 4664 8482 4720
rect 8538 4664 8543 4720
rect 6729 4662 8543 4664
rect 6729 4659 6795 4662
rect 8477 4659 8543 4662
rect 9949 4722 10015 4725
rect 16297 4722 16363 4725
rect 19425 4722 19491 4725
rect 9949 4720 19491 4722
rect 9949 4664 9954 4720
rect 10010 4664 16302 4720
rect 16358 4664 19430 4720
rect 19486 4664 19491 4720
rect 9949 4662 19491 4664
rect 9949 4659 10015 4662
rect 16297 4659 16363 4662
rect 19425 4659 19491 4662
rect 5809 4586 5875 4589
rect 8937 4586 9003 4589
rect 15653 4586 15719 4589
rect 18965 4586 19031 4589
rect 5809 4584 7068 4586
rect 5809 4528 5814 4584
rect 5870 4528 7068 4584
rect 5809 4526 7068 4528
rect 5809 4523 5875 4526
rect 0 4450 800 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 7008 4450 7068 4526
rect 8937 4584 15719 4586
rect 8937 4528 8942 4584
rect 8998 4528 15658 4584
rect 15714 4528 15719 4584
rect 8937 4526 15719 4528
rect 8937 4523 9003 4526
rect 15653 4523 15719 4526
rect 15840 4584 19031 4586
rect 15840 4528 18970 4584
rect 19026 4528 19031 4584
rect 15840 4526 19031 4528
rect 14825 4450 14891 4453
rect 15142 4450 15148 4452
rect 7008 4390 9506 4450
rect 0 4360 800 4390
rect 4061 4387 4127 4390
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 5901 4314 5967 4317
rect 8661 4314 8727 4317
rect 5901 4312 8727 4314
rect 5901 4256 5906 4312
rect 5962 4256 8666 4312
rect 8722 4256 8727 4312
rect 5901 4254 8727 4256
rect 5901 4251 5967 4254
rect 8661 4251 8727 4254
rect 4521 4178 4587 4181
rect 5809 4178 5875 4181
rect 4521 4176 5875 4178
rect 4521 4120 4526 4176
rect 4582 4120 5814 4176
rect 5870 4120 5875 4176
rect 4521 4118 5875 4120
rect 4521 4115 4587 4118
rect 5809 4115 5875 4118
rect 7649 4178 7715 4181
rect 8661 4178 8727 4181
rect 7649 4176 8727 4178
rect 7649 4120 7654 4176
rect 7710 4120 8666 4176
rect 8722 4120 8727 4176
rect 7649 4118 8727 4120
rect 9446 4178 9506 4390
rect 14825 4448 15148 4450
rect 14825 4392 14830 4448
rect 14886 4392 15148 4448
rect 14825 4390 15148 4392
rect 14825 4387 14891 4390
rect 15142 4388 15148 4390
rect 15212 4450 15218 4452
rect 15840 4450 15900 4526
rect 18965 4523 19031 4526
rect 15212 4390 15900 4450
rect 18965 4450 19031 4453
rect 22000 4450 22800 4480
rect 18965 4448 22800 4450
rect 18965 4392 18970 4448
rect 19026 4392 22800 4448
rect 18965 4390 22800 4392
rect 15212 4388 15218 4390
rect 18965 4387 19031 4390
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 22000 4360 22800 4390
rect 18104 4319 18424 4320
rect 15561 4178 15627 4181
rect 15837 4178 15903 4181
rect 9446 4176 15903 4178
rect 9446 4120 15566 4176
rect 15622 4120 15842 4176
rect 15898 4120 15903 4176
rect 9446 4118 15903 4120
rect 7649 4115 7715 4118
rect 8661 4115 8727 4118
rect 15561 4115 15627 4118
rect 15837 4115 15903 4118
rect 0 4042 800 4072
rect 13905 4042 13971 4045
rect 0 4040 13971 4042
rect 0 3984 13910 4040
rect 13966 3984 13971 4040
rect 0 3982 13971 3984
rect 0 3952 800 3982
rect 13905 3979 13971 3982
rect 17953 4042 18019 4045
rect 22000 4042 22800 4072
rect 17953 4040 22800 4042
rect 17953 3984 17958 4040
rect 18014 3984 22800 4040
rect 17953 3982 22800 3984
rect 17953 3979 18019 3982
rect 22000 3952 22800 3982
rect 5441 3906 5507 3909
rect 7005 3906 7071 3909
rect 5441 3904 7071 3906
rect 5441 3848 5446 3904
rect 5502 3848 7010 3904
rect 7066 3848 7071 3904
rect 5441 3846 7071 3848
rect 5441 3843 5507 3846
rect 7005 3843 7071 3846
rect 8661 3906 8727 3909
rect 10593 3906 10659 3909
rect 8661 3904 10659 3906
rect 8661 3848 8666 3904
rect 8722 3848 10598 3904
rect 10654 3848 10659 3904
rect 8661 3846 10659 3848
rect 8661 3843 8727 3846
rect 10593 3843 10659 3846
rect 7808 3840 8128 3841
rect 0 3770 800 3800
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 4981 3770 5047 3773
rect 5625 3770 5691 3773
rect 0 3710 4906 3770
rect 0 3680 800 3710
rect 4846 3634 4906 3710
rect 4981 3768 5691 3770
rect 4981 3712 4986 3768
rect 5042 3712 5630 3768
rect 5686 3712 5691 3768
rect 4981 3710 5691 3712
rect 4981 3707 5047 3710
rect 5625 3707 5691 3710
rect 8845 3770 8911 3773
rect 9581 3770 9647 3773
rect 8845 3768 9647 3770
rect 8845 3712 8850 3768
rect 8906 3712 9586 3768
rect 9642 3712 9647 3768
rect 8845 3710 9647 3712
rect 8845 3707 8911 3710
rect 9581 3707 9647 3710
rect 11094 3708 11100 3772
rect 11164 3770 11170 3772
rect 11697 3770 11763 3773
rect 11164 3768 11763 3770
rect 11164 3712 11702 3768
rect 11758 3712 11763 3768
rect 11164 3710 11763 3712
rect 11164 3708 11170 3710
rect 11697 3707 11763 3710
rect 15285 3770 15351 3773
rect 22000 3770 22800 3800
rect 15285 3768 22800 3770
rect 15285 3712 15290 3768
rect 15346 3712 22800 3768
rect 15285 3710 22800 3712
rect 15285 3707 15351 3710
rect 22000 3680 22800 3710
rect 13261 3634 13327 3637
rect 4846 3632 13327 3634
rect 4846 3576 13266 3632
rect 13322 3576 13327 3632
rect 4846 3574 13327 3576
rect 13261 3571 13327 3574
rect 8569 3498 8635 3501
rect 9622 3498 9628 3500
rect 8569 3496 9628 3498
rect 8569 3440 8574 3496
rect 8630 3440 9628 3496
rect 8569 3438 9628 3440
rect 8569 3435 8635 3438
rect 9622 3436 9628 3438
rect 9692 3498 9698 3500
rect 14273 3498 14339 3501
rect 9692 3496 14339 3498
rect 9692 3440 14278 3496
rect 14334 3440 14339 3496
rect 9692 3438 14339 3440
rect 9692 3436 9698 3438
rect 14273 3435 14339 3438
rect 0 3362 800 3392
rect 4061 3362 4127 3365
rect 0 3360 4127 3362
rect 0 3304 4066 3360
rect 4122 3304 4127 3360
rect 0 3302 4127 3304
rect 0 3272 800 3302
rect 4061 3299 4127 3302
rect 8201 3362 8267 3365
rect 8569 3362 8635 3365
rect 8201 3360 8635 3362
rect 8201 3304 8206 3360
rect 8262 3304 8574 3360
rect 8630 3304 8635 3360
rect 8201 3302 8635 3304
rect 8201 3299 8267 3302
rect 8569 3299 8635 3302
rect 18822 3300 18828 3364
rect 18892 3362 18898 3364
rect 22000 3362 22800 3392
rect 18892 3302 22800 3362
rect 18892 3300 18898 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 22000 3272 22800 3302
rect 18104 3231 18424 3232
rect 4838 3164 4844 3228
rect 4908 3226 4914 3228
rect 10593 3226 10659 3229
rect 4908 3224 10659 3226
rect 4908 3168 10598 3224
rect 10654 3168 10659 3224
rect 4908 3166 10659 3168
rect 4908 3164 4914 3166
rect 10593 3163 10659 3166
rect 3325 3090 3391 3093
rect 1350 3088 3391 3090
rect 1350 3032 3330 3088
rect 3386 3032 3391 3088
rect 1350 3030 3391 3032
rect 0 2954 800 2984
rect 1350 2954 1410 3030
rect 3325 3027 3391 3030
rect 7097 3090 7163 3093
rect 9397 3090 9463 3093
rect 11973 3090 12039 3093
rect 7097 3088 12039 3090
rect 7097 3032 7102 3088
rect 7158 3032 9402 3088
rect 9458 3032 11978 3088
rect 12034 3032 12039 3088
rect 7097 3030 12039 3032
rect 7097 3027 7163 3030
rect 9397 3027 9463 3030
rect 11973 3027 12039 3030
rect 0 2894 1410 2954
rect 2957 2954 3023 2957
rect 12985 2954 13051 2957
rect 18413 2954 18479 2957
rect 2957 2952 13051 2954
rect 2957 2896 2962 2952
rect 3018 2896 12990 2952
rect 13046 2896 13051 2952
rect 2957 2894 13051 2896
rect 0 2864 800 2894
rect 2957 2891 3023 2894
rect 8526 2821 8586 2894
rect 12985 2891 13051 2894
rect 13126 2952 18479 2954
rect 13126 2896 18418 2952
rect 18474 2896 18479 2952
rect 13126 2894 18479 2896
rect 8526 2816 8635 2821
rect 8526 2760 8574 2816
rect 8630 2760 8635 2816
rect 8526 2758 8635 2760
rect 8569 2755 8635 2758
rect 10593 2818 10659 2821
rect 13126 2818 13186 2894
rect 18413 2891 18479 2894
rect 20253 2954 20319 2957
rect 22000 2954 22800 2984
rect 20253 2952 22800 2954
rect 20253 2896 20258 2952
rect 20314 2896 22800 2952
rect 20253 2894 22800 2896
rect 20253 2891 20319 2894
rect 22000 2864 22800 2894
rect 10593 2816 13186 2818
rect 10593 2760 10598 2816
rect 10654 2760 13186 2816
rect 10593 2758 13186 2760
rect 17493 2818 17559 2821
rect 18689 2818 18755 2821
rect 17493 2816 18755 2818
rect 17493 2760 17498 2816
rect 17554 2760 18694 2816
rect 18750 2760 18755 2816
rect 17493 2758 18755 2760
rect 10593 2755 10659 2758
rect 17493 2755 17559 2758
rect 18689 2755 18755 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 800 2576
rect 2313 2546 2379 2549
rect 0 2544 2379 2546
rect 0 2488 2318 2544
rect 2374 2488 2379 2544
rect 0 2486 2379 2488
rect 0 2456 800 2486
rect 2313 2483 2379 2486
rect 2773 2546 2839 2549
rect 4889 2546 4955 2549
rect 6821 2546 6887 2549
rect 2773 2544 6887 2546
rect 2773 2488 2778 2544
rect 2834 2488 4894 2544
rect 4950 2488 6826 2544
rect 6882 2488 6887 2544
rect 2773 2486 6887 2488
rect 2773 2483 2839 2486
rect 4889 2483 4955 2486
rect 6821 2483 6887 2486
rect 18597 2546 18663 2549
rect 19241 2546 19307 2549
rect 22000 2546 22800 2576
rect 18597 2544 22800 2546
rect 18597 2488 18602 2544
rect 18658 2488 19246 2544
rect 19302 2488 22800 2544
rect 18597 2486 22800 2488
rect 18597 2483 18663 2486
rect 19241 2483 19307 2486
rect 22000 2456 22800 2486
rect 4376 2208 4696 2209
rect 0 2138 800 2168
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 3233 2138 3299 2141
rect 0 2136 3299 2138
rect 0 2080 3238 2136
rect 3294 2080 3299 2136
rect 0 2078 3299 2080
rect 0 2048 800 2078
rect 3233 2075 3299 2078
rect 20161 2138 20227 2141
rect 22000 2138 22800 2168
rect 20161 2136 22800 2138
rect 20161 2080 20166 2136
rect 20222 2080 22800 2136
rect 20161 2078 22800 2080
rect 20161 2075 20227 2078
rect 22000 2048 22800 2078
rect 4613 2002 4679 2005
rect 4838 2002 4844 2004
rect 4613 2000 4844 2002
rect 4613 1944 4618 2000
rect 4674 1944 4844 2000
rect 4613 1942 4844 1944
rect 4613 1939 4679 1942
rect 4838 1940 4844 1942
rect 4908 1940 4914 2004
rect 0 1730 800 1760
rect 2497 1730 2563 1733
rect 0 1728 2563 1730
rect 0 1672 2502 1728
rect 2558 1672 2563 1728
rect 0 1670 2563 1672
rect 0 1640 800 1670
rect 2497 1667 2563 1670
rect 18689 1730 18755 1733
rect 22000 1730 22800 1760
rect 18689 1728 22800 1730
rect 18689 1672 18694 1728
rect 18750 1672 22800 1728
rect 18689 1670 22800 1672
rect 18689 1667 18755 1670
rect 22000 1640 22800 1670
rect 0 1322 800 1352
rect 3325 1322 3391 1325
rect 0 1320 3391 1322
rect 0 1264 3330 1320
rect 3386 1264 3391 1320
rect 0 1262 3391 1264
rect 0 1232 800 1262
rect 3325 1259 3391 1262
rect 20621 1322 20687 1325
rect 22000 1322 22800 1352
rect 20621 1320 22800 1322
rect 20621 1264 20626 1320
rect 20682 1264 22800 1320
rect 20621 1262 22800 1264
rect 20621 1259 20687 1262
rect 22000 1232 22800 1262
rect 0 914 800 944
rect 1761 914 1827 917
rect 0 912 1827 914
rect 0 856 1766 912
rect 1822 856 1827 912
rect 0 854 1827 856
rect 0 824 800 854
rect 1761 851 1827 854
rect 18781 914 18847 917
rect 22000 914 22800 944
rect 18781 912 22800 914
rect 18781 856 18786 912
rect 18842 856 22800 912
rect 18781 854 22800 856
rect 18781 851 18847 854
rect 22000 824 22800 854
rect 0 506 800 536
rect 3785 506 3851 509
rect 0 504 3851 506
rect 0 448 3790 504
rect 3846 448 3851 504
rect 0 446 3851 448
rect 0 416 800 446
rect 3785 443 3851 446
rect 19149 506 19215 509
rect 22000 506 22800 536
rect 19149 504 22800 506
rect 19149 448 19154 504
rect 19210 448 22800 504
rect 19149 446 22800 448
rect 19149 443 19215 446
rect 22000 416 22800 446
rect 0 234 800 264
rect 4153 234 4219 237
rect 0 232 4219 234
rect 0 176 4158 232
rect 4214 176 4219 232
rect 0 174 4219 176
rect 0 144 800 174
rect 4153 171 4219 174
rect 17677 234 17743 237
rect 22000 234 22800 264
rect 17677 232 22800 234
rect 17677 176 17682 232
rect 17738 176 22800 232
rect 17677 174 22800 176
rect 17677 171 17743 174
rect 22000 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 5028 19076 5092 19140
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 8524 17912 8588 17916
rect 8524 17856 8538 17912
rect 8538 17856 8588 17912
rect 8524 17852 8588 17856
rect 8340 17580 8404 17644
rect 9076 17580 9140 17644
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 9812 17172 9876 17236
rect 7604 17036 7668 17100
rect 8708 17096 8772 17100
rect 8708 17040 8758 17096
rect 8758 17040 8772 17096
rect 8708 17036 8772 17040
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 8892 16492 8956 16556
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 5212 15812 5276 15876
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 12940 15540 13004 15604
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 4844 15192 4908 15196
rect 4844 15136 4858 15192
rect 4858 15136 4908 15192
rect 4844 15132 4908 15136
rect 11836 15464 11900 15468
rect 11836 15408 11850 15464
rect 11850 15408 11900 15464
rect 11836 15404 11900 15408
rect 13676 15328 13740 15332
rect 13676 15272 13690 15328
rect 13690 15272 13740 15328
rect 13676 15268 13740 15272
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 15148 15132 15212 15196
rect 7052 14724 7116 14788
rect 8340 14784 8404 14788
rect 8340 14728 8390 14784
rect 8390 14728 8404 14784
rect 8340 14724 8404 14728
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 9628 14588 9692 14652
rect 12020 14724 12084 14788
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 20116 13908 20180 13972
rect 10364 13772 10428 13836
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 11652 13500 11716 13564
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 6868 12548 6932 12612
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 10180 12548 10244 12612
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 12204 12276 12268 12340
rect 7420 12140 7484 12204
rect 6868 12004 6932 12068
rect 10180 12064 10244 12068
rect 10180 12008 10230 12064
rect 10230 12008 10244 12064
rect 10180 12004 10244 12008
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 5028 11732 5092 11796
rect 4844 11596 4908 11660
rect 5028 11656 5092 11660
rect 5028 11600 5042 11656
rect 5042 11600 5092 11656
rect 5028 11596 5092 11600
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 12388 11324 12452 11388
rect 9812 11248 9876 11252
rect 9812 11192 9826 11248
rect 9826 11192 9876 11248
rect 9812 11188 9876 11192
rect 9444 11052 9508 11116
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7604 10780 7668 10844
rect 8524 10644 8588 10708
rect 18644 10508 18708 10572
rect 8892 10372 8956 10436
rect 10364 10372 10428 10436
rect 14044 10432 14108 10436
rect 14044 10376 14058 10432
rect 14058 10376 14108 10432
rect 14044 10372 14108 10376
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 5212 10296 5276 10300
rect 5212 10240 5226 10296
rect 5226 10240 5276 10296
rect 5212 10236 5276 10240
rect 20116 10100 20180 10164
rect 13676 10024 13740 10028
rect 13676 9968 13726 10024
rect 13726 9968 13740 10024
rect 13676 9964 13740 9968
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 11652 9556 11716 9620
rect 12940 9556 13004 9620
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 7236 9148 7300 9212
rect 13676 9420 13740 9484
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 8708 9148 8772 9212
rect 11836 9208 11900 9212
rect 11836 9152 11886 9208
rect 11886 9152 11900 9208
rect 11836 9148 11900 9152
rect 9628 8876 9692 8940
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 9076 8740 9140 8804
rect 10180 8740 10244 8804
rect 10548 8800 10612 8804
rect 10548 8744 10562 8800
rect 10562 8744 10612 8800
rect 10548 8740 10612 8744
rect 12020 8740 12084 8804
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 12204 8060 12268 8124
rect 15148 7788 15212 7852
rect 7236 7652 7300 7716
rect 11100 7652 11164 7716
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 10548 7516 10612 7580
rect 9444 7244 9508 7308
rect 9812 7244 9876 7308
rect 14044 7244 14108 7308
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 18828 6972 18892 7036
rect 12388 6836 12452 6900
rect 13676 6836 13740 6900
rect 12204 6700 12268 6764
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7420 6428 7484 6492
rect 18644 6428 18708 6492
rect 12388 6292 12452 6356
rect 12204 6156 12268 6220
rect 4844 6020 4908 6084
rect 7052 6020 7116 6084
rect 10180 6080 10244 6084
rect 10180 6024 10230 6080
rect 10230 6024 10244 6080
rect 10180 6020 10244 6024
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 5028 5204 5092 5268
rect 8524 5264 8588 5268
rect 8524 5208 8574 5264
rect 8574 5208 8588 5264
rect 8524 5204 8588 5208
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 15148 4388 15212 4452
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 11100 3708 11164 3772
rect 9628 3436 9692 3500
rect 18828 3300 18892 3364
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 4844 3164 4908 3228
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 4844 1940 4908 2004
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 5027 19140 5093 19141
rect 5027 19076 5028 19140
rect 5092 19076 5093 19140
rect 5027 19075 5093 19076
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4843 15196 4909 15197
rect 4843 15132 4844 15196
rect 4908 15132 4909 15196
rect 4843 15131 4909 15132
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4846 11661 4906 15131
rect 5030 11797 5090 19075
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7603 17100 7669 17101
rect 7603 17036 7604 17100
rect 7668 17036 7669 17100
rect 7603 17035 7669 17036
rect 5211 15876 5277 15877
rect 5211 15812 5212 15876
rect 5276 15812 5277 15876
rect 5211 15811 5277 15812
rect 5027 11796 5093 11797
rect 5027 11732 5028 11796
rect 5092 11732 5093 11796
rect 5027 11731 5093 11732
rect 4843 11660 4909 11661
rect 4843 11596 4844 11660
rect 4908 11596 4909 11660
rect 4843 11595 4909 11596
rect 5027 11660 5093 11661
rect 5027 11596 5028 11660
rect 5092 11596 5093 11660
rect 5027 11595 5093 11596
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4843 6084 4909 6085
rect 4843 6020 4844 6084
rect 4908 6020 4909 6084
rect 4843 6019 4909 6020
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4846 3229 4906 6019
rect 5030 5269 5090 11595
rect 5214 10301 5274 15811
rect 7051 14788 7117 14789
rect 7051 14724 7052 14788
rect 7116 14724 7117 14788
rect 7051 14723 7117 14724
rect 6867 12612 6933 12613
rect 6867 12548 6868 12612
rect 6932 12548 6933 12612
rect 6867 12547 6933 12548
rect 6870 12069 6930 12547
rect 6867 12068 6933 12069
rect 6867 12004 6868 12068
rect 6932 12004 6933 12068
rect 6867 12003 6933 12004
rect 5211 10300 5277 10301
rect 5211 10236 5212 10300
rect 5276 10236 5277 10300
rect 5211 10235 5277 10236
rect 7054 6085 7114 14723
rect 7419 12204 7485 12205
rect 7419 12140 7420 12204
rect 7484 12140 7485 12204
rect 7419 12139 7485 12140
rect 7235 9212 7301 9213
rect 7235 9148 7236 9212
rect 7300 9148 7301 9212
rect 7235 9147 7301 9148
rect 7238 7717 7298 9147
rect 7235 7716 7301 7717
rect 7235 7652 7236 7716
rect 7300 7652 7301 7716
rect 7235 7651 7301 7652
rect 7422 6493 7482 12139
rect 7606 10845 7666 17035
rect 7808 16896 8128 17920
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 8523 17916 8589 17917
rect 8523 17852 8524 17916
rect 8588 17852 8589 17916
rect 8523 17851 8589 17852
rect 8339 17644 8405 17645
rect 8339 17580 8340 17644
rect 8404 17580 8405 17644
rect 8339 17579 8405 17580
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 8342 14789 8402 17579
rect 8339 14788 8405 14789
rect 8339 14724 8340 14788
rect 8404 14724 8405 14788
rect 8339 14723 8405 14724
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7603 10844 7669 10845
rect 7603 10780 7604 10844
rect 7668 10780 7669 10844
rect 7603 10779 7669 10780
rect 7808 10368 8128 11392
rect 8526 10709 8586 17851
rect 9075 17644 9141 17645
rect 9075 17580 9076 17644
rect 9140 17580 9141 17644
rect 9075 17579 9141 17580
rect 8707 17100 8773 17101
rect 8707 17036 8708 17100
rect 8772 17036 8773 17100
rect 8707 17035 8773 17036
rect 8523 10708 8589 10709
rect 8523 10644 8524 10708
rect 8588 10644 8589 10708
rect 8523 10643 8589 10644
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7419 6492 7485 6493
rect 7419 6428 7420 6492
rect 7484 6428 7485 6492
rect 7419 6427 7485 6428
rect 7051 6084 7117 6085
rect 7051 6020 7052 6084
rect 7116 6020 7117 6084
rect 7051 6019 7117 6020
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 5027 5268 5093 5269
rect 5027 5204 5028 5268
rect 5092 5204 5093 5268
rect 5027 5203 5093 5204
rect 7808 4928 8128 5952
rect 8526 5269 8586 10643
rect 8710 9213 8770 17035
rect 8891 16556 8957 16557
rect 8891 16492 8892 16556
rect 8956 16492 8957 16556
rect 8891 16491 8957 16492
rect 8894 10437 8954 16491
rect 8891 10436 8957 10437
rect 8891 10372 8892 10436
rect 8956 10372 8957 10436
rect 8891 10371 8957 10372
rect 8707 9212 8773 9213
rect 8707 9148 8708 9212
rect 8772 9148 8773 9212
rect 8707 9147 8773 9148
rect 9078 8805 9138 17579
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 9811 17236 9877 17237
rect 9811 17172 9812 17236
rect 9876 17172 9877 17236
rect 9811 17171 9877 17172
rect 9627 14652 9693 14653
rect 9627 14588 9628 14652
rect 9692 14588 9693 14652
rect 9627 14587 9693 14588
rect 9443 11116 9509 11117
rect 9443 11052 9444 11116
rect 9508 11052 9509 11116
rect 9443 11051 9509 11052
rect 9075 8804 9141 8805
rect 9075 8740 9076 8804
rect 9140 8740 9141 8804
rect 9075 8739 9141 8740
rect 9446 7309 9506 11051
rect 9630 10570 9690 14587
rect 9814 11253 9874 17171
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 12939 15604 13005 15605
rect 12939 15540 12940 15604
rect 13004 15540 13005 15604
rect 12939 15539 13005 15540
rect 11835 15468 11901 15469
rect 11835 15404 11836 15468
rect 11900 15404 11901 15468
rect 11835 15403 11901 15404
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 10363 13836 10429 13837
rect 10363 13772 10364 13836
rect 10428 13772 10429 13836
rect 10363 13771 10429 13772
rect 10179 12612 10245 12613
rect 10179 12548 10180 12612
rect 10244 12548 10245 12612
rect 10179 12547 10245 12548
rect 10182 12069 10242 12547
rect 10179 12068 10245 12069
rect 10179 12004 10180 12068
rect 10244 12004 10245 12068
rect 10179 12003 10245 12004
rect 9811 11252 9877 11253
rect 9811 11188 9812 11252
rect 9876 11188 9877 11252
rect 9811 11187 9877 11188
rect 9630 10510 9874 10570
rect 9627 8940 9693 8941
rect 9627 8876 9628 8940
rect 9692 8876 9693 8940
rect 9627 8875 9693 8876
rect 9443 7308 9509 7309
rect 9443 7244 9444 7308
rect 9508 7244 9509 7308
rect 9443 7243 9509 7244
rect 8523 5268 8589 5269
rect 8523 5204 8524 5268
rect 8588 5204 8589 5268
rect 8523 5203 8589 5204
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 4843 3228 4909 3229
rect 4843 3164 4844 3228
rect 4908 3164 4909 3228
rect 4843 3163 4909 3164
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 4846 2005 4906 3163
rect 7808 2752 8128 3776
rect 9630 3501 9690 8875
rect 9814 7309 9874 10510
rect 10366 10437 10426 13771
rect 11240 13088 11560 14112
rect 11651 13564 11717 13565
rect 11651 13500 11652 13564
rect 11716 13500 11717 13564
rect 11651 13499 11717 13500
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 10363 10436 10429 10437
rect 10363 10372 10364 10436
rect 10428 10372 10429 10436
rect 10363 10371 10429 10372
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 10179 8804 10245 8805
rect 10179 8740 10180 8804
rect 10244 8740 10245 8804
rect 10179 8739 10245 8740
rect 10547 8804 10613 8805
rect 10547 8740 10548 8804
rect 10612 8740 10613 8804
rect 10547 8739 10613 8740
rect 9811 7308 9877 7309
rect 9811 7244 9812 7308
rect 9876 7244 9877 7308
rect 9811 7243 9877 7244
rect 10182 6085 10242 8739
rect 10550 7581 10610 8739
rect 11240 8736 11560 9760
rect 11654 9621 11714 13499
rect 11651 9620 11717 9621
rect 11651 9556 11652 9620
rect 11716 9556 11717 9620
rect 11651 9555 11717 9556
rect 11838 9213 11898 15403
rect 12019 14788 12085 14789
rect 12019 14724 12020 14788
rect 12084 14724 12085 14788
rect 12019 14723 12085 14724
rect 11835 9212 11901 9213
rect 11835 9148 11836 9212
rect 11900 9148 11901 9212
rect 11835 9147 11901 9148
rect 12022 8805 12082 14723
rect 12203 12340 12269 12341
rect 12203 12276 12204 12340
rect 12268 12276 12269 12340
rect 12203 12275 12269 12276
rect 12019 8804 12085 8805
rect 12019 8740 12020 8804
rect 12084 8740 12085 8804
rect 12019 8739 12085 8740
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11099 7716 11165 7717
rect 11099 7652 11100 7716
rect 11164 7652 11165 7716
rect 11099 7651 11165 7652
rect 10547 7580 10613 7581
rect 10547 7516 10548 7580
rect 10612 7516 10613 7580
rect 10547 7515 10613 7516
rect 10179 6084 10245 6085
rect 10179 6020 10180 6084
rect 10244 6020 10245 6084
rect 10179 6019 10245 6020
rect 11102 3773 11162 7651
rect 11240 7648 11560 8672
rect 12206 8125 12266 12275
rect 12387 11388 12453 11389
rect 12387 11324 12388 11388
rect 12452 11324 12453 11388
rect 12387 11323 12453 11324
rect 12203 8124 12269 8125
rect 12203 8060 12204 8124
rect 12268 8060 12269 8124
rect 12203 8059 12269 8060
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 12390 6901 12450 11323
rect 12942 9621 13002 15539
rect 13675 15332 13741 15333
rect 13675 15268 13676 15332
rect 13740 15268 13741 15332
rect 13675 15267 13741 15268
rect 13678 10029 13738 15267
rect 14672 14720 14992 15744
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 15147 15196 15213 15197
rect 15147 15132 15148 15196
rect 15212 15132 15213 15196
rect 15147 15131 15213 15132
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14043 10436 14109 10437
rect 14043 10372 14044 10436
rect 14108 10372 14109 10436
rect 14043 10371 14109 10372
rect 13675 10028 13741 10029
rect 13675 9964 13676 10028
rect 13740 9964 13741 10028
rect 13675 9963 13741 9964
rect 12939 9620 13005 9621
rect 12939 9556 12940 9620
rect 13004 9556 13005 9620
rect 12939 9555 13005 9556
rect 13678 9485 13738 9963
rect 13675 9484 13741 9485
rect 13675 9420 13676 9484
rect 13740 9420 13741 9484
rect 13675 9419 13741 9420
rect 13678 6901 13738 9419
rect 14046 7309 14106 10371
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14043 7308 14109 7309
rect 14043 7244 14044 7308
rect 14108 7244 14109 7308
rect 14043 7243 14109 7244
rect 14672 7104 14992 8128
rect 15150 7853 15210 15131
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 20115 13972 20181 13973
rect 20115 13908 20116 13972
rect 20180 13908 20181 13972
rect 20115 13907 20181 13908
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18643 10572 18709 10573
rect 18643 10508 18644 10572
rect 18708 10508 18709 10572
rect 18643 10507 18709 10508
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 15147 7852 15213 7853
rect 15147 7788 15148 7852
rect 15212 7788 15213 7852
rect 15147 7787 15213 7788
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 12387 6900 12453 6901
rect 12387 6836 12388 6900
rect 12452 6836 12453 6900
rect 12387 6835 12453 6836
rect 13675 6900 13741 6901
rect 13675 6836 13676 6900
rect 13740 6836 13741 6900
rect 13675 6835 13741 6836
rect 12203 6764 12269 6765
rect 12203 6700 12204 6764
rect 12268 6700 12269 6764
rect 12203 6699 12269 6700
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 12206 6221 12266 6699
rect 12390 6357 12450 6835
rect 12387 6356 12453 6357
rect 12387 6292 12388 6356
rect 12452 6292 12453 6356
rect 12387 6291 12453 6292
rect 12203 6220 12269 6221
rect 12203 6156 12204 6220
rect 12268 6156 12269 6220
rect 12203 6155 12269 6156
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11099 3772 11165 3773
rect 11099 3708 11100 3772
rect 11164 3708 11165 3772
rect 11099 3707 11165 3708
rect 9627 3500 9693 3501
rect 9627 3436 9628 3500
rect 9692 3436 9693 3500
rect 9627 3435 9693 3436
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 15150 4453 15210 7787
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18646 6493 18706 10507
rect 20118 10165 20178 13907
rect 20115 10164 20181 10165
rect 20115 10100 20116 10164
rect 20180 10100 20181 10164
rect 20115 10099 20181 10100
rect 18827 7036 18893 7037
rect 18827 6972 18828 7036
rect 18892 6972 18893 7036
rect 18827 6971 18893 6972
rect 18643 6492 18709 6493
rect 18643 6428 18644 6492
rect 18708 6428 18709 6492
rect 18643 6427 18709 6428
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 15147 4452 15213 4453
rect 15147 4388 15148 4452
rect 15212 4388 15213 4452
rect 15147 4387 15213 4388
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18830 3365 18890 6971
rect 18827 3364 18893 3365
rect 18827 3300 18828 3364
rect 18892 3300 18893 3364
rect 18827 3299 18893 3300
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 4843 2004 4909 2005
rect 4843 1940 4844 2004
rect 4908 1940 4909 2004
rect 4843 1939 4909 1940
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1608762545
transform 1 0 20424 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608762545
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608762545
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_216
timestamp 1608762545
transform 1 0 20976 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608762545
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1608762545
transform 1 0 19872 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1608762545
transform 1 0 19320 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_193
timestamp 1608762545
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1608762545
transform 1 0 19228 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1608762545
transform 1 0 18308 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608762545
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_176
timestamp 1608762545
transform 1 0 17296 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1608762545
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1608762545
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1608762545
transform 1 0 15824 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608762545
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_148
timestamp 1608762545
transform 1 0 14720 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1608762545
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_164
timestamp 1608762545
transform 1 0 16192 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1608762545
transform 1 0 13248 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_131
timestamp 1608762545
transform 1 0 13156 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_136
timestamp 1608762545
transform 1 0 13616 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608762545
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1608762545
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1608762545
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_125
timestamp 1608762545
transform 1 0 12604 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608762545
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1608762545
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1608762545
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 6900 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1608762545
transform 1 0 7544 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_69
timestamp 1608762545
transform 1 0 7452 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_79
timestamp 1608762545
transform 1 0 8372 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608762545
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_50
timestamp 1608762545
transform 1 0 5704 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1608762545
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 4232 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608762545
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1608762545
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608762545
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608762545
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608762545
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1608762545
transform 1 0 20424 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608762545
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_209
timestamp 1608762545
transform 1 0 20332 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_216
timestamp 1608762545
transform 1 0 20976 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608762545
transform 1 0 18860 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1608762545
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1608762545
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_E_FTB01
timestamp 1608762545
transform 1 0 18308 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1608762545
transform 1 0 17388 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1608762545
transform 1 0 16836 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608762545
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_184
timestamp 1608762545
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1608762545
transform 1 0 14536 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1608762545
transform 1 0 14904 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1608762545
transform 1 0 15272 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_W_FTB01
timestamp 1608762545
transform 1 0 15916 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_158
timestamp 1608762545
transform 1 0 15640 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1608762545
transform 1 0 13064 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1608762545
transform 1 0 13432 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1608762545
transform 1 0 13800 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1608762545
transform 1 0 14168 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1608762545
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1608762545
transform 1 0 11408 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 12512 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608762545
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1608762545
transform 1 0 10856 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1608762545
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1608762545
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608762545
transform 1 0 10120 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1608762545
transform 1 0 10488 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 9568 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1608762545
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 6900 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608762545
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1608762545
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608762545
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1608762545
transform 1 0 6348 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_62
timestamp 1608762545
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 4876 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608762545
transform 1 0 4048 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1608762545
transform 1 0 3128 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_21
timestamp 1608762545
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_31
timestamp 1608762545
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608762545
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1608762545
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_15
timestamp 1608762545
transform 1 0 2484 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608762545
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608762545
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608762545
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608762545
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1608762545
transform 1 0 18492 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1608762545
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1608762545
transform 1 0 19688 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1608762545
transform 1 0 19136 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1608762545
transform 1 0 19044 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1608762545
transform 1 0 16560 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_W_FTB01
timestamp 1608762545
transform 1 0 17940 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_172
timestamp 1608762545
transform 1 0 16928 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_180
timestamp 1608762545
transform 1 0 17664 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608762545
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1608762545
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_160
timestamp 1608762545
transform 1 0 15824 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 12788 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 14260 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 11316 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_109
timestamp 1608762545
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608762545
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 10580 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608762545
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608762545
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_102
timestamp 1608762545
transform 1 0 10488 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 7912 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_72
timestamp 1608762545
transform 1 0 7728 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 6256 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1608762545
transform 1 0 5428 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608762545
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 4876 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608762545
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608762545
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1608762545
transform 1 0 2760 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608762545
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1608762545
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_15
timestamp 1608762545
transform 1 0 2484 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_E_FTB01
timestamp 1608762545
transform 1 0 20424 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608762545
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_216
timestamp 1608762545
transform 1 0 20976 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1608762545
transform 1 0 19872 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1608762545
transform 1 0 19320 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_196
timestamp 1608762545
transform 1 0 19136 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1608762545
transform 1 0 17020 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608762545
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_177
timestamp 1608762545
transform 1 0 17388 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1608762545
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_153
timestamp 1608762545
transform 1 0 15180 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_165
timestamp 1608762545
transform 1 0 16284 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1608762545
transform 1 0 13248 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_141
timestamp 1608762545
transform 1 0 14076 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1608762545
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608762545
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_115
timestamp 1608762545
transform 1 0 11684 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1608762545
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 10212 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608762545
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_85
timestamp 1608762545
transform 1 0 8924 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1608762545
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608762545
transform 1 0 8096 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608762545
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_66
timestamp 1608762545
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608762545
transform 1 0 5612 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608762545
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_45
timestamp 1608762545
transform 1 0 5244 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1608762545
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1608762545
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608762545
transform 1 0 4416 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608762545
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608762545
transform 1 0 2944 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608762545
transform 1 0 2116 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608762545
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608762545
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608762545
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608762545
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608762545
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608762545
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1608762545
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1608762545
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1608762545
transform 1 0 19688 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1608762545
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608762545
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1608762545
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1608762545
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1608762545
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 13432 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1608762545
transform 1 0 11776 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608762545
transform 1 0 10948 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608762545
transform 1 0 12604 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1608762545
transform 1 0 10120 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608762545
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1608762545
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1608762545
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_97
timestamp 1608762545
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1608762545
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1608762545
transform 1 0 7176 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608762545
transform 1 0 5980 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_62
timestamp 1608762545
transform 1 0 6808 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 4508 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608762545
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_24
timestamp 1608762545
transform 1 0 3312 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1608762545
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1608762545
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_36
timestamp 1608762545
transform 1 0 4416 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608762545
transform 1 0 1472 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 1840 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608762545
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1608762545
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608762545
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608762545
transform 1 0 20976 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1608762545
transform 1 0 20424 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608762545
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608762545
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608762545
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608762545
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608762545
transform 1 0 20056 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608762545
transform 1 0 19688 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1608762545
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_198
timestamp 1608762545
transform 1 0 19320 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1608762545
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_196
timestamp 1608762545
transform 1 0 19136 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1608762545
transform 1 0 16744 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608762545
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_174
timestamp 1608762545
transform 1 0 17112 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_186
timestamp 1608762545
transform 1 0 18216 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_176
timestamp 1608762545
transform 1 0 17296 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1608762545
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608762545
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 14720 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608762545
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1608762545
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_164
timestamp 1608762545
transform 1 0 16192 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 13248 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1608762545
transform 1 0 13432 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1608762545
transform 1 0 14260 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1608762545
transform 1 0 12604 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_26_124
timestamp 1608762545
transform 1 0 12512 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1608762545
transform 1 0 11684 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1608762545
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608762545
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1608762545
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608762545
transform 1 0 11132 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1608762545
transform 1 0 11408 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1608762545
transform 1 0 10856 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_108
timestamp 1608762545
transform 1 0 11040 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 9568 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608762545
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608762545
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1608762545
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1608762545
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1608762545
transform 1 0 9200 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608762545
transform 1 0 8096 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 7176 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1608762545
transform 1 0 8648 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1608762545
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1608762545
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1608762545
transform 1 0 7636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_75
timestamp 1608762545
transform 1 0 8004 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608762545
transform 1 0 5520 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608762545
transform 1 0 6164 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1608762545
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608762545
transform 1 0 5336 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608762545
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_47
timestamp 1608762545
transform 1 0 5428 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1608762545
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608762545
transform 1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1608762545
transform 1 0 4508 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1608762545
transform 1 0 3772 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1608762545
transform 1 0 4600 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608762545
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1608762545
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1608762545
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_36
timestamp 1608762545
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608762545
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608762545
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1608762545
transform 1 0 2944 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1608762545
transform 1 0 2116 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1608762545
transform 1 0 2576 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1608762545
transform 1 0 1748 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608762545
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608762545
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608762545
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608762545
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608762545
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608762545
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1608762545
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608762545
transform 1 0 20148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 19504 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_188
timestamp 1608762545
transform 1 0 18400 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_206
timestamp 1608762545
transform 1 0 20056 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1608762545
transform 1 0 17204 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1608762545
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608762545
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1608762545
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1608762545
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1608762545
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1608762545
transform 1 0 14720 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1608762545
transform 1 0 15548 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_165
timestamp 1608762545
transform 1 0 16284 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608762545
transform 1 0 13064 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1608762545
transform 1 0 13892 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1608762545
transform 1 0 12972 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 10856 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608762545
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_105
timestamp 1608762545
transform 1 0 10764 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_123
timestamp 1608762545
transform 1 0 12420 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1608762545
transform 1 0 8832 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1608762545
transform 1 0 9936 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_93
timestamp 1608762545
transform 1 0 9660 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1608762545
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1608762545
transform 1 0 8280 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 5244 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608762545
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1608762545
transform 1 0 4416 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1608762545
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_29
timestamp 1608762545
transform 1 0 3772 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1608762545
transform 1 0 4140 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608762545
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608762545
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 2300 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608762545
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1608762545
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608762545
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608762545
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608762545
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608762545
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608762545
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1608762545
transform 1 0 18492 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608762545
transform 1 0 20056 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_195
timestamp 1608762545
transform 1 0 19044 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_203
timestamp 1608762545
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1608762545
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608762545
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 16192 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608762545
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608762545
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_157
timestamp 1608762545
transform 1 0 15548 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_163
timestamp 1608762545
transform 1 0 16100 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608762545
transform 1 0 13340 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1608762545
transform 1 0 14168 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1608762545
transform 1 0 12880 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_132
timestamp 1608762545
transform 1 0 13248 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608762545
transform 1 0 12052 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_111
timestamp 1608762545
transform 1 0 11316 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 9844 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608762545
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1608762545
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608762545
transform 1 0 7636 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1608762545
transform 1 0 8740 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1608762545
transform 1 0 7912 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_82
timestamp 1608762545
transform 1 0 8648 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608762545
transform 1 0 6808 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1608762545
transform 1 0 5980 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_52
timestamp 1608762545
transform 1 0 5888 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608762545
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 4416 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608762545
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1608762545
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 1472 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1608762545
transform 1 0 2852 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1608762545
transform 1 0 2024 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608762545
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608762545
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608762545
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608762545
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608762545
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1608762545
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608762545
transform 1 0 20148 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608762545
transform 1 0 19780 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608762545
transform 1 0 19412 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_193
timestamp 1608762545
transform 1 0 18860 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1608762545
transform 1 0 17020 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1608762545
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608762545
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1608762545
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 15548 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_156
timestamp 1608762545
transform 1 0 15456 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1608762545
transform 1 0 13524 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1608762545
transform 1 0 12696 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_144
timestamp 1608762545
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608762545
transform 1 0 11500 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608762545
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1608762545
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 8832 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1608762545
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1608762545
transform 1 0 10304 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1608762545
transform 1 0 7176 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1608762545
transform 1 0 8004 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608762545
transform 1 0 5336 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608762545
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_43
timestamp 1608762545
transform 1 0 5060 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_55
timestamp 1608762545
transform 1 0 6164 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1608762545
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608762545
transform 1 0 4232 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1608762545
transform 1 0 3404 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1608762545
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1608762545
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1608762545
transform 1 0 2116 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608762545
transform 1 0 2484 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608762545
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608762545
transform 1 0 2852 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608762545
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608762545
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608762545
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608762545
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1608762545
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1608762545
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 19596 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 20148 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_191
timestamp 1608762545
transform 1 0 18676 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1608762545
transform 1 0 19412 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 17204 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_168
timestamp 1608762545
transform 1 0 16560 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_174
timestamp 1608762545
transform 1 0 17112 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608762545
transform 1 0 15732 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608762545
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1608762545
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1608762545
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1608762545
transform 1 0 14352 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 13984 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_143
timestamp 1608762545
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 12512 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1608762545
transform 1 0 10764 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1608762545
transform 1 0 11592 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_123
timestamp 1608762545
transform 1 0 12420 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608762545
transform 1 0 9936 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608762545
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1608762545
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1608762545
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 7912 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 7636 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608762545
transform 1 0 5980 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1608762545
transform 1 0 6808 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_48
timestamp 1608762545
transform 1 0 5520 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_52
timestamp 1608762545
transform 1 0 5888 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1608762545
transform 1 0 3128 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608762545
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1608762545
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1608762545
transform 1 0 1564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 1932 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608762545
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1608762545
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_19
timestamp 1608762545
transform 1 0 2852 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 20516 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608762545
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1608762545
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1608762545
transform 1 0 18860 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1608762545
transform 1 0 19688 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608762545
transform 1 0 17020 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608762545
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608762545
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1608762545
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608762545
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 15364 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 13892 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608762545
transform 1 0 11132 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1608762545
transform 1 0 11500 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608762545
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_112
timestamp 1608762545
transform 1 0 11408 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608762545
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1608762545
transform 1 0 9476 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_90
timestamp 1608762545
transform 1 0 9384 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1608762545
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608762545
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 5980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_56
timestamp 1608762545
transform 1 0 6256 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1608762545
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 4508 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_34
timestamp 1608762545
transform 1 0 4232 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1608762545
transform 1 0 1564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 2760 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 1932 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608762545
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608762545
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_15
timestamp 1608762545
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608762545
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1608762545
transform 1 0 20516 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608762545
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608762545
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608762545
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608762545
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608762545
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 19136 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608762545
transform 1 0 18860 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1608762545
transform 1 0 19688 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 17664 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608762545
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608762545
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 16928 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1608762545
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1608762545
transform 1 0 17204 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_179
timestamp 1608762545
transform 1 0 17572 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608762545
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608762545
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1608762545
transform 1 0 16100 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1608762545
transform 1 0 15456 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1608762545
transform 1 0 14628 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608762545
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_165
timestamp 1608762545
transform 1 0 16284 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1608762545
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608762545
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1608762545
transform 1 0 13432 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1608762545
transform 1 0 13156 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1608762545
transform 1 0 14260 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1608762545
transform 1 0 14260 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608762545
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1608762545
transform 1 0 11224 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1608762545
transform 1 0 12604 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608762545
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1608762545
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_123
timestamp 1608762545
transform 1 0 12420 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_113
timestamp 1608762545
transform 1 0 11500 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1608762545
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1608762545
transform 1 0 10396 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1608762545
transform 1 0 10672 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608762545
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608762545
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1608762545
transform 1 0 10304 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1608762545
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_93
timestamp 1608762545
transform 1 0 9660 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_101
timestamp 1608762545
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 8004 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608762545
transform 1 0 8648 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608762545
transform 1 0 7820 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_74
timestamp 1608762545
transform 1 0 7912 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1608762545
transform 1 0 7360 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_72
timestamp 1608762545
transform 1 0 7728 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1608762545
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1608762545
transform 1 0 6532 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1608762545
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1608762545
transform 1 0 5244 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608762545
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_54
timestamp 1608762545
transform 1 0 6072 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1608762545
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 3220 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608762545
transform 1 0 4876 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1608762545
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608762545
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_39
timestamp 1608762545
transform 1 0 4692 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1608762545
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1608762545
transform 1 0 2944 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1608762545
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1608762545
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_18
timestamp 1608762545
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1608762545
transform 1 0 1564 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1608762545
transform 1 0 1932 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 1564 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608762545
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608762545
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1608762545
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1608762545
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608762545
transform 1 0 20976 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608762545
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608762545
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_215
timestamp 1608762545
transform 1 0 20884 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608762545
transform 1 0 19044 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 19320 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 17572 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1608762545
transform 1 0 16744 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608762545
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608762545
transform 1 0 14352 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 13708 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_130
timestamp 1608762545
transform 1 0 13064 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_136
timestamp 1608762545
transform 1 0 13616 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_140
timestamp 1608762545
transform 1 0 13984 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 11592 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 10120 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608762545
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608762545
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1608762545
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1608762545
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1608762545
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1608762545
transform 1 0 7728 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_70
timestamp 1608762545
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 6072 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_44
timestamp 1608762545
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1608762545
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1608762545
transform 1 0 4324 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 3312 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608762545
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608762545
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1608762545
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1608762545
transform 1 0 1472 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608762545
transform 1 0 1840 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608762545
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1608762545
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 20516 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608762545
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1608762545
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1608762545
transform 1 0 18860 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1608762545
transform 1 0 19688 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608762545
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608762545
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1608762545
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 15732 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 14260 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1608762545
transform 1 0 13892 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1608762545
transform 1 0 11040 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608762545
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1608762545
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608762545
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608762545
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608762545
transform 1 0 9108 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_96
timestamp 1608762545
transform 1 0 9936 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1608762545
transform 1 0 8280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608762545
transform 1 0 5612 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1608762545
transform 1 0 5888 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608762545
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_46
timestamp 1608762545
transform 1 0 5336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1608762545
transform 1 0 4508 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608762545
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_23
timestamp 1608762545
transform 1 0 3220 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1608762545
transform 1 0 3588 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1608762545
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 1748 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608762545
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608762545
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608762545
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608762545
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608762545
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 19320 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1608762545
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1608762545
transform 1 0 19228 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608762545
transform 1 0 16928 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1608762545
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1608762545
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_175
timestamp 1608762545
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608762545
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1608762545
transform 1 0 16100 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608762545
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608762545
transform 1 0 14352 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1608762545
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 12604 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_122
timestamp 1608762545
transform 1 0 12328 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608762545
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 10488 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1608762545
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1608762545
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1608762545
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 7544 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 7268 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_63
timestamp 1608762545
transform 1 0 6900 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1608762545
transform 1 0 6072 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_49
timestamp 1608762545
transform 1 0 5612 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_53
timestamp 1608762545
transform 1 0 5980 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608762545
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608762545
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_32
timestamp 1608762545
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 2484 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1608762545
transform 1 0 1656 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608762545
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1608762545
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 20792 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608762545
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608762545
transform 1 0 18492 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1608762545
transform 1 0 19964 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1608762545
transform 1 0 18400 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1608762545
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608762545
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608762545
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1608762545
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608762545
transform 1 0 14628 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1608762545
transform 1 0 16100 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_156
timestamp 1608762545
transform 1 0 15456 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_162
timestamp 1608762545
transform 1 0 16008 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608762545
transform 1 0 14076 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1608762545
transform 1 0 13248 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 14352 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608762545
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1608762545
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608762545
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1608762545
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 9844 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1608762545
transform 1 0 9016 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608762545
transform 1 0 8188 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1608762545
transform 1 0 6992 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1608762545
transform 1 0 7820 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1608762545
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608762545
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608762545
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1608762545
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608762545
transform 1 0 4876 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608762545
transform 1 0 4048 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1608762545
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1608762545
transform 1 0 2392 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1608762545
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608762545
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1608762545
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608762545
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608762545
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608762545
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_217
timestamp 1608762545
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1608762545
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608762545
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608762545
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1608762545
transform 1 0 20240 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1608762545
transform 1 0 19412 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1608762545
transform 1 0 19596 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_193
timestamp 1608762545
transform 1 0 18860 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_194
timestamp 1608762545
transform 1 0 18952 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_200
timestamp 1608762545
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 17480 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1608762545
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608762545
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_175
timestamp 1608762545
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_170
timestamp 1608762545
transform 1 0 16744 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608762545
transform 1 0 14720 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608762545
transform 1 0 15548 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1608762545
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608762545
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608762545
transform 1 0 13892 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608762545
transform 1 0 13524 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1608762545
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1608762545
transform 1 0 13432 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1608762545
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1608762545
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1608762545
transform 1 0 11500 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608762545
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_119
timestamp 1608762545
transform 1 0 12052 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608762545
transform 1 0 10396 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1608762545
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1608762545
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608762545
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_90
timestamp 1608762545
transform 1 0 9384 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_100
timestamp 1608762545
transform 1 0 10304 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1608762545
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1608762545
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 7728 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608762545
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608762545
transform 1 0 6900 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 8280 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608762545
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1608762545
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608762545
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608762545
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1608762545
transform 1 0 5520 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_61
timestamp 1608762545
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1608762545
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 4784 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608762545
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_36
timestamp 1608762545
transform 1 0 4416 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1608762545
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1608762545
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1608762545
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 2944 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1608762545
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1608762545
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1608762545
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608762545
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608762545
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1608762545
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1608762545
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608762545
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608762545
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608762545
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608762545
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1608762545
transform 1 0 19964 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1608762545
transform 1 0 19136 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1608762545
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 16652 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608762545
transform 1 0 18124 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1608762545
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608762545
transform 1 0 15364 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608762545
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 16192 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1608762545
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1608762545
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1608762545
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608762545
transform 1 0 13984 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 11684 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_109
timestamp 1608762545
transform 1 0 11132 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608762545
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1608762545
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1608762545
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1608762545
transform 1 0 8096 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1608762545
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1608762545
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1608762545
transform 1 0 6256 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1608762545
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_44
timestamp 1608762545
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_55
timestamp 1608762545
transform 1 0 6164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608762545
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1608762545
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608762545
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1608762545
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608762545
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1608762545
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_11
timestamp 1608762545
transform 1 0 2116 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608762545
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_217
timestamp 1608762545
transform 1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608762545
transform 1 0 19872 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1608762545
transform 1 0 18860 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1608762545
transform 1 0 20240 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_202
timestamp 1608762545
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_207
timestamp 1608762545
transform 1 0 20148 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1608762545
transform 1 0 16928 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608762545
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608762545
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1608762545
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608762545
transform 1 0 14536 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1608762545
transform 1 0 16100 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_155
timestamp 1608762545
transform 1 0 15364 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 13708 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_134
timestamp 1608762545
transform 1 0 13432 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_140
timestamp 1608762545
transform 1 0 13984 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608762545
transform 1 0 11592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608762545
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608762545
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1608762545
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608762545
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1608762545
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 10120 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1608762545
transform 1 0 7636 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1608762545
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608762545
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608762545
transform 1 0 5428 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608762545
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_44
timestamp 1608762545
transform 1 0 5152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_56
timestamp 1608762545
transform 1 0 6256 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1608762545
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1608762545
transform 1 0 3220 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1608762545
transform 1 0 4048 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1608762545
transform 1 0 1472 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1608762545
transform 1 0 2392 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 1840 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608762545
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1608762545
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608762545
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608762545
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1608762545
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608762545
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608762545
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 19136 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1608762545
transform 1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608762545
transform 1 0 16744 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1608762545
transform 1 0 18032 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_179
timestamp 1608762545
transform 1 0 17572 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_183
timestamp 1608762545
transform 1 0 17940 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608762545
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1608762545
transform 1 0 14352 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_140
timestamp 1608762545
transform 1 0 13984 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 12512 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1608762545
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_123
timestamp 1608762545
transform 1 0 12420 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1608762545
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1608762545
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608762545
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608762545
transform 1 0 8740 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1608762545
transform 1 0 7912 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608762545
transform 1 0 7084 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608762545
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 5704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1608762545
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_53
timestamp 1608762545
transform 1 0 5980 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 4140 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1608762545
transform 1 0 3128 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608762545
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_21
timestamp 1608762545
transform 1 0 3036 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1608762545
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 1564 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608762545
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1608762545
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608762545
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_213
timestamp 1608762545
transform 1 0 20700 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1608762545
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 18400 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1608762545
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608762545
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1608762545
transform 1 0 17020 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608762545
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1608762545
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_187
timestamp 1608762545
transform 1 0 18308 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 15548 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1608762545
transform 1 0 14720 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608762545
transform 1 0 12696 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1608762545
transform 1 0 13064 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1608762545
transform 1 0 13892 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp 1608762545
transform 1 0 12972 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 10856 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608762545
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608762545
transform 1 0 10028 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1608762545
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1608762545
transform 1 0 8372 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608762545
transform 1 0 7084 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762545
transform 1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1608762545
transform 1 0 6900 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1608762545
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608762545
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1608762545
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1608762545
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 4508 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1608762545
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1608762545
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1608762545
transform 1 0 1932 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1608762545
transform 1 0 2760 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608762545
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608762545
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608762545
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1608762545
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608762545
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608762545
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1608762545
transform 1 0 19780 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 18308 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608762545
transform 1 0 17020 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_182
timestamp 1608762545
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_186
timestamp 1608762545
transform 1 0 18216 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608762545
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608762545
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1608762545
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_146
timestamp 1608762545
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1608762545
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_165
timestamp 1608762545
transform 1 0 16284 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608762545
transform 1 0 13708 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1608762545
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_127
timestamp 1608762545
transform 1 0 12788 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 11316 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_110
timestamp 1608762545
transform 1 0 11224 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1608762545
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608762545
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1608762545
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_104
timestamp 1608762545
transform 1 0 10672 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608762545
transform 1 0 8740 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1608762545
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_78
timestamp 1608762545
transform 1 0 8280 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_82
timestamp 1608762545
transform 1 0 8648 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1608762545
transform 1 0 6624 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1608762545
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_56
timestamp 1608762545
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608762545
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 4784 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608762545
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_35
timestamp 1608762545
transform 1 0 4324 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_39
timestamp 1608762545
transform 1 0 4692 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 2484 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1608762545
transform 1 0 1656 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608762545
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1608762545
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608762545
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608762545
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608762545
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608762545
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608762545
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 1608762545
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1608762545
transform 1 0 19964 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1608762545
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1608762545
transform 1 0 19964 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608762545
transform 1 0 19136 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1608762545
transform 1 0 19044 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1608762545
transform 1 0 19504 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_204
timestamp 1608762545
transform 1 0 19872 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 16744 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 18032 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608762545
transform 1 0 18216 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608762545
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1608762545
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_176
timestamp 1608762545
transform 1 0 17296 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1608762545
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 15824 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608762545
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608762545
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_163
timestamp 1608762545
transform 1 0 16100 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1608762545
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 13984 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608762545
transform 1 0 12880 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608762545
transform 1 0 14352 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_6_137
timestamp 1608762545
transform 1 0 13708 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_143
timestamp 1608762545
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_133
timestamp 1608762545
transform 1 0 13340 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_139
timestamp 1608762545
transform 1 0 13892 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608762545
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1608762545
transform 1 0 12512 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1608762545
transform 1 0 11500 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608762545
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1608762545
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_122
timestamp 1608762545
transform 1 0 12328 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_111
timestamp 1608762545
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1608762545
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1608762545
transform 1 0 10488 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1608762545
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1608762545
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608762545
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1608762545
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608762545
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1608762545
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608762545
transform 1 0 7268 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1608762545
transform 1 0 8096 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1608762545
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1608762545
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1608762545
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1608762545
transform 1 0 6072 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608762545
transform 1 0 5244 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1608762545
transform 1 0 5428 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608762545
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_56
timestamp 1608762545
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1608762545
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608762545
transform 1 0 4416 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608762545
transform 1 0 4600 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1608762545
transform 1 0 3036 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608762545
transform 1 0 3772 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608762545
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1608762545
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1608762545
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1608762545
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 1564 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 1472 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608762545
transform 1 0 2944 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608762545
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608762545
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1608762545
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1608762545
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 20516 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608762545
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp 1608762545
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1608762545
transform 1 0 18860 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608762545
transform 1 0 19688 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608762545
transform 1 0 16468 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1608762545
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608762545
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_176
timestamp 1608762545
transform 1 0 17296 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1608762545
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608762545
transform 1 0 15180 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_162
timestamp 1608762545
transform 1 0 16008 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_166
timestamp 1608762545
transform 1 0 16376 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1608762545
transform 1 0 14352 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1608762545
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1608762545
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1608762545
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608762545
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1608762545
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608762545
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_123
timestamp 1608762545
transform 1 0 12420 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608762545
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 10396 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1608762545
transform 1 0 9568 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_85
timestamp 1608762545
transform 1 0 8924 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 7452 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_65
timestamp 1608762545
transform 1 0 7084 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608762545
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1608762545
transform 1 0 5888 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608762545
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_47
timestamp 1608762545
transform 1 0 5428 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_51
timestamp 1608762545
transform 1 0 5796 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 3128 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608762545
transform 1 0 4600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608762545
transform 1 0 1840 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1608762545
transform 1 0 2116 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608762545
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1608762545
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1608762545
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_20
timestamp 1608762545
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608762545
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608762545
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608762545
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608762545
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 19320 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1608762545
transform 1 0 18492 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 17020 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_171
timestamp 1608762545
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1608762545
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608762545
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1608762545
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1608762545
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1608762545
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 13064 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608762545
transform 1 0 12236 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608762545
transform 1 0 11132 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_118
timestamp 1608762545
transform 1 0 11960 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1608762545
transform 1 0 10304 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608762545
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_93
timestamp 1608762545
transform 1 0 9660 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_99
timestamp 1608762545
transform 1 0 10212 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1608762545
transform 1 0 8740 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608762545
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_78
timestamp 1608762545
transform 1 0 8280 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_82
timestamp 1608762545
transform 1 0 8648 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608762545
transform 1 0 6624 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1608762545
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608762545
transform 1 0 4968 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1608762545
transform 1 0 3036 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608762545
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1608762545
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1608762545
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1608762545
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1608762545
transform 1 0 1840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608762545
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1608762545
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1608762545
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1608762545
transform 1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608762545
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1608762545
transform 1 0 20884 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1608762545
transform 1 0 21252 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_203
timestamp 1608762545
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1608762545
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 18308 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608762545
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1608762545
transform 1 0 17204 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608762545
transform 1 0 15180 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608762545
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_156
timestamp 1608762545
transform 1 0 15456 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_164
timestamp 1608762545
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1608762545
transform 1 0 13340 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1608762545
transform 1 0 14352 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_142
timestamp 1608762545
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1608762545
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608762545
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608762545
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608762545
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1608762545
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1608762545
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp 1608762545
transform 1 0 10212 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 8740 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1608762545
transform 1 0 6900 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1608762545
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1608762545
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1608762545
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608762545
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1608762545
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1608762545
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608762545
transform 1 0 4324 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 2852 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1608762545
transform 1 0 2024 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608762545
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1608762545
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1608762545
transform 1 0 1932 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608762545
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608762545
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1608762545
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1608762545
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608762545
transform 1 0 18400 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1608762545
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1608762545
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608762545
transform 1 0 17572 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1608762545
transform 1 0 16744 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_169
timestamp 1608762545
transform 1 0 16652 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608762545
transform 1 0 16284 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608762545
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608762545
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1608762545
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1608762545
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 13432 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608762545
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1608762545
transform 1 0 12604 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608762545
transform 1 0 11500 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_122
timestamp 1608762545
transform 1 0 12328 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608762545
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608762545
transform 1 0 7912 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1608762545
transform 1 0 8740 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 4968 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608762545
transform 1 0 6440 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608762545
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1608762545
transform 1 0 4140 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608762545
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1608762545
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1608762545
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 2024 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608762545
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1608762545
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1608762545
transform 1 0 1932 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608762545
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608762545
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608762545
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1608762545
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608762545
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_209
timestamp 1608762545
transform 1 0 20332 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp 1608762545
transform 1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608762545
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608762545
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608762545
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608762545
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_208
timestamp 1608762545
transform 1 0 20240 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_197
timestamp 1608762545
transform 1 0 19228 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608762545
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608762545
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608762545
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1608762545
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608762545
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608762545
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608762545
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1608762545
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608762545
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608762545
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608762545
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 15916 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608762545
transform 1 0 16192 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 15640 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_160
timestamp 1608762545
transform 1 0 15824 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608762545
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608762545
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1608762545
transform 1 0 14996 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608762545
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1608762545
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_150
timestamp 1608762545
transform 1 0 14904 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608762545
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608762545
transform 1 0 13524 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608762545
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608762545
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608762545
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 14352 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_143
timestamp 1608762545
transform 1 0 14260 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 12420 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608762545
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608762545
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608762545
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115
timestamp 1608762545
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1608762545
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 11224 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 11132 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762545
transform 1 0 8924 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608762545
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1608762545
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762545
transform 1 0 10580 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608762545
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608762545
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762545
transform 1 0 7452 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1608762545
transform 1 0 7452 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1608762545
transform 1 0 8280 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1608762545
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68
timestamp 1608762545
transform 1 0 7360 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1608762545
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608762545
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608762545
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55
timestamp 1608762545
transform 1 0 6164 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1608762545
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1608762545
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_62
timestamp 1608762545
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762545
transform 1 0 4876 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762545
transform 1 0 3036 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1608762545
transform 1 0 4508 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1608762545
transform 1 0 3128 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608762545
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21
timestamp 1608762545
transform 1 0 3036 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1608762545
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36
timestamp 1608762545
transform 1 0 4416 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1608762545
transform 1 0 4508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1608762545
transform 1 0 2208 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608762545
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608762545
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608762545
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15
timestamp 1608762545
transform 1 0 2484 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1608762545
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp 1608762545
transform 1 0 2116 0 1 2720
box -38 -48 130 592
<< labels >>
rlabel metal2 s 18418 22000 18474 22800 4 Test_en_N_out
port 1 nsew
rlabel metal2 s 18878 0 18934 800 4 Test_en_S_in
port 2 nsew
rlabel metal2 s 202 0 258 800 4 bottom_left_grid_pin_42_
port 3 nsew
rlabel metal2 s 570 0 626 800 4 bottom_left_grid_pin_43_
port 4 nsew
rlabel metal2 s 938 0 994 800 4 bottom_left_grid_pin_44_
port 5 nsew
rlabel metal2 s 1306 0 1362 800 4 bottom_left_grid_pin_45_
port 6 nsew
rlabel metal2 s 1674 0 1730 800 4 bottom_left_grid_pin_46_
port 7 nsew
rlabel metal2 s 2042 0 2098 800 4 bottom_left_grid_pin_47_
port 8 nsew
rlabel metal2 s 2410 0 2466 800 4 bottom_left_grid_pin_48_
port 9 nsew
rlabel metal2 s 2778 0 2834 800 4 bottom_left_grid_pin_49_
port 10 nsew
rlabel metal2 s 3146 0 3202 800 4 ccff_head
port 11 nsew
rlabel metal2 s 3514 0 3570 800 4 ccff_tail
port 12 nsew
rlabel metal3 s 0 3272 800 3392 4 chanx_left_in[0]
port 13 nsew
rlabel metal3 s 0 7216 800 7336 4 chanx_left_in[10]
port 14 nsew
rlabel metal3 s 0 7624 800 7744 4 chanx_left_in[11]
port 15 nsew
rlabel metal3 s 0 7896 800 8016 4 chanx_left_in[12]
port 16 nsew
rlabel metal3 s 0 8304 800 8424 4 chanx_left_in[13]
port 17 nsew
rlabel metal3 s 0 8712 800 8832 4 chanx_left_in[14]
port 18 nsew
rlabel metal3 s 0 9120 800 9240 4 chanx_left_in[15]
port 19 nsew
rlabel metal3 s 0 9528 800 9648 4 chanx_left_in[16]
port 20 nsew
rlabel metal3 s 0 9936 800 10056 4 chanx_left_in[17]
port 21 nsew
rlabel metal3 s 0 10344 800 10464 4 chanx_left_in[18]
port 22 nsew
rlabel metal3 s 0 10752 800 10872 4 chanx_left_in[19]
port 23 nsew
rlabel metal3 s 0 3680 800 3800 4 chanx_left_in[1]
port 24 nsew
rlabel metal3 s 0 3952 800 4072 4 chanx_left_in[2]
port 25 nsew
rlabel metal3 s 0 4360 800 4480 4 chanx_left_in[3]
port 26 nsew
rlabel metal3 s 0 4768 800 4888 4 chanx_left_in[4]
port 27 nsew
rlabel metal3 s 0 5176 800 5296 4 chanx_left_in[5]
port 28 nsew
rlabel metal3 s 0 5584 800 5704 4 chanx_left_in[6]
port 29 nsew
rlabel metal3 s 0 5992 800 6112 4 chanx_left_in[7]
port 30 nsew
rlabel metal3 s 0 6400 800 6520 4 chanx_left_in[8]
port 31 nsew
rlabel metal3 s 0 6808 800 6928 4 chanx_left_in[9]
port 32 nsew
rlabel metal3 s 0 11160 800 11280 4 chanx_left_out[0]
port 33 nsew
rlabel metal3 s 0 15104 800 15224 4 chanx_left_out[10]
port 34 nsew
rlabel metal3 s 0 15376 800 15496 4 chanx_left_out[11]
port 35 nsew
rlabel metal3 s 0 15784 800 15904 4 chanx_left_out[12]
port 36 nsew
rlabel metal3 s 0 16192 800 16312 4 chanx_left_out[13]
port 37 nsew
rlabel metal3 s 0 16600 800 16720 4 chanx_left_out[14]
port 38 nsew
rlabel metal3 s 0 17008 800 17128 4 chanx_left_out[15]
port 39 nsew
rlabel metal3 s 0 17416 800 17536 4 chanx_left_out[16]
port 40 nsew
rlabel metal3 s 0 17824 800 17944 4 chanx_left_out[17]
port 41 nsew
rlabel metal3 s 0 18232 800 18352 4 chanx_left_out[18]
port 42 nsew
rlabel metal3 s 0 18640 800 18760 4 chanx_left_out[19]
port 43 nsew
rlabel metal3 s 0 11568 800 11688 4 chanx_left_out[1]
port 44 nsew
rlabel metal3 s 0 11840 800 11960 4 chanx_left_out[2]
port 45 nsew
rlabel metal3 s 0 12248 800 12368 4 chanx_left_out[3]
port 46 nsew
rlabel metal3 s 0 12656 800 12776 4 chanx_left_out[4]
port 47 nsew
rlabel metal3 s 0 13064 800 13184 4 chanx_left_out[5]
port 48 nsew
rlabel metal3 s 0 13472 800 13592 4 chanx_left_out[6]
port 49 nsew
rlabel metal3 s 0 13880 800 14000 4 chanx_left_out[7]
port 50 nsew
rlabel metal3 s 0 14288 800 14408 4 chanx_left_out[8]
port 51 nsew
rlabel metal3 s 0 14696 800 14816 4 chanx_left_out[9]
port 52 nsew
rlabel metal3 s 22000 3272 22800 3392 4 chanx_right_in[0]
port 53 nsew
rlabel metal3 s 22000 7216 22800 7336 4 chanx_right_in[10]
port 54 nsew
rlabel metal3 s 22000 7624 22800 7744 4 chanx_right_in[11]
port 55 nsew
rlabel metal3 s 22000 7896 22800 8016 4 chanx_right_in[12]
port 56 nsew
rlabel metal3 s 22000 8304 22800 8424 4 chanx_right_in[13]
port 57 nsew
rlabel metal3 s 22000 8712 22800 8832 4 chanx_right_in[14]
port 58 nsew
rlabel metal3 s 22000 9120 22800 9240 4 chanx_right_in[15]
port 59 nsew
rlabel metal3 s 22000 9528 22800 9648 4 chanx_right_in[16]
port 60 nsew
rlabel metal3 s 22000 9936 22800 10056 4 chanx_right_in[17]
port 61 nsew
rlabel metal3 s 22000 10344 22800 10464 4 chanx_right_in[18]
port 62 nsew
rlabel metal3 s 22000 10752 22800 10872 4 chanx_right_in[19]
port 63 nsew
rlabel metal3 s 22000 3680 22800 3800 4 chanx_right_in[1]
port 64 nsew
rlabel metal3 s 22000 3952 22800 4072 4 chanx_right_in[2]
port 65 nsew
rlabel metal3 s 22000 4360 22800 4480 4 chanx_right_in[3]
port 66 nsew
rlabel metal3 s 22000 4768 22800 4888 4 chanx_right_in[4]
port 67 nsew
rlabel metal3 s 22000 5176 22800 5296 4 chanx_right_in[5]
port 68 nsew
rlabel metal3 s 22000 5584 22800 5704 4 chanx_right_in[6]
port 69 nsew
rlabel metal3 s 22000 5992 22800 6112 4 chanx_right_in[7]
port 70 nsew
rlabel metal3 s 22000 6400 22800 6520 4 chanx_right_in[8]
port 71 nsew
rlabel metal3 s 22000 6808 22800 6928 4 chanx_right_in[9]
port 72 nsew
rlabel metal3 s 22000 11160 22800 11280 4 chanx_right_out[0]
port 73 nsew
rlabel metal3 s 22000 15104 22800 15224 4 chanx_right_out[10]
port 74 nsew
rlabel metal3 s 22000 15376 22800 15496 4 chanx_right_out[11]
port 75 nsew
rlabel metal3 s 22000 15784 22800 15904 4 chanx_right_out[12]
port 76 nsew
rlabel metal3 s 22000 16192 22800 16312 4 chanx_right_out[13]
port 77 nsew
rlabel metal3 s 22000 16600 22800 16720 4 chanx_right_out[14]
port 78 nsew
rlabel metal3 s 22000 17008 22800 17128 4 chanx_right_out[15]
port 79 nsew
rlabel metal3 s 22000 17416 22800 17536 4 chanx_right_out[16]
port 80 nsew
rlabel metal3 s 22000 17824 22800 17944 4 chanx_right_out[17]
port 81 nsew
rlabel metal3 s 22000 18232 22800 18352 4 chanx_right_out[18]
port 82 nsew
rlabel metal3 s 22000 18640 22800 18760 4 chanx_right_out[19]
port 83 nsew
rlabel metal3 s 22000 11568 22800 11688 4 chanx_right_out[1]
port 84 nsew
rlabel metal3 s 22000 11840 22800 11960 4 chanx_right_out[2]
port 85 nsew
rlabel metal3 s 22000 12248 22800 12368 4 chanx_right_out[3]
port 86 nsew
rlabel metal3 s 22000 12656 22800 12776 4 chanx_right_out[4]
port 87 nsew
rlabel metal3 s 22000 13064 22800 13184 4 chanx_right_out[5]
port 88 nsew
rlabel metal3 s 22000 13472 22800 13592 4 chanx_right_out[6]
port 89 nsew
rlabel metal3 s 22000 13880 22800 14000 4 chanx_right_out[7]
port 90 nsew
rlabel metal3 s 22000 14288 22800 14408 4 chanx_right_out[8]
port 91 nsew
rlabel metal3 s 22000 14696 22800 14816 4 chanx_right_out[9]
port 92 nsew
rlabel metal2 s 3882 0 3938 800 4 chany_bottom_in[0]
port 93 nsew
rlabel metal2 s 7654 0 7710 800 4 chany_bottom_in[10]
port 94 nsew
rlabel metal2 s 8022 0 8078 800 4 chany_bottom_in[11]
port 95 nsew
rlabel metal2 s 8390 0 8446 800 4 chany_bottom_in[12]
port 96 nsew
rlabel metal2 s 8758 0 8814 800 4 chany_bottom_in[13]
port 97 nsew
rlabel metal2 s 9126 0 9182 800 4 chany_bottom_in[14]
port 98 nsew
rlabel metal2 s 9494 0 9550 800 4 chany_bottom_in[15]
port 99 nsew
rlabel metal2 s 9862 0 9918 800 4 chany_bottom_in[16]
port 100 nsew
rlabel metal2 s 10230 0 10286 800 4 chany_bottom_in[17]
port 101 nsew
rlabel metal2 s 10598 0 10654 800 4 chany_bottom_in[18]
port 102 nsew
rlabel metal2 s 10966 0 11022 800 4 chany_bottom_in[19]
port 103 nsew
rlabel metal2 s 4250 0 4306 800 4 chany_bottom_in[1]
port 104 nsew
rlabel metal2 s 4618 0 4674 800 4 chany_bottom_in[2]
port 105 nsew
rlabel metal2 s 4986 0 5042 800 4 chany_bottom_in[3]
port 106 nsew
rlabel metal2 s 5354 0 5410 800 4 chany_bottom_in[4]
port 107 nsew
rlabel metal2 s 5722 0 5778 800 4 chany_bottom_in[5]
port 108 nsew
rlabel metal2 s 6182 0 6238 800 4 chany_bottom_in[6]
port 109 nsew
rlabel metal2 s 6550 0 6606 800 4 chany_bottom_in[7]
port 110 nsew
rlabel metal2 s 6918 0 6974 800 4 chany_bottom_in[8]
port 111 nsew
rlabel metal2 s 7286 0 7342 800 4 chany_bottom_in[9]
port 112 nsew
rlabel metal2 s 11334 0 11390 800 4 chany_bottom_out[0]
port 113 nsew
rlabel metal2 s 15106 0 15162 800 4 chany_bottom_out[10]
port 114 nsew
rlabel metal2 s 15474 0 15530 800 4 chany_bottom_out[11]
port 115 nsew
rlabel metal2 s 15842 0 15898 800 4 chany_bottom_out[12]
port 116 nsew
rlabel metal2 s 16210 0 16266 800 4 chany_bottom_out[13]
port 117 nsew
rlabel metal2 s 16578 0 16634 800 4 chany_bottom_out[14]
port 118 nsew
rlabel metal2 s 16946 0 17002 800 4 chany_bottom_out[15]
port 119 nsew
rlabel metal2 s 17406 0 17462 800 4 chany_bottom_out[16]
port 120 nsew
rlabel metal2 s 17774 0 17830 800 4 chany_bottom_out[17]
port 121 nsew
rlabel metal2 s 18142 0 18198 800 4 chany_bottom_out[18]
port 122 nsew
rlabel metal2 s 18510 0 18566 800 4 chany_bottom_out[19]
port 123 nsew
rlabel metal2 s 11794 0 11850 800 4 chany_bottom_out[1]
port 124 nsew
rlabel metal2 s 12162 0 12218 800 4 chany_bottom_out[2]
port 125 nsew
rlabel metal2 s 12530 0 12586 800 4 chany_bottom_out[3]
port 126 nsew
rlabel metal2 s 12898 0 12954 800 4 chany_bottom_out[4]
port 127 nsew
rlabel metal2 s 13266 0 13322 800 4 chany_bottom_out[5]
port 128 nsew
rlabel metal2 s 13634 0 13690 800 4 chany_bottom_out[6]
port 129 nsew
rlabel metal2 s 14002 0 14058 800 4 chany_bottom_out[7]
port 130 nsew
rlabel metal2 s 14370 0 14426 800 4 chany_bottom_out[8]
port 131 nsew
rlabel metal2 s 14738 0 14794 800 4 chany_bottom_out[9]
port 132 nsew
rlabel metal2 s 3238 22000 3294 22800 4 chany_top_in[0]
port 133 nsew
rlabel metal2 s 7010 22000 7066 22800 4 chany_top_in[10]
port 134 nsew
rlabel metal2 s 7378 22000 7434 22800 4 chany_top_in[11]
port 135 nsew
rlabel metal2 s 7746 22000 7802 22800 4 chany_top_in[12]
port 136 nsew
rlabel metal2 s 8114 22000 8170 22800 4 chany_top_in[13]
port 137 nsew
rlabel metal2 s 8482 22000 8538 22800 4 chany_top_in[14]
port 138 nsew
rlabel metal2 s 8942 22000 8998 22800 4 chany_top_in[15]
port 139 nsew
rlabel metal2 s 9310 22000 9366 22800 4 chany_top_in[16]
port 140 nsew
rlabel metal2 s 9678 22000 9734 22800 4 chany_top_in[17]
port 141 nsew
rlabel metal2 s 10046 22000 10102 22800 4 chany_top_in[18]
port 142 nsew
rlabel metal2 s 10414 22000 10470 22800 4 chany_top_in[19]
port 143 nsew
rlabel metal2 s 3606 22000 3662 22800 4 chany_top_in[1]
port 144 nsew
rlabel metal2 s 3974 22000 4030 22800 4 chany_top_in[2]
port 145 nsew
rlabel metal2 s 4342 22000 4398 22800 4 chany_top_in[3]
port 146 nsew
rlabel metal2 s 4710 22000 4766 22800 4 chany_top_in[4]
port 147 nsew
rlabel metal2 s 5078 22000 5134 22800 4 chany_top_in[5]
port 148 nsew
rlabel metal2 s 5446 22000 5502 22800 4 chany_top_in[6]
port 149 nsew
rlabel metal2 s 5906 22000 5962 22800 4 chany_top_in[7]
port 150 nsew
rlabel metal2 s 6274 22000 6330 22800 4 chany_top_in[8]
port 151 nsew
rlabel metal2 s 6642 22000 6698 22800 4 chany_top_in[9]
port 152 nsew
rlabel metal2 s 10782 22000 10838 22800 4 chany_top_out[0]
port 153 nsew
rlabel metal2 s 14646 22000 14702 22800 4 chany_top_out[10]
port 154 nsew
rlabel metal2 s 15014 22000 15070 22800 4 chany_top_out[11]
port 155 nsew
rlabel metal2 s 15382 22000 15438 22800 4 chany_top_out[12]
port 156 nsew
rlabel metal2 s 15750 22000 15806 22800 4 chany_top_out[13]
port 157 nsew
rlabel metal2 s 16118 22000 16174 22800 4 chany_top_out[14]
port 158 nsew
rlabel metal2 s 16486 22000 16542 22800 4 chany_top_out[15]
port 159 nsew
rlabel metal2 s 16854 22000 16910 22800 4 chany_top_out[16]
port 160 nsew
rlabel metal2 s 17314 22000 17370 22800 4 chany_top_out[17]
port 161 nsew
rlabel metal2 s 17682 22000 17738 22800 4 chany_top_out[18]
port 162 nsew
rlabel metal2 s 18050 22000 18106 22800 4 chany_top_out[19]
port 163 nsew
rlabel metal2 s 11150 22000 11206 22800 4 chany_top_out[1]
port 164 nsew
rlabel metal2 s 11610 22000 11666 22800 4 chany_top_out[2]
port 165 nsew
rlabel metal2 s 11978 22000 12034 22800 4 chany_top_out[3]
port 166 nsew
rlabel metal2 s 12346 22000 12402 22800 4 chany_top_out[4]
port 167 nsew
rlabel metal2 s 12714 22000 12770 22800 4 chany_top_out[5]
port 168 nsew
rlabel metal2 s 13082 22000 13138 22800 4 chany_top_out[6]
port 169 nsew
rlabel metal2 s 13450 22000 13506 22800 4 chany_top_out[7]
port 170 nsew
rlabel metal2 s 13818 22000 13874 22800 4 chany_top_out[8]
port 171 nsew
rlabel metal2 s 14186 22000 14242 22800 4 chany_top_out[9]
port 172 nsew
rlabel metal3 s 22000 20544 22800 20664 4 clk_1_E_out
port 173 nsew
rlabel metal2 s 18786 22000 18842 22800 4 clk_1_N_in
port 174 nsew
rlabel metal2 s 19246 0 19302 800 4 clk_1_S_in
port 175 nsew
rlabel metal3 s 0 19048 800 19168 4 clk_1_W_out
port 176 nsew
rlabel metal3 s 22000 19048 22800 19168 4 clk_2_E_in
port 177 nsew
rlabel metal3 s 22000 20952 22800 21072 4 clk_2_E_out
port 178 nsew
rlabel metal2 s 19154 22000 19210 22800 4 clk_2_N_in
port 179 nsew
rlabel metal2 s 21454 22000 21510 22800 4 clk_2_N_out
port 180 nsew
rlabel metal2 s 19614 0 19670 800 4 clk_2_S_in
port 181 nsew
rlabel metal2 s 20350 0 20406 800 4 clk_2_S_out
port 182 nsew
rlabel metal3 s 0 21360 800 21480 4 clk_2_W_in
port 183 nsew
rlabel metal3 s 0 19320 800 19440 4 clk_2_W_out
port 184 nsew
rlabel metal3 s 22000 19320 22800 19440 4 clk_3_E_in
port 185 nsew
rlabel metal3 s 22000 21360 22800 21480 4 clk_3_E_out
port 186 nsew
rlabel metal2 s 19522 22000 19578 22800 4 clk_3_N_in
port 187 nsew
rlabel metal2 s 21822 22000 21878 22800 4 clk_3_N_out
port 188 nsew
rlabel metal2 s 19982 0 20038 800 4 clk_3_S_in
port 189 nsew
rlabel metal2 s 20718 0 20774 800 4 clk_3_S_out
port 190 nsew
rlabel metal3 s 0 21768 800 21888 4 clk_3_W_in
port 191 nsew
rlabel metal3 s 0 19728 800 19848 4 clk_3_W_out
port 192 nsew
rlabel metal3 s 0 144 800 264 4 left_bottom_grid_pin_34_
port 193 nsew
rlabel metal3 s 0 416 800 536 4 left_bottom_grid_pin_35_
port 194 nsew
rlabel metal3 s 0 824 800 944 4 left_bottom_grid_pin_36_
port 195 nsew
rlabel metal3 s 0 1232 800 1352 4 left_bottom_grid_pin_37_
port 196 nsew
rlabel metal3 s 0 1640 800 1760 4 left_bottom_grid_pin_38_
port 197 nsew
rlabel metal3 s 0 2048 800 2168 4 left_bottom_grid_pin_39_
port 198 nsew
rlabel metal3 s 0 2456 800 2576 4 left_bottom_grid_pin_40_
port 199 nsew
rlabel metal3 s 0 2864 800 2984 4 left_bottom_grid_pin_41_
port 200 nsew
rlabel metal2 s 19890 22000 19946 22800 4 prog_clk_0_N_in
port 201 nsew
rlabel metal3 s 22000 21768 22800 21888 4 prog_clk_1_E_out
port 202 nsew
rlabel metal2 s 20350 22000 20406 22800 4 prog_clk_1_N_in
port 203 nsew
rlabel metal2 s 21086 0 21142 800 4 prog_clk_1_S_in
port 204 nsew
rlabel metal3 s 0 20136 800 20256 4 prog_clk_1_W_out
port 205 nsew
rlabel metal3 s 22000 19728 22800 19848 4 prog_clk_2_E_in
port 206 nsew
rlabel metal3 s 22000 22176 22800 22296 4 prog_clk_2_E_out
port 207 nsew
rlabel metal2 s 20718 22000 20774 22800 4 prog_clk_2_N_in
port 208 nsew
rlabel metal2 s 22190 22000 22246 22800 4 prog_clk_2_N_out
port 209 nsew
rlabel metal2 s 21454 0 21510 800 4 prog_clk_2_S_in
port 210 nsew
rlabel metal2 s 22190 0 22246 800 4 prog_clk_2_S_out
port 211 nsew
rlabel metal3 s 0 22176 800 22296 4 prog_clk_2_W_in
port 212 nsew
rlabel metal3 s 0 20544 800 20664 4 prog_clk_2_W_out
port 213 nsew
rlabel metal3 s 22000 20136 22800 20256 4 prog_clk_3_E_in
port 214 nsew
rlabel metal3 s 22000 22584 22800 22704 4 prog_clk_3_E_out
port 215 nsew
rlabel metal2 s 21086 22000 21142 22800 4 prog_clk_3_N_in
port 216 nsew
rlabel metal2 s 22558 22000 22614 22800 4 prog_clk_3_N_out
port 217 nsew
rlabel metal2 s 21822 0 21878 800 4 prog_clk_3_S_in
port 218 nsew
rlabel metal2 s 22558 0 22614 800 4 prog_clk_3_S_out
port 219 nsew
rlabel metal3 s 0 22584 800 22704 4 prog_clk_3_W_in
port 220 nsew
rlabel metal3 s 0 20952 800 21072 4 prog_clk_3_W_out
port 221 nsew
rlabel metal3 s 22000 144 22800 264 4 right_bottom_grid_pin_34_
port 222 nsew
rlabel metal3 s 22000 416 22800 536 4 right_bottom_grid_pin_35_
port 223 nsew
rlabel metal3 s 22000 824 22800 944 4 right_bottom_grid_pin_36_
port 224 nsew
rlabel metal3 s 22000 1232 22800 1352 4 right_bottom_grid_pin_37_
port 225 nsew
rlabel metal3 s 22000 1640 22800 1760 4 right_bottom_grid_pin_38_
port 226 nsew
rlabel metal3 s 22000 2048 22800 2168 4 right_bottom_grid_pin_39_
port 227 nsew
rlabel metal3 s 22000 2456 22800 2576 4 right_bottom_grid_pin_40_
port 228 nsew
rlabel metal3 s 22000 2864 22800 2984 4 right_bottom_grid_pin_41_
port 229 nsew
rlabel metal2 s 202 22000 258 22800 4 top_left_grid_pin_42_
port 230 nsew
rlabel metal2 s 570 22000 626 22800 4 top_left_grid_pin_43_
port 231 nsew
rlabel metal2 s 938 22000 994 22800 4 top_left_grid_pin_44_
port 232 nsew
rlabel metal2 s 1306 22000 1362 22800 4 top_left_grid_pin_45_
port 233 nsew
rlabel metal2 s 1674 22000 1730 22800 4 top_left_grid_pin_46_
port 234 nsew
rlabel metal2 s 2042 22000 2098 22800 4 top_left_grid_pin_47_
port 235 nsew
rlabel metal2 s 2410 22000 2466 22800 4 top_left_grid_pin_48_
port 236 nsew
rlabel metal2 s 2778 22000 2834 22800 4 top_left_grid_pin_49_
port 237 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 238 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 239 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22800
string GDS_FILE /ef/openfpga/openlane/runs/sb_1__1_/results/magic/sb_1__1_.gds
string GDS_END 1788730
string GDS_START 81916
<< end >>
