magic
tech sky130A
magscale 1 2
timestamp 1605121875
<< locali >>
rect 21649 20247 21683 20349
rect 14289 19159 14323 19397
rect 20637 16983 20671 17085
rect 24869 16439 24903 16677
rect 16681 14399 16715 14569
rect 18705 12087 18739 12257
rect 12265 11611 12299 11849
rect 14289 9571 14323 9673
rect 23489 8959 23523 9129
rect 13093 2499 13127 2601
<< viali >>
rect 16681 25449 16715 25483
rect 19073 25449 19107 25483
rect 22109 25449 22143 25483
rect 14289 25313 14323 25347
rect 16497 25313 16531 25347
rect 18889 25313 18923 25347
rect 19993 25313 20027 25347
rect 21925 25313 21959 25347
rect 24593 25313 24627 25347
rect 15485 25245 15519 25279
rect 14473 25177 14507 25211
rect 20177 25177 20211 25211
rect 24777 25109 24811 25143
rect 20637 24905 20671 24939
rect 16865 24769 16899 24803
rect 13553 24701 13587 24735
rect 14657 24701 14691 24735
rect 15393 24701 15427 24735
rect 15945 24701 15979 24735
rect 18061 24701 18095 24735
rect 19349 24701 19383 24735
rect 20453 24701 20487 24735
rect 21005 24701 21039 24735
rect 21557 24701 21591 24735
rect 22201 24701 22235 24735
rect 24593 24701 24627 24735
rect 25145 24701 25179 24735
rect 14933 24633 14967 24667
rect 13461 24565 13495 24599
rect 13737 24565 13771 24599
rect 14289 24565 14323 24599
rect 16129 24565 16163 24599
rect 16589 24565 16623 24599
rect 17785 24565 17819 24599
rect 18245 24565 18279 24599
rect 18981 24565 19015 24599
rect 19533 24565 19567 24599
rect 19993 24565 20027 24599
rect 21741 24565 21775 24599
rect 22569 24565 22603 24599
rect 24409 24565 24443 24599
rect 24777 24565 24811 24599
rect 12817 24361 12851 24395
rect 14013 24361 14047 24395
rect 15485 24361 15519 24395
rect 16221 24361 16255 24395
rect 18153 24361 18187 24395
rect 18889 24361 18923 24395
rect 21097 24361 21131 24395
rect 22569 24361 22603 24395
rect 23673 24361 23707 24395
rect 16742 24293 16776 24327
rect 12633 24225 12667 24259
rect 13829 24225 13863 24259
rect 14381 24225 14415 24259
rect 15301 24225 15335 24259
rect 18705 24225 18739 24259
rect 20913 24225 20947 24259
rect 22385 24225 22419 24259
rect 23489 24225 23523 24259
rect 24593 24225 24627 24259
rect 14841 24157 14875 24191
rect 16497 24157 16531 24191
rect 19809 24157 19843 24191
rect 17877 24089 17911 24123
rect 12541 24021 12575 24055
rect 15853 24021 15887 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 24777 24021 24811 24055
rect 12173 23817 12207 23851
rect 13461 23817 13495 23851
rect 16037 23817 16071 23851
rect 19809 23817 19843 23851
rect 21557 23817 21591 23851
rect 22661 23817 22695 23851
rect 23489 23817 23523 23851
rect 13001 23681 13035 23715
rect 15761 23681 15795 23715
rect 16773 23681 16807 23715
rect 17233 23681 17267 23715
rect 18613 23681 18647 23715
rect 20913 23681 20947 23715
rect 23857 23681 23891 23715
rect 12817 23613 12851 23647
rect 14013 23613 14047 23647
rect 16589 23613 16623 23647
rect 18429 23613 18463 23647
rect 19625 23613 19659 23647
rect 20177 23613 20211 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 22477 23613 22511 23647
rect 23673 23613 23707 23647
rect 24961 23613 24995 23647
rect 12909 23545 12943 23579
rect 13921 23545 13955 23579
rect 14280 23545 14314 23579
rect 16681 23545 16715 23579
rect 18521 23545 18555 23579
rect 12449 23477 12483 23511
rect 15393 23477 15427 23511
rect 16221 23477 16255 23511
rect 17785 23477 17819 23511
rect 18061 23477 18095 23511
rect 19073 23477 19107 23511
rect 19533 23477 19567 23511
rect 22385 23477 22419 23511
rect 23029 23477 23063 23511
rect 24593 23477 24627 23511
rect 25145 23477 25179 23511
rect 25513 23477 25547 23511
rect 12449 23273 12483 23307
rect 12909 23273 12943 23307
rect 15025 23273 15059 23307
rect 16957 23273 16991 23307
rect 21281 23273 21315 23307
rect 22753 23273 22787 23307
rect 13246 23205 13280 23239
rect 17325 23205 17359 23239
rect 17868 23205 17902 23239
rect 25237 23205 25271 23239
rect 15301 23137 15335 23171
rect 15568 23137 15602 23171
rect 17601 23137 17635 23171
rect 19349 23137 19383 23171
rect 19717 23137 19751 23171
rect 20361 23137 20395 23171
rect 22569 23137 22603 23171
rect 23673 23137 23707 23171
rect 24961 23137 24995 23171
rect 11989 23069 12023 23103
rect 13001 23069 13035 23103
rect 19809 23069 19843 23103
rect 21373 23069 21407 23103
rect 21465 23069 21499 23103
rect 22477 23069 22511 23103
rect 23857 23069 23891 23103
rect 16681 23001 16715 23035
rect 21925 23001 21959 23035
rect 14381 22933 14415 22967
rect 14657 22933 14691 22967
rect 18981 22933 19015 22967
rect 20637 22933 20671 22967
rect 20913 22933 20947 22967
rect 14657 22729 14691 22763
rect 17693 22729 17727 22763
rect 21005 22729 21039 22763
rect 24869 22729 24903 22763
rect 11897 22593 11931 22627
rect 12449 22593 12483 22627
rect 14565 22593 14599 22627
rect 15209 22593 15243 22627
rect 15669 22593 15703 22627
rect 16865 22593 16899 22627
rect 17049 22593 17083 22627
rect 18337 22593 18371 22627
rect 23949 22593 23983 22627
rect 18797 22525 18831 22559
rect 18981 22525 19015 22559
rect 21189 22525 21223 22559
rect 22845 22525 22879 22559
rect 23673 22525 23707 22559
rect 24961 22525 24995 22559
rect 25513 22525 25547 22559
rect 12694 22457 12728 22491
rect 14197 22457 14231 22491
rect 15025 22457 15059 22491
rect 16313 22457 16347 22491
rect 16773 22457 16807 22491
rect 19226 22457 19260 22491
rect 21434 22457 21468 22491
rect 12265 22389 12299 22423
rect 13829 22389 13863 22423
rect 15117 22389 15151 22423
rect 16405 22389 16439 22423
rect 20361 22389 20395 22423
rect 22569 22389 22603 22423
rect 23489 22389 23523 22423
rect 24409 22389 24443 22423
rect 25145 22389 25179 22423
rect 10885 22185 10919 22219
rect 12357 22185 12391 22219
rect 13001 22185 13035 22219
rect 13645 22185 13679 22219
rect 16773 22185 16807 22219
rect 18061 22185 18095 22219
rect 20729 22185 20763 22219
rect 14013 22117 14047 22151
rect 10977 22049 11011 22083
rect 11244 22049 11278 22083
rect 13461 22049 13495 22083
rect 14657 22049 14691 22083
rect 16037 22049 16071 22083
rect 17601 22049 17635 22083
rect 18153 22049 18187 22083
rect 19625 22049 19659 22083
rect 20361 22049 20395 22083
rect 21364 22049 21398 22083
rect 23857 22049 23891 22083
rect 24133 22049 24167 22083
rect 25145 22049 25179 22083
rect 25421 22049 25455 22083
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 16129 21981 16163 22015
rect 16313 21981 16347 22015
rect 18245 21981 18279 22015
rect 19717 21981 19751 22015
rect 19809 21981 19843 22015
rect 21097 21981 21131 22015
rect 15117 21913 15151 21947
rect 17693 21913 17727 21947
rect 10333 21845 10367 21879
rect 15577 21845 15611 21879
rect 15669 21845 15703 21879
rect 18705 21845 18739 21879
rect 19073 21845 19107 21879
rect 19257 21845 19291 21879
rect 22477 21845 22511 21879
rect 22753 21845 22787 21879
rect 10057 21641 10091 21675
rect 11253 21641 11287 21675
rect 14197 21641 14231 21675
rect 15301 21641 15335 21675
rect 15669 21641 15703 21675
rect 17509 21641 17543 21675
rect 19717 21641 19751 21675
rect 23857 21641 23891 21675
rect 10241 21573 10275 21607
rect 20453 21573 20487 21607
rect 21465 21573 21499 21607
rect 25145 21573 25179 21607
rect 10793 21505 10827 21539
rect 12265 21505 12299 21539
rect 13001 21505 13035 21539
rect 14749 21505 14783 21539
rect 16313 21505 16347 21539
rect 16497 21505 16531 21539
rect 18889 21505 18923 21539
rect 19441 21505 19475 21539
rect 20361 21505 20395 21539
rect 21097 21505 21131 21539
rect 22569 21505 22603 21539
rect 23029 21505 23063 21539
rect 10609 21437 10643 21471
rect 14565 21437 14599 21471
rect 20821 21437 20855 21471
rect 23489 21437 23523 21471
rect 24225 21437 24259 21471
rect 25513 21437 25547 21471
rect 26065 21437 26099 21471
rect 12817 21369 12851 21403
rect 17877 21369 17911 21403
rect 18797 21369 18831 21403
rect 21833 21369 21867 21403
rect 22477 21369 22511 21403
rect 24501 21369 24535 21403
rect 10701 21301 10735 21335
rect 11805 21301 11839 21335
rect 12449 21301 12483 21335
rect 12909 21301 12943 21335
rect 13645 21301 13679 21335
rect 14013 21301 14047 21335
rect 14657 21301 14691 21335
rect 15853 21301 15887 21335
rect 16221 21301 16255 21335
rect 16957 21301 16991 21335
rect 18337 21301 18371 21335
rect 18705 21301 18739 21335
rect 20913 21301 20947 21335
rect 22017 21301 22051 21335
rect 22385 21301 22419 21335
rect 25697 21301 25731 21335
rect 11897 21097 11931 21131
rect 12541 21097 12575 21131
rect 12725 21097 12759 21131
rect 13185 21097 13219 21131
rect 13829 21097 13863 21131
rect 14749 21097 14783 21131
rect 17785 21097 17819 21131
rect 19349 21097 19383 21131
rect 19901 21097 19935 21131
rect 20453 21097 20487 21131
rect 21189 21097 21223 21131
rect 24041 21097 24075 21131
rect 10762 21029 10796 21063
rect 10517 20961 10551 20995
rect 13093 20961 13127 20995
rect 14473 20961 14507 20995
rect 15761 20961 15795 20995
rect 16120 20961 16154 20995
rect 18429 20961 18463 20995
rect 19717 20961 19751 20995
rect 21465 20961 21499 20995
rect 21732 20961 21766 20995
rect 25237 20961 25271 20995
rect 13277 20893 13311 20927
rect 15853 20893 15887 20927
rect 18521 20893 18555 20927
rect 18705 20893 18739 20927
rect 24133 20893 24167 20927
rect 24225 20893 24259 20927
rect 14289 20825 14323 20859
rect 22845 20825 22879 20859
rect 23673 20825 23707 20859
rect 10333 20757 10367 20791
rect 14105 20757 14139 20791
rect 17233 20757 17267 20791
rect 18061 20757 18095 20791
rect 23121 20757 23155 20791
rect 23489 20757 23523 20791
rect 25421 20757 25455 20791
rect 9413 20553 9447 20587
rect 10793 20553 10827 20587
rect 11805 20553 11839 20587
rect 15577 20553 15611 20587
rect 17509 20553 17543 20587
rect 18245 20553 18279 20587
rect 21373 20553 21407 20587
rect 22017 20553 22051 20587
rect 25053 20553 25087 20587
rect 25973 20553 26007 20587
rect 17049 20485 17083 20519
rect 23489 20485 23523 20519
rect 9781 20417 9815 20451
rect 11345 20417 11379 20451
rect 12173 20417 12207 20451
rect 13277 20417 13311 20451
rect 13645 20417 13679 20451
rect 16497 20417 16531 20451
rect 16589 20417 16623 20451
rect 20913 20417 20947 20451
rect 21189 20417 21223 20451
rect 22569 20417 22603 20451
rect 24133 20417 24167 20451
rect 24225 20417 24259 20451
rect 25421 20417 25455 20451
rect 9505 20349 9539 20383
rect 13912 20349 13946 20383
rect 15945 20349 15979 20383
rect 18061 20349 18095 20383
rect 19165 20349 19199 20383
rect 21557 20349 21591 20383
rect 21649 20349 21683 20383
rect 22477 20349 22511 20383
rect 24685 20349 24719 20383
rect 25237 20349 25271 20383
rect 10333 20281 10367 20315
rect 11161 20281 11195 20315
rect 12449 20281 12483 20315
rect 19073 20281 19107 20315
rect 19410 20281 19444 20315
rect 24041 20281 24075 20315
rect 10609 20213 10643 20247
rect 11253 20213 11287 20247
rect 13001 20213 13035 20247
rect 15025 20213 15059 20247
rect 16037 20213 16071 20247
rect 16405 20213 16439 20247
rect 17785 20213 17819 20247
rect 18705 20213 18739 20247
rect 20545 20213 20579 20247
rect 21649 20213 21683 20247
rect 21833 20213 21867 20247
rect 22385 20213 22419 20247
rect 23029 20213 23063 20247
rect 23673 20213 23707 20247
rect 11529 20009 11563 20043
rect 12817 20009 12851 20043
rect 15025 20009 15059 20043
rect 17233 20009 17267 20043
rect 17785 20009 17819 20043
rect 18153 20009 18187 20043
rect 18245 20009 18279 20043
rect 18889 20009 18923 20043
rect 19901 20009 19935 20043
rect 20361 20009 20395 20043
rect 20729 20009 20763 20043
rect 21373 20009 21407 20043
rect 23673 20009 23707 20043
rect 24317 20009 24351 20043
rect 25513 20009 25547 20043
rect 10057 19941 10091 19975
rect 12081 19941 12115 19975
rect 12449 19941 12483 19975
rect 17601 19941 17635 19975
rect 24869 19941 24903 19975
rect 10149 19873 10183 19907
rect 10405 19873 10439 19907
rect 13165 19873 13199 19907
rect 15577 19873 15611 19907
rect 15833 19873 15867 19907
rect 19717 19873 19751 19907
rect 21189 19873 21223 19907
rect 22560 19873 22594 19907
rect 24041 19873 24075 19907
rect 24961 19873 24995 19907
rect 12909 19805 12943 19839
rect 18337 19805 18371 19839
rect 19625 19805 19659 19839
rect 22293 19805 22327 19839
rect 25053 19805 25087 19839
rect 14657 19737 14691 19771
rect 16957 19737 16991 19771
rect 24501 19737 24535 19771
rect 14289 19669 14323 19703
rect 19257 19669 19291 19703
rect 22109 19669 22143 19703
rect 10609 19465 10643 19499
rect 11805 19465 11839 19499
rect 12265 19465 12299 19499
rect 14105 19465 14139 19499
rect 18521 19465 18555 19499
rect 21925 19465 21959 19499
rect 24777 19465 24811 19499
rect 25973 19465 26007 19499
rect 14289 19397 14323 19431
rect 17509 19397 17543 19431
rect 23673 19397 23707 19431
rect 12449 19329 12483 19363
rect 10241 19261 10275 19295
rect 12694 19193 12728 19227
rect 15209 19329 15243 19363
rect 17049 19329 17083 19363
rect 19165 19329 19199 19363
rect 22569 19329 22603 19363
rect 24225 19329 24259 19363
rect 14473 19261 14507 19295
rect 15117 19261 15151 19295
rect 15945 19261 15979 19295
rect 16773 19261 16807 19295
rect 18061 19261 18095 19295
rect 20913 19261 20947 19295
rect 23489 19261 23523 19295
rect 24133 19261 24167 19295
rect 25237 19261 25271 19295
rect 15025 19193 15059 19227
rect 17785 19193 17819 19227
rect 19410 19193 19444 19227
rect 22385 19193 22419 19227
rect 25513 19193 25547 19227
rect 11345 19125 11379 19159
rect 13829 19125 13863 19159
rect 14289 19125 14323 19159
rect 14657 19125 14691 19159
rect 16221 19125 16255 19159
rect 16405 19125 16439 19159
rect 16865 19125 16899 19159
rect 18981 19125 19015 19159
rect 20545 19125 20579 19159
rect 21281 19125 21315 19159
rect 22017 19125 22051 19159
rect 22477 19125 22511 19159
rect 23121 19125 23155 19159
rect 24041 19125 24075 19159
rect 25145 19125 25179 19159
rect 14381 18921 14415 18955
rect 14565 18921 14599 18955
rect 15669 18921 15703 18955
rect 17141 18921 17175 18955
rect 17877 18921 17911 18955
rect 19809 18921 19843 18955
rect 20729 18921 20763 18955
rect 21373 18921 21407 18955
rect 22109 18921 22143 18955
rect 23673 18921 23707 18955
rect 25513 18921 25547 18955
rect 13461 18853 13495 18887
rect 24869 18853 24903 18887
rect 11805 18785 11839 18819
rect 13369 18785 13403 18819
rect 14749 18785 14783 18819
rect 16497 18785 16531 18819
rect 18429 18785 18463 18819
rect 18685 18785 18719 18819
rect 21189 18785 21223 18819
rect 22549 18785 22583 18819
rect 23949 18785 23983 18819
rect 24317 18785 24351 18819
rect 11897 18717 11931 18751
rect 12081 18717 12115 18751
rect 13645 18717 13679 18751
rect 16589 18717 16623 18751
rect 16681 18717 16715 18751
rect 22293 18717 22327 18751
rect 24961 18717 24995 18751
rect 25145 18717 25179 18751
rect 11437 18649 11471 18683
rect 12541 18649 12575 18683
rect 24501 18649 24535 18683
rect 12909 18581 12943 18615
rect 13001 18581 13035 18615
rect 14013 18581 14047 18615
rect 15117 18581 15151 18615
rect 15945 18581 15979 18615
rect 16129 18581 16163 18615
rect 18153 18581 18187 18615
rect 20085 18581 20119 18615
rect 12725 18377 12759 18411
rect 13921 18377 13955 18411
rect 14197 18377 14231 18411
rect 14841 18377 14875 18411
rect 19073 18377 19107 18411
rect 20637 18377 20671 18411
rect 22385 18377 22419 18411
rect 22661 18377 22695 18411
rect 23673 18377 23707 18411
rect 24685 18377 24719 18411
rect 11805 18309 11839 18343
rect 12817 18309 12851 18343
rect 19257 18309 19291 18343
rect 20821 18309 20855 18343
rect 13277 18241 13311 18275
rect 13461 18241 13495 18275
rect 15485 18241 15519 18275
rect 15577 18241 15611 18275
rect 17325 18241 17359 18275
rect 19809 18241 19843 18275
rect 20269 18241 20303 18275
rect 21373 18241 21407 18275
rect 21833 18241 21867 18275
rect 24225 18241 24259 18275
rect 11437 18173 11471 18207
rect 13185 18173 13219 18207
rect 16589 18173 16623 18207
rect 19717 18173 19751 18207
rect 21189 18173 21223 18207
rect 22477 18173 22511 18207
rect 23029 18173 23063 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 15393 18105 15427 18139
rect 16865 18105 16899 18139
rect 18705 18105 18739 18139
rect 21281 18105 21315 18139
rect 24041 18105 24075 18139
rect 12265 18037 12299 18071
rect 15025 18037 15059 18071
rect 16221 18037 16255 18071
rect 17877 18037 17911 18071
rect 18245 18037 18279 18071
rect 19625 18037 19659 18071
rect 23397 18037 23431 18071
rect 24133 18037 24167 18071
rect 25053 18037 25087 18071
rect 25421 18037 25455 18071
rect 13001 17833 13035 17867
rect 13461 17833 13495 17867
rect 14105 17833 14139 17867
rect 15025 17833 15059 17867
rect 16221 17833 16255 17867
rect 17969 17833 18003 17867
rect 18889 17833 18923 17867
rect 19625 17833 19659 17867
rect 20913 17833 20947 17867
rect 22109 17833 22143 17867
rect 24317 17833 24351 17867
rect 24685 17833 24719 17867
rect 14565 17765 14599 17799
rect 16856 17765 16890 17799
rect 19717 17765 19751 17799
rect 23204 17765 23238 17799
rect 11713 17697 11747 17731
rect 13369 17697 13403 17731
rect 15301 17697 15335 17731
rect 19165 17697 19199 17731
rect 20729 17697 20763 17731
rect 21281 17697 21315 17731
rect 25145 17697 25179 17731
rect 11989 17629 12023 17663
rect 12909 17629 12943 17663
rect 13645 17629 13679 17663
rect 15577 17629 15611 17663
rect 16589 17629 16623 17663
rect 19901 17629 19935 17663
rect 21373 17629 21407 17663
rect 21465 17629 21499 17663
rect 22937 17629 22971 17663
rect 12541 17561 12575 17595
rect 19257 17561 19291 17595
rect 20269 17561 20303 17595
rect 11621 17493 11655 17527
rect 18245 17493 18279 17527
rect 18981 17493 19015 17527
rect 22477 17493 22511 17527
rect 25329 17493 25363 17527
rect 10977 17289 11011 17323
rect 14197 17289 14231 17323
rect 19349 17289 19383 17323
rect 22385 17289 22419 17323
rect 23121 17289 23155 17323
rect 14657 17221 14691 17255
rect 22017 17221 22051 17255
rect 25329 17221 25363 17255
rect 11345 17153 11379 17187
rect 18613 17153 18647 17187
rect 19993 17153 20027 17187
rect 21557 17153 21591 17187
rect 22569 17153 22603 17187
rect 11069 17085 11103 17119
rect 12449 17085 12483 17119
rect 14841 17085 14875 17119
rect 15577 17085 15611 17119
rect 17877 17085 17911 17119
rect 19717 17085 19751 17119
rect 20637 17085 20671 17119
rect 21373 17085 21407 17119
rect 23673 17085 23707 17119
rect 11897 17017 11931 17051
rect 12716 17017 12750 17051
rect 14565 17017 14599 17051
rect 15485 17017 15519 17051
rect 15822 17017 15856 17051
rect 18429 17017 18463 17051
rect 20821 17017 20855 17051
rect 21465 17017 21499 17051
rect 23489 17017 23523 17051
rect 23940 17017 23974 17051
rect 12173 16949 12207 16983
rect 13829 16949 13863 16983
rect 16957 16949 16991 16983
rect 17417 16949 17451 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 20453 16949 20487 16983
rect 20637 16949 20671 16983
rect 21005 16949 21039 16983
rect 25053 16949 25087 16983
rect 10885 16745 10919 16779
rect 14473 16745 14507 16779
rect 14841 16745 14875 16779
rect 16681 16745 16715 16779
rect 16957 16745 16991 16779
rect 17877 16745 17911 16779
rect 18153 16745 18187 16779
rect 18521 16745 18555 16779
rect 19349 16745 19383 16779
rect 20269 16745 20303 16779
rect 20729 16745 20763 16779
rect 22293 16745 22327 16779
rect 23949 16745 23983 16779
rect 24317 16745 24351 16779
rect 11989 16677 12023 16711
rect 15568 16677 15602 16711
rect 17417 16677 17451 16711
rect 23857 16677 23891 16711
rect 24869 16677 24903 16711
rect 11253 16609 11287 16643
rect 11345 16609 11379 16643
rect 12716 16609 12750 16643
rect 15301 16609 15335 16643
rect 17693 16609 17727 16643
rect 18061 16609 18095 16643
rect 18613 16609 18647 16643
rect 19717 16609 19751 16643
rect 21281 16609 21315 16643
rect 22661 16609 22695 16643
rect 23397 16609 23431 16643
rect 11529 16541 11563 16575
rect 12449 16541 12483 16575
rect 18705 16541 18739 16575
rect 21373 16541 21407 16575
rect 21465 16541 21499 16575
rect 22937 16541 22971 16575
rect 24409 16541 24443 16575
rect 24501 16541 24535 16575
rect 12357 16405 12391 16439
rect 13829 16405 13863 16439
rect 14105 16405 14139 16439
rect 19901 16405 19935 16439
rect 20913 16405 20947 16439
rect 22017 16405 22051 16439
rect 24869 16405 24903 16439
rect 25053 16405 25087 16439
rect 11253 16201 11287 16235
rect 11713 16201 11747 16235
rect 12449 16201 12483 16235
rect 13553 16201 13587 16235
rect 15393 16201 15427 16235
rect 15761 16201 15795 16235
rect 19441 16201 19475 16235
rect 23029 16201 23063 16235
rect 23489 16201 23523 16235
rect 24041 16201 24075 16235
rect 25053 16201 25087 16235
rect 14013 16133 14047 16167
rect 16773 16133 16807 16167
rect 22661 16133 22695 16167
rect 25421 16133 25455 16167
rect 12909 16065 12943 16099
rect 13093 16065 13127 16099
rect 14473 16065 14507 16099
rect 14565 16065 14599 16099
rect 16221 16065 16255 16099
rect 16405 16065 16439 16099
rect 23857 16065 23891 16099
rect 24593 16065 24627 16099
rect 25605 16065 25639 16099
rect 18061 15997 18095 16031
rect 20269 15997 20303 16031
rect 22293 15997 22327 16031
rect 22477 15997 22511 16031
rect 24501 15997 24535 16031
rect 12265 15929 12299 15963
rect 18328 15929 18362 15963
rect 20536 15929 20570 15963
rect 21925 15929 21959 15963
rect 10977 15861 11011 15895
rect 12817 15861 12851 15895
rect 13829 15861 13863 15895
rect 14381 15861 14415 15895
rect 16129 15861 16163 15895
rect 17509 15861 17543 15895
rect 17877 15861 17911 15895
rect 19809 15861 19843 15895
rect 20177 15861 20211 15895
rect 21649 15861 21683 15895
rect 24409 15861 24443 15895
rect 13277 15657 13311 15691
rect 14013 15657 14047 15691
rect 14657 15657 14691 15691
rect 15025 15657 15059 15691
rect 16589 15657 16623 15691
rect 18153 15657 18187 15691
rect 19257 15657 19291 15691
rect 20361 15657 20395 15691
rect 24409 15657 24443 15691
rect 25605 15657 25639 15691
rect 15669 15589 15703 15623
rect 16221 15589 16255 15623
rect 17141 15589 17175 15623
rect 21373 15589 21407 15623
rect 12164 15521 12198 15555
rect 15393 15521 15427 15555
rect 17049 15521 17083 15555
rect 18245 15521 18279 15555
rect 19625 15521 19659 15555
rect 19717 15521 19751 15555
rect 21097 15521 21131 15555
rect 22652 15521 22686 15555
rect 24961 15521 24995 15555
rect 11897 15453 11931 15487
rect 14105 15453 14139 15487
rect 17233 15453 17267 15487
rect 19165 15453 19199 15487
rect 19809 15453 19843 15487
rect 21833 15453 21867 15487
rect 22293 15453 22327 15487
rect 22385 15453 22419 15487
rect 25053 15453 25087 15487
rect 25145 15453 25179 15487
rect 18705 15385 18739 15419
rect 24593 15385 24627 15419
rect 10885 15317 10919 15351
rect 11345 15317 11379 15351
rect 11713 15317 11747 15351
rect 13553 15317 13587 15351
rect 16681 15317 16715 15351
rect 17693 15317 17727 15351
rect 20729 15317 20763 15351
rect 23765 15317 23799 15351
rect 24133 15317 24167 15351
rect 12633 15113 12667 15147
rect 15853 15113 15887 15147
rect 16313 15113 16347 15147
rect 21557 15113 21591 15147
rect 22201 15113 22235 15147
rect 25513 15113 25547 15147
rect 26249 15113 26283 15147
rect 15577 15045 15611 15079
rect 16405 15045 16439 15079
rect 21281 15045 21315 15079
rect 23029 15045 23063 15079
rect 23949 15045 23983 15079
rect 10701 14977 10735 15011
rect 11437 14977 11471 15011
rect 11897 14977 11931 15011
rect 13185 14977 13219 15011
rect 13645 14977 13679 15011
rect 14197 14977 14231 15011
rect 16957 14977 16991 15011
rect 18613 14977 18647 15011
rect 22477 14977 22511 15011
rect 11253 14909 11287 14943
rect 13001 14909 13035 14943
rect 16773 14909 16807 14943
rect 16865 14909 16899 14943
rect 19901 14909 19935 14943
rect 22293 14909 22327 14943
rect 24133 14909 24167 14943
rect 10333 14841 10367 14875
rect 11161 14841 11195 14875
rect 14105 14841 14139 14875
rect 14442 14841 14476 14875
rect 18429 14841 18463 14875
rect 19717 14841 19751 14875
rect 20168 14841 20202 14875
rect 23489 14841 23523 14875
rect 24400 14841 24434 14875
rect 25789 14841 25823 14875
rect 10793 14773 10827 14807
rect 12265 14773 12299 14807
rect 13093 14773 13127 14807
rect 17417 14773 17451 14807
rect 17785 14773 17819 14807
rect 18061 14773 18095 14807
rect 18521 14773 18555 14807
rect 19349 14773 19383 14807
rect 9965 14569 9999 14603
rect 12725 14569 12759 14603
rect 13645 14569 13679 14603
rect 15117 14569 15151 14603
rect 16405 14569 16439 14603
rect 16681 14569 16715 14603
rect 20913 14569 20947 14603
rect 21373 14569 21407 14603
rect 22477 14569 22511 14603
rect 22845 14569 22879 14603
rect 24041 14569 24075 14603
rect 11244 14501 11278 14535
rect 14013 14501 14047 14535
rect 15577 14501 15611 14535
rect 16129 14501 16163 14535
rect 10517 14433 10551 14467
rect 10977 14433 11011 14467
rect 14105 14433 14139 14467
rect 15301 14433 15335 14467
rect 22937 14501 22971 14535
rect 24501 14501 24535 14535
rect 17029 14433 17063 14467
rect 19625 14433 19659 14467
rect 19717 14433 19751 14467
rect 21281 14433 21315 14467
rect 24409 14433 24443 14467
rect 14197 14365 14231 14399
rect 16681 14365 16715 14399
rect 16773 14365 16807 14399
rect 19809 14365 19843 14399
rect 20729 14365 20763 14399
rect 21557 14365 21591 14399
rect 23121 14365 23155 14399
rect 24685 14365 24719 14399
rect 25145 14365 25179 14399
rect 19165 14297 19199 14331
rect 23949 14297 23983 14331
rect 10885 14229 10919 14263
rect 12357 14229 12391 14263
rect 13185 14229 13219 14263
rect 13461 14229 13495 14263
rect 14749 14229 14783 14263
rect 18153 14229 18187 14263
rect 18429 14229 18463 14263
rect 19257 14229 19291 14263
rect 20361 14229 20395 14263
rect 22109 14229 22143 14263
rect 23581 14229 23615 14263
rect 25421 14229 25455 14263
rect 11897 14025 11931 14059
rect 12265 14025 12299 14059
rect 13645 14025 13679 14059
rect 14657 14025 14691 14059
rect 15117 14025 15151 14059
rect 17877 14025 17911 14059
rect 20085 14025 20119 14059
rect 20269 14025 20303 14059
rect 21373 14025 21407 14059
rect 23397 14025 23431 14059
rect 24041 14025 24075 14059
rect 24593 14025 24627 14059
rect 25605 14025 25639 14059
rect 9413 13957 9447 13991
rect 10793 13957 10827 13991
rect 13553 13957 13587 13991
rect 16589 13957 16623 13991
rect 17417 13957 17451 13991
rect 19809 13957 19843 13991
rect 21833 13957 21867 13991
rect 9781 13889 9815 13923
rect 11345 13889 11379 13923
rect 14105 13889 14139 13923
rect 14197 13889 14231 13923
rect 20821 13889 20855 13923
rect 22569 13889 22603 13923
rect 25237 13889 25271 13923
rect 9505 13821 9539 13855
rect 10333 13821 10367 13855
rect 11253 13821 11287 13855
rect 13185 13821 13219 13855
rect 15209 13821 15243 13855
rect 15476 13821 15510 13855
rect 18061 13821 18095 13855
rect 23029 13821 23063 13855
rect 24409 13821 24443 13855
rect 25053 13821 25087 13855
rect 18306 13753 18340 13787
rect 20637 13753 20671 13787
rect 22385 13753 22419 13787
rect 22477 13753 22511 13787
rect 24961 13753 24995 13787
rect 10701 13685 10735 13719
rect 11161 13685 11195 13719
rect 12633 13685 12667 13719
rect 14013 13685 14047 13719
rect 17141 13685 17175 13719
rect 19441 13685 19475 13719
rect 20729 13685 20763 13719
rect 22017 13685 22051 13719
rect 10057 13481 10091 13515
rect 10149 13481 10183 13515
rect 12541 13481 12575 13515
rect 13185 13481 13219 13515
rect 15485 13481 15519 13515
rect 16589 13481 16623 13515
rect 16865 13481 16899 13515
rect 18337 13481 18371 13515
rect 20729 13481 20763 13515
rect 21649 13481 21683 13515
rect 23305 13481 23339 13515
rect 11428 13413 11462 13447
rect 15853 13413 15887 13447
rect 17049 13413 17083 13447
rect 19134 13413 19168 13447
rect 24102 13413 24136 13447
rect 14013 13345 14047 13379
rect 14105 13345 14139 13379
rect 18889 13345 18923 13379
rect 20913 13345 20947 13379
rect 22661 13345 22695 13379
rect 11161 13277 11195 13311
rect 13553 13277 13587 13311
rect 14289 13277 14323 13311
rect 15945 13277 15979 13311
rect 16037 13277 16071 13311
rect 21097 13277 21131 13311
rect 22753 13277 22787 13311
rect 22937 13277 22971 13311
rect 23857 13277 23891 13311
rect 13645 13209 13679 13243
rect 14749 13209 14783 13243
rect 10885 13141 10919 13175
rect 15025 13141 15059 13175
rect 20269 13141 20303 13175
rect 22109 13141 22143 13175
rect 22293 13141 22327 13175
rect 23673 13141 23707 13175
rect 25237 13141 25271 13175
rect 10793 12937 10827 12971
rect 11805 12937 11839 12971
rect 14105 12937 14139 12971
rect 16037 12937 16071 12971
rect 17049 12937 17083 12971
rect 19441 12937 19475 12971
rect 22937 12937 22971 12971
rect 23489 12937 23523 12971
rect 25053 12937 25087 12971
rect 12173 12869 12207 12903
rect 18337 12869 18371 12903
rect 19717 12869 19751 12903
rect 10333 12801 10367 12835
rect 11437 12801 11471 12835
rect 16773 12801 16807 12835
rect 17601 12801 17635 12835
rect 18797 12801 18831 12835
rect 18889 12801 18923 12835
rect 19901 12801 19935 12835
rect 22385 12801 22419 12835
rect 12449 12733 12483 12767
rect 12705 12733 12739 12767
rect 14657 12733 14691 12767
rect 17417 12733 17451 12767
rect 20157 12733 20191 12767
rect 21557 12733 21591 12767
rect 22109 12733 22143 12767
rect 23673 12733 23707 12767
rect 25329 12733 25363 12767
rect 25697 12733 25731 12767
rect 10701 12665 10735 12699
rect 11161 12665 11195 12699
rect 14565 12665 14599 12699
rect 14902 12665 14936 12699
rect 16681 12665 16715 12699
rect 17509 12665 17543 12699
rect 18705 12665 18739 12699
rect 21925 12665 21959 12699
rect 23918 12665 23952 12699
rect 11253 12597 11287 12631
rect 13829 12597 13863 12631
rect 21281 12597 21315 12631
rect 10517 12393 10551 12427
rect 11529 12393 11563 12427
rect 12081 12393 12115 12427
rect 13645 12393 13679 12427
rect 15301 12393 15335 12427
rect 16773 12393 16807 12427
rect 19257 12393 19291 12427
rect 20545 12393 20579 12427
rect 22569 12393 22603 12427
rect 22937 12393 22971 12427
rect 25605 12393 25639 12427
rect 10885 12325 10919 12359
rect 14749 12325 14783 12359
rect 18889 12325 18923 12359
rect 24492 12325 24526 12359
rect 12449 12257 12483 12291
rect 13185 12257 13219 12291
rect 14013 12257 14047 12291
rect 14105 12257 14139 12291
rect 15669 12257 15703 12291
rect 17233 12257 17267 12291
rect 18705 12257 18739 12291
rect 19625 12257 19659 12291
rect 21180 12257 21214 12291
rect 23121 12257 23155 12291
rect 10977 12189 11011 12223
rect 11161 12189 11195 12223
rect 12541 12189 12575 12223
rect 12725 12189 12759 12223
rect 14289 12189 14323 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 17325 12189 17359 12223
rect 17417 12189 17451 12223
rect 13553 12121 13587 12155
rect 16865 12121 16899 12155
rect 18153 12121 18187 12155
rect 19717 12189 19751 12223
rect 19901 12189 19935 12223
rect 20913 12189 20947 12223
rect 24041 12189 24075 12223
rect 24225 12189 24259 12223
rect 11989 12053 12023 12087
rect 15025 12053 15059 12087
rect 16313 12053 16347 12087
rect 18429 12053 18463 12087
rect 18705 12053 18739 12087
rect 22293 12053 22327 12087
rect 23765 12053 23799 12087
rect 10609 11849 10643 11883
rect 12173 11849 12207 11883
rect 12265 11849 12299 11883
rect 13369 11849 13403 11883
rect 16037 11849 16071 11883
rect 19533 11849 19567 11883
rect 20361 11849 20395 11883
rect 20453 11849 20487 11883
rect 21465 11849 21499 11883
rect 22017 11849 22051 11883
rect 10885 11781 10919 11815
rect 11805 11713 11839 11747
rect 15209 11781 15243 11815
rect 15577 11781 15611 11815
rect 12817 11713 12851 11747
rect 16589 11713 16623 11747
rect 17785 11713 17819 11747
rect 18613 11713 18647 11747
rect 21097 11713 21131 11747
rect 22661 11713 22695 11747
rect 24225 11713 24259 11747
rect 24777 11713 24811 11747
rect 24869 11713 24903 11747
rect 12541 11645 12575 11679
rect 13829 11645 13863 11679
rect 16405 11645 16439 11679
rect 18429 11645 18463 11679
rect 20821 11645 20855 11679
rect 21925 11645 21959 11679
rect 23489 11645 23523 11679
rect 11345 11577 11379 11611
rect 12265 11577 12299 11611
rect 14074 11577 14108 11611
rect 19073 11577 19107 11611
rect 20913 11577 20947 11611
rect 23029 11577 23063 11611
rect 25329 11577 25363 11611
rect 25697 11577 25731 11611
rect 13737 11509 13771 11543
rect 15945 11509 15979 11543
rect 16497 11509 16531 11543
rect 17049 11509 17083 11543
rect 17417 11509 17451 11543
rect 18061 11509 18095 11543
rect 18521 11509 18555 11543
rect 19901 11509 19935 11543
rect 22385 11509 22419 11543
rect 22477 11509 22511 11543
rect 24317 11509 24351 11543
rect 24685 11509 24719 11543
rect 12173 11305 12207 11339
rect 13461 11305 13495 11339
rect 14749 11305 14783 11339
rect 15301 11305 15335 11339
rect 18061 11305 18095 11339
rect 19165 11305 19199 11339
rect 19257 11305 19291 11339
rect 19625 11305 19659 11339
rect 20269 11305 20303 11339
rect 20729 11305 20763 11339
rect 21005 11305 21039 11339
rect 21373 11305 21407 11339
rect 22109 11305 22143 11339
rect 22477 11305 22511 11339
rect 24133 11305 24167 11339
rect 24869 11305 24903 11339
rect 25145 11305 25179 11339
rect 16313 11237 16347 11271
rect 16681 11237 16715 11271
rect 22998 11237 23032 11271
rect 13921 11169 13955 11203
rect 15669 11169 15703 11203
rect 17509 11169 17543 11203
rect 17969 11169 18003 11203
rect 19717 11169 19751 11203
rect 24961 11169 24995 11203
rect 14013 11101 14047 11135
rect 14197 11101 14231 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 18245 11101 18279 11135
rect 19901 11101 19935 11135
rect 21465 11101 21499 11135
rect 21557 11101 21591 11135
rect 22753 11101 22787 11135
rect 12633 11033 12667 11067
rect 13553 11033 13587 11067
rect 15025 11033 15059 11067
rect 17601 11033 17635 11067
rect 24501 11033 24535 11067
rect 13093 10965 13127 10999
rect 17141 10965 17175 10999
rect 18613 10965 18647 10999
rect 14657 10761 14691 10795
rect 15761 10761 15795 10795
rect 17601 10761 17635 10795
rect 19441 10761 19475 10795
rect 19809 10761 19843 10795
rect 20177 10761 20211 10795
rect 21097 10761 21131 10795
rect 23397 10761 23431 10795
rect 25789 10761 25823 10795
rect 22753 10693 22787 10727
rect 15209 10625 15243 10659
rect 16313 10625 16347 10659
rect 16957 10625 16991 10659
rect 20269 10625 20303 10659
rect 24317 10625 24351 10659
rect 25329 10625 25363 10659
rect 13001 10557 13035 10591
rect 13268 10557 13302 10591
rect 16773 10557 16807 10591
rect 18061 10557 18095 10591
rect 21373 10557 21407 10591
rect 21640 10557 21674 10591
rect 23029 10557 23063 10591
rect 24133 10557 24167 10591
rect 25145 10557 25179 10591
rect 12265 10489 12299 10523
rect 18328 10489 18362 10523
rect 12817 10421 12851 10455
rect 14381 10421 14415 10455
rect 15025 10421 15059 10455
rect 16405 10421 16439 10455
rect 16865 10421 16899 10455
rect 23765 10421 23799 10455
rect 24225 10421 24259 10455
rect 24777 10421 24811 10455
rect 26157 10421 26191 10455
rect 12633 10217 12667 10251
rect 14105 10217 14139 10251
rect 14473 10217 14507 10251
rect 15577 10217 15611 10251
rect 16681 10217 16715 10251
rect 17049 10217 17083 10251
rect 18797 10217 18831 10251
rect 19349 10217 19383 10251
rect 21373 10217 21407 10251
rect 22753 10217 22787 10251
rect 23581 10217 23615 10251
rect 25145 10217 25179 10251
rect 12970 10149 13004 10183
rect 17386 10149 17420 10183
rect 19257 10149 19291 10183
rect 20361 10149 20395 10183
rect 22293 10149 22327 10183
rect 24010 10149 24044 10183
rect 11529 10081 11563 10115
rect 11621 10081 11655 10115
rect 12725 10081 12759 10115
rect 15945 10081 15979 10115
rect 20729 10081 20763 10115
rect 21281 10081 21315 10115
rect 23213 10081 23247 10115
rect 23765 10081 23799 10115
rect 25421 10081 25455 10115
rect 11805 10013 11839 10047
rect 16037 10013 16071 10047
rect 16221 10013 16255 10047
rect 17141 10013 17175 10047
rect 21557 10013 21591 10047
rect 10885 9877 10919 9911
rect 11161 9877 11195 9911
rect 15025 9877 15059 9911
rect 18521 9877 18555 9911
rect 19901 9877 19935 9911
rect 20545 9877 20579 9911
rect 20913 9877 20947 9911
rect 21925 9877 21959 9911
rect 11897 9673 11931 9707
rect 12265 9673 12299 9707
rect 14289 9673 14323 9707
rect 15025 9673 15059 9707
rect 21649 9673 21683 9707
rect 23857 9673 23891 9707
rect 10793 9605 10827 9639
rect 13461 9605 13495 9639
rect 16497 9605 16531 9639
rect 17325 9605 17359 9639
rect 21281 9605 21315 9639
rect 9965 9537 9999 9571
rect 10333 9537 10367 9571
rect 11437 9537 11471 9571
rect 12909 9537 12943 9571
rect 13369 9537 13403 9571
rect 14013 9537 14047 9571
rect 14289 9537 14323 9571
rect 15945 9537 15979 9571
rect 16129 9537 16163 9571
rect 17877 9537 17911 9571
rect 18613 9537 18647 9571
rect 19625 9537 19659 9571
rect 22385 9537 22419 9571
rect 24501 9537 24535 9571
rect 24869 9537 24903 9571
rect 25237 9537 25271 9571
rect 13829 9469 13863 9503
rect 13921 9469 13955 9503
rect 15209 9469 15243 9503
rect 16865 9469 16899 9503
rect 18429 9469 18463 9503
rect 19073 9469 19107 9503
rect 22201 9469 22235 9503
rect 22293 9469 22327 9503
rect 10701 9401 10735 9435
rect 15853 9401 15887 9435
rect 18521 9401 18555 9435
rect 19533 9401 19567 9435
rect 19870 9401 19904 9435
rect 24317 9401 24351 9435
rect 11161 9333 11195 9367
rect 11253 9333 11287 9367
rect 12449 9333 12483 9367
rect 14473 9333 14507 9367
rect 14841 9333 14875 9367
rect 15485 9333 15519 9367
rect 18061 9333 18095 9367
rect 21005 9333 21039 9367
rect 21833 9333 21867 9367
rect 23029 9333 23063 9367
rect 23489 9333 23523 9367
rect 24225 9333 24259 9367
rect 25421 9333 25455 9367
rect 13185 9129 13219 9163
rect 13829 9129 13863 9163
rect 15117 9129 15151 9163
rect 17233 9129 17267 9163
rect 17969 9129 18003 9163
rect 18337 9129 18371 9163
rect 20729 9129 20763 9163
rect 23029 9129 23063 9163
rect 23489 9129 23523 9163
rect 23581 9129 23615 9163
rect 25145 9129 25179 9163
rect 10793 9061 10827 9095
rect 11713 9061 11747 9095
rect 13553 9061 13587 9095
rect 14749 9061 14783 9095
rect 18797 9061 18831 9095
rect 19625 9061 19659 9095
rect 10517 8993 10551 9027
rect 11805 8993 11839 9027
rect 12072 8993 12106 9027
rect 15669 8993 15703 9027
rect 15761 8993 15795 9027
rect 19717 8993 19751 9027
rect 20913 8993 20947 9027
rect 21180 8993 21214 9027
rect 24021 8993 24055 9027
rect 14197 8925 14231 8959
rect 15945 8925 15979 8959
rect 17325 8925 17359 8959
rect 17509 8925 17543 8959
rect 19165 8925 19199 8959
rect 19901 8925 19935 8959
rect 23489 8925 23523 8959
rect 23765 8925 23799 8959
rect 16865 8857 16899 8891
rect 11253 8789 11287 8823
rect 15301 8789 15335 8823
rect 16405 8789 16439 8823
rect 16681 8789 16715 8823
rect 19257 8789 19291 8823
rect 20269 8789 20303 8823
rect 22293 8789 22327 8823
rect 22661 8789 22695 8823
rect 11529 8585 11563 8619
rect 11897 8585 11931 8619
rect 12173 8585 12207 8619
rect 13829 8585 13863 8619
rect 17417 8585 17451 8619
rect 17877 8585 17911 8619
rect 19441 8585 19475 8619
rect 19809 8585 19843 8619
rect 20361 8585 20395 8619
rect 24225 8585 24259 8619
rect 12449 8517 12483 8551
rect 14289 8517 14323 8551
rect 22109 8517 22143 8551
rect 22385 8517 22419 8551
rect 24317 8517 24351 8551
rect 13001 8449 13035 8483
rect 24777 8449 24811 8483
rect 24961 8449 24995 8483
rect 25329 8449 25363 8483
rect 10149 8381 10183 8415
rect 14473 8381 14507 8415
rect 14565 8381 14599 8415
rect 14832 8381 14866 8415
rect 16497 8381 16531 8415
rect 18061 8381 18095 8415
rect 18317 8381 18351 8415
rect 20545 8381 20579 8415
rect 20729 8381 20763 8415
rect 23489 8381 23523 8415
rect 24685 8381 24719 8415
rect 10057 8313 10091 8347
rect 10394 8313 10428 8347
rect 14197 8313 14231 8347
rect 16773 8313 16807 8347
rect 16957 8313 16991 8347
rect 20974 8313 21008 8347
rect 23121 8313 23155 8347
rect 12817 8245 12851 8279
rect 12909 8245 12943 8279
rect 15945 8245 15979 8279
rect 20269 8245 20303 8279
rect 10609 8041 10643 8075
rect 12173 8041 12207 8075
rect 12817 8041 12851 8075
rect 13001 8041 13035 8075
rect 14289 8041 14323 8075
rect 15669 8041 15703 8075
rect 16865 8041 16899 8075
rect 19257 8041 19291 8075
rect 21373 8041 21407 8075
rect 21925 8041 21959 8075
rect 22293 8041 22327 8075
rect 25053 8041 25087 8075
rect 12541 7973 12575 8007
rect 16681 7973 16715 8007
rect 18061 7973 18095 8007
rect 19717 7973 19751 8007
rect 20637 7973 20671 8007
rect 11060 7905 11094 7939
rect 13369 7905 13403 7939
rect 17233 7905 17267 7939
rect 18889 7905 18923 7939
rect 19625 7905 19659 7939
rect 21281 7905 21315 7939
rect 23940 7905 23974 7939
rect 10241 7837 10275 7871
rect 10793 7837 10827 7871
rect 13461 7837 13495 7871
rect 13553 7837 13587 7871
rect 15761 7837 15795 7871
rect 15853 7837 15887 7871
rect 17325 7837 17359 7871
rect 17509 7837 17543 7871
rect 19901 7837 19935 7871
rect 21557 7837 21591 7871
rect 22569 7837 22603 7871
rect 23673 7837 23707 7871
rect 15301 7769 15335 7803
rect 20913 7769 20947 7803
rect 14657 7701 14691 7735
rect 15025 7701 15059 7735
rect 16313 7701 16347 7735
rect 18521 7701 18555 7735
rect 23489 7701 23523 7735
rect 12725 7497 12759 7531
rect 13093 7497 13127 7531
rect 15577 7497 15611 7531
rect 17601 7497 17635 7531
rect 18705 7497 18739 7531
rect 19809 7497 19843 7531
rect 20545 7497 20579 7531
rect 21557 7497 21591 7531
rect 21925 7497 21959 7531
rect 25053 7497 25087 7531
rect 10793 7429 10827 7463
rect 12173 7429 12207 7463
rect 11437 7361 11471 7395
rect 16313 7361 16347 7395
rect 16957 7361 16991 7395
rect 18337 7361 18371 7395
rect 19349 7361 19383 7395
rect 21005 7361 21039 7395
rect 21189 7361 21223 7395
rect 9781 7293 9815 7327
rect 13369 7293 13403 7327
rect 16129 7293 16163 7327
rect 16221 7293 16255 7327
rect 19165 7293 19199 7327
rect 22385 7293 22419 7327
rect 23673 7293 23707 7327
rect 25329 7293 25363 7327
rect 10333 7225 10367 7259
rect 11253 7225 11287 7259
rect 13614 7225 13648 7259
rect 15301 7225 15335 7259
rect 19257 7225 19291 7259
rect 20913 7225 20947 7259
rect 23489 7225 23523 7259
rect 23940 7225 23974 7259
rect 10609 7157 10643 7191
rect 11161 7157 11195 7191
rect 11897 7157 11931 7191
rect 14749 7157 14783 7191
rect 15761 7157 15795 7191
rect 17233 7157 17267 7191
rect 18797 7157 18831 7191
rect 20269 7157 20303 7191
rect 22569 7157 22603 7191
rect 23029 7157 23063 7191
rect 11161 6953 11195 6987
rect 11529 6953 11563 6987
rect 12081 6953 12115 6987
rect 13461 6953 13495 6987
rect 14013 6953 14047 6987
rect 14749 6953 14783 6987
rect 18153 6953 18187 6987
rect 19625 6953 19659 6987
rect 20637 6953 20671 6987
rect 21189 6953 21223 6987
rect 22661 6953 22695 6987
rect 23765 6953 23799 6987
rect 12449 6885 12483 6919
rect 15853 6885 15887 6919
rect 16497 6885 16531 6919
rect 18061 6885 18095 6919
rect 9781 6817 9815 6851
rect 10037 6817 10071 6851
rect 11989 6817 12023 6851
rect 15025 6817 15059 6851
rect 17233 6817 17267 6851
rect 17509 6817 17543 6851
rect 19717 6817 19751 6851
rect 21537 6817 21571 6851
rect 24225 6817 24259 6851
rect 12541 6749 12575 6783
rect 12725 6749 12759 6783
rect 14105 6749 14139 6783
rect 14289 6749 14323 6783
rect 15945 6749 15979 6783
rect 16129 6749 16163 6783
rect 18245 6749 18279 6783
rect 19901 6749 19935 6783
rect 21281 6749 21315 6783
rect 24317 6749 24351 6783
rect 24409 6749 24443 6783
rect 25421 6749 25455 6783
rect 13645 6681 13679 6715
rect 16865 6681 16899 6715
rect 17693 6681 17727 6715
rect 15485 6613 15519 6647
rect 17049 6613 17083 6647
rect 18797 6613 18831 6647
rect 19257 6613 19291 6647
rect 22937 6613 22971 6647
rect 23305 6613 23339 6647
rect 23857 6613 23891 6647
rect 9873 6409 9907 6443
rect 10241 6409 10275 6443
rect 10793 6409 10827 6443
rect 12173 6409 12207 6443
rect 12909 6409 12943 6443
rect 15117 6409 15151 6443
rect 17785 6409 17819 6443
rect 18337 6409 18371 6443
rect 20361 6409 20395 6443
rect 23121 6409 23155 6443
rect 23489 6409 23523 6443
rect 24501 6409 24535 6443
rect 25513 6409 25547 6443
rect 11437 6341 11471 6375
rect 13277 6341 13311 6375
rect 21005 6341 21039 6375
rect 22753 6341 22787 6375
rect 11805 6273 11839 6307
rect 13645 6273 13679 6307
rect 16405 6273 16439 6307
rect 16589 6273 16623 6307
rect 16957 6273 16991 6307
rect 18705 6273 18739 6307
rect 21373 6273 21407 6307
rect 25145 6273 25179 6307
rect 13737 6205 13771 6239
rect 14004 6205 14038 6239
rect 15485 6205 15519 6239
rect 21189 6205 21223 6239
rect 16313 6137 16347 6171
rect 17417 6137 17451 6171
rect 18950 6137 18984 6171
rect 20913 6137 20947 6171
rect 21640 6137 21674 6171
rect 23949 6137 23983 6171
rect 24869 6137 24903 6171
rect 15761 6069 15795 6103
rect 15945 6069 15979 6103
rect 20085 6069 20119 6103
rect 24409 6069 24443 6103
rect 24961 6069 24995 6103
rect 12081 5865 12115 5899
rect 13829 5865 13863 5899
rect 15117 5865 15151 5899
rect 17141 5865 17175 5899
rect 18889 5865 18923 5899
rect 19349 5865 19383 5899
rect 20729 5865 20763 5899
rect 21281 5865 21315 5899
rect 22293 5865 22327 5899
rect 23581 5865 23615 5899
rect 15568 5797 15602 5831
rect 24041 5797 24075 5831
rect 13001 5729 13035 5763
rect 14105 5729 14139 5763
rect 14657 5729 14691 5763
rect 17765 5729 17799 5763
rect 19717 5729 19751 5763
rect 22477 5729 22511 5763
rect 23949 5729 23983 5763
rect 25145 5729 25179 5763
rect 13093 5661 13127 5695
rect 15301 5661 15335 5695
rect 17509 5661 17543 5695
rect 21373 5661 21407 5695
rect 21557 5661 21591 5695
rect 21925 5661 21959 5695
rect 24225 5661 24259 5695
rect 22661 5593 22695 5627
rect 24685 5593 24719 5627
rect 14289 5525 14323 5559
rect 16681 5525 16715 5559
rect 19901 5525 19935 5559
rect 20269 5525 20303 5559
rect 20913 5525 20947 5559
rect 23029 5525 23063 5559
rect 23397 5525 23431 5559
rect 24961 5525 24995 5559
rect 25329 5525 25363 5559
rect 13737 5321 13771 5355
rect 14197 5321 14231 5355
rect 15393 5321 15427 5355
rect 19717 5321 19751 5355
rect 21373 5321 21407 5355
rect 21649 5321 21683 5355
rect 22293 5321 22327 5355
rect 23029 5321 23063 5355
rect 23397 5321 23431 5355
rect 25329 5321 25363 5355
rect 25053 5253 25087 5287
rect 14657 5185 14691 5219
rect 14841 5185 14875 5219
rect 18981 5185 19015 5219
rect 19993 5185 20027 5219
rect 23673 5185 23707 5219
rect 13093 5117 13127 5151
rect 14105 5117 14139 5151
rect 14565 5117 14599 5151
rect 15761 5117 15795 5151
rect 18337 5117 18371 5151
rect 18797 5117 18831 5151
rect 22477 5117 22511 5151
rect 16028 5049 16062 5083
rect 20238 5049 20272 5083
rect 23918 5049 23952 5083
rect 12909 4981 12943 5015
rect 13277 4981 13311 5015
rect 17141 4981 17175 5015
rect 17509 4981 17543 5015
rect 18429 4981 18463 5015
rect 18889 4981 18923 5015
rect 22661 4981 22695 5015
rect 25697 4981 25731 5015
rect 13001 4777 13035 4811
rect 14749 4777 14783 4811
rect 15117 4777 15151 4811
rect 15945 4777 15979 4811
rect 16037 4777 16071 4811
rect 16681 4777 16715 4811
rect 17325 4777 17359 4811
rect 17693 4777 17727 4811
rect 18889 4777 18923 4811
rect 21649 4777 21683 4811
rect 22109 4777 22143 4811
rect 24685 4777 24719 4811
rect 25053 4777 25087 4811
rect 14197 4709 14231 4743
rect 17785 4709 17819 4743
rect 19257 4709 19291 4743
rect 20361 4709 20395 4743
rect 12817 4641 12851 4675
rect 13921 4641 13955 4675
rect 20913 4641 20947 4675
rect 22744 4641 22778 4675
rect 25145 4641 25179 4675
rect 11805 4573 11839 4607
rect 13461 4573 13495 4607
rect 13829 4573 13863 4607
rect 16129 4573 16163 4607
rect 17877 4573 17911 4607
rect 19349 4573 19383 4607
rect 19441 4573 19475 4607
rect 19993 4573 20027 4607
rect 21097 4573 21131 4607
rect 22477 4573 22511 4607
rect 25237 4573 25271 4607
rect 24501 4505 24535 4539
rect 15577 4437 15611 4471
rect 17141 4437 17175 4471
rect 18429 4437 18463 4471
rect 23857 4437 23891 4471
rect 24133 4437 24167 4471
rect 14381 4233 14415 4267
rect 15669 4233 15703 4267
rect 17417 4233 17451 4267
rect 17785 4233 17819 4267
rect 18521 4233 18555 4267
rect 19441 4233 19475 4267
rect 20913 4233 20947 4267
rect 23489 4233 23523 4267
rect 25053 4233 25087 4267
rect 17049 4165 17083 4199
rect 19901 4165 19935 4199
rect 12265 4097 12299 4131
rect 13737 4097 13771 4131
rect 13921 4097 13955 4131
rect 14841 4097 14875 4131
rect 15209 4097 15243 4131
rect 16221 4097 16255 4131
rect 19717 4097 19751 4131
rect 20453 4097 20487 4131
rect 21557 4097 21591 4131
rect 22569 4097 22603 4131
rect 24133 4097 24167 4131
rect 24225 4097 24259 4131
rect 24777 4097 24811 4131
rect 11253 4029 11287 4063
rect 12817 4029 12851 4063
rect 15577 4029 15611 4063
rect 16129 4029 16163 4063
rect 18613 4029 18647 4063
rect 25237 4029 25271 4063
rect 25789 4029 25823 4063
rect 13645 3961 13679 3995
rect 16037 3961 16071 3995
rect 18889 3961 18923 3995
rect 20269 3961 20303 3995
rect 21833 3961 21867 3995
rect 22385 3961 22419 3995
rect 22477 3961 22511 3995
rect 24041 3961 24075 3995
rect 11437 3893 11471 3927
rect 11897 3893 11931 3927
rect 13093 3893 13127 3927
rect 13277 3893 13311 3927
rect 20361 3893 20395 3927
rect 22017 3893 22051 3927
rect 23029 3893 23063 3927
rect 23673 3893 23707 3927
rect 25421 3893 25455 3927
rect 14105 3689 14139 3723
rect 14657 3689 14691 3723
rect 16405 3689 16439 3723
rect 18337 3689 18371 3723
rect 18613 3689 18647 3723
rect 19257 3689 19291 3723
rect 21097 3689 21131 3723
rect 23765 3689 23799 3723
rect 24961 3689 24995 3723
rect 25329 3689 25363 3723
rect 12633 3621 12667 3655
rect 14013 3621 14047 3655
rect 15577 3621 15611 3655
rect 16129 3621 16163 3655
rect 24317 3621 24351 3655
rect 11253 3553 11287 3587
rect 12357 3553 12391 3587
rect 13369 3553 13403 3587
rect 15117 3553 15151 3587
rect 15301 3553 15335 3587
rect 16589 3553 16623 3587
rect 16856 3553 16890 3587
rect 19625 3553 19659 3587
rect 19717 3553 19751 3587
rect 22008 3553 22042 3587
rect 10241 3485 10275 3519
rect 14197 3485 14231 3519
rect 19809 3485 19843 3519
rect 21741 3485 21775 3519
rect 24409 3485 24443 3519
rect 24593 3485 24627 3519
rect 11437 3417 11471 3451
rect 13645 3417 13679 3451
rect 12265 3349 12299 3383
rect 17969 3349 18003 3383
rect 19165 3349 19199 3383
rect 20269 3349 20303 3383
rect 20637 3349 20671 3383
rect 21557 3349 21591 3383
rect 23121 3349 23155 3383
rect 23949 3349 23983 3383
rect 10701 3145 10735 3179
rect 12265 3145 12299 3179
rect 12817 3145 12851 3179
rect 14657 3145 14691 3179
rect 15301 3145 15335 3179
rect 16865 3145 16899 3179
rect 17141 3145 17175 3179
rect 17877 3145 17911 3179
rect 19533 3145 19567 3179
rect 19809 3145 19843 3179
rect 21925 3145 21959 3179
rect 22201 3145 22235 3179
rect 22569 3145 22603 3179
rect 23121 3145 23155 3179
rect 23489 3145 23523 3179
rect 24409 3145 24443 3179
rect 24777 3145 24811 3179
rect 10333 3077 10367 3111
rect 13185 3077 13219 3111
rect 14933 3077 14967 3111
rect 25145 3077 25179 3111
rect 11897 3009 11931 3043
rect 18153 3009 18187 3043
rect 20269 3009 20303 3043
rect 10149 2941 10183 2975
rect 11161 2941 11195 2975
rect 11253 2941 11287 2975
rect 13277 2941 13311 2975
rect 13544 2941 13578 2975
rect 15485 2941 15519 2975
rect 15741 2941 15775 2975
rect 20545 2941 20579 2975
rect 23673 2941 23707 2975
rect 24961 2941 24995 2975
rect 25513 2941 25547 2975
rect 18398 2873 18432 2907
rect 20790 2873 20824 2907
rect 23949 2873 23983 2907
rect 11437 2805 11471 2839
rect 10977 2601 11011 2635
rect 12449 2601 12483 2635
rect 13093 2601 13127 2635
rect 13369 2601 13403 2635
rect 14289 2601 14323 2635
rect 14933 2601 14967 2635
rect 16589 2601 16623 2635
rect 17049 2601 17083 2635
rect 17785 2601 17819 2635
rect 20269 2601 20303 2635
rect 20545 2601 20579 2635
rect 21465 2601 21499 2635
rect 22845 2601 22879 2635
rect 23213 2601 23247 2635
rect 23581 2601 23615 2635
rect 21925 2533 21959 2567
rect 24317 2533 24351 2567
rect 8585 2465 8619 2499
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 12725 2465 12759 2499
rect 13093 2465 13127 2499
rect 14197 2465 14231 2499
rect 15577 2465 15611 2499
rect 16129 2465 16163 2499
rect 18889 2465 18923 2499
rect 19156 2465 19190 2499
rect 20913 2465 20947 2499
rect 21833 2465 21867 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25329 2465 25363 2499
rect 25881 2465 25915 2499
rect 14473 2397 14507 2431
rect 15301 2397 15335 2431
rect 17141 2397 17175 2431
rect 17325 2397 17359 2431
rect 18797 2397 18831 2431
rect 22017 2397 22051 2431
rect 22477 2397 22511 2431
rect 12909 2329 12943 2363
rect 13829 2329 13863 2363
rect 18061 2329 18095 2363
rect 25513 2329 25547 2363
rect 8769 2261 8803 2295
rect 9229 2261 9263 2295
rect 10517 2261 10551 2295
rect 11621 2261 11655 2295
rect 13645 2261 13679 2295
rect 15761 2261 15795 2295
rect 16681 2261 16715 2295
<< metal1 >>
rect 16942 26800 16948 26852
rect 17000 26840 17006 26852
rect 23750 26840 23756 26852
rect 17000 26812 23756 26840
rect 17000 26800 17006 26812
rect 23750 26800 23756 26812
rect 23808 26800 23814 26852
rect 21542 26596 21548 26648
rect 21600 26636 21606 26648
rect 24762 26636 24768 26648
rect 21600 26608 24768 26636
rect 21600 26596 21606 26608
rect 24762 26596 24768 26608
rect 24820 26596 24826 26648
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 16669 25483 16727 25489
rect 16669 25449 16681 25483
rect 16715 25480 16727 25483
rect 17310 25480 17316 25492
rect 16715 25452 17316 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 17310 25440 17316 25452
rect 17368 25440 17374 25492
rect 19061 25483 19119 25489
rect 19061 25449 19073 25483
rect 19107 25449 19119 25483
rect 19061 25443 19119 25449
rect 22097 25483 22155 25489
rect 22097 25449 22109 25483
rect 22143 25480 22155 25483
rect 22738 25480 22744 25492
rect 22143 25452 22744 25480
rect 22143 25449 22155 25452
rect 22097 25443 22155 25449
rect 19076 25412 19104 25443
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 24670 25412 24676 25424
rect 19076 25384 24676 25412
rect 24670 25372 24676 25384
rect 24728 25372 24734 25424
rect 13998 25304 14004 25356
rect 14056 25344 14062 25356
rect 14277 25347 14335 25353
rect 14277 25344 14289 25347
rect 14056 25316 14289 25344
rect 14056 25304 14062 25316
rect 14277 25313 14289 25316
rect 14323 25313 14335 25347
rect 16482 25344 16488 25356
rect 16443 25316 16488 25344
rect 14277 25307 14335 25313
rect 16482 25304 16488 25316
rect 16540 25304 16546 25356
rect 18877 25347 18935 25353
rect 18877 25313 18889 25347
rect 18923 25344 18935 25347
rect 19242 25344 19248 25356
rect 18923 25316 19248 25344
rect 18923 25313 18935 25316
rect 18877 25307 18935 25313
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 19978 25344 19984 25356
rect 19939 25316 19984 25344
rect 19978 25304 19984 25316
rect 20036 25304 20042 25356
rect 21913 25347 21971 25353
rect 21913 25313 21925 25347
rect 21959 25344 21971 25347
rect 22554 25344 22560 25356
rect 21959 25316 22560 25344
rect 21959 25313 21971 25316
rect 21913 25307 21971 25313
rect 22554 25304 22560 25316
rect 22612 25304 22618 25356
rect 24210 25304 24216 25356
rect 24268 25344 24274 25356
rect 24581 25347 24639 25353
rect 24581 25344 24593 25347
rect 24268 25316 24593 25344
rect 24268 25304 24274 25316
rect 24581 25313 24593 25316
rect 24627 25313 24639 25347
rect 24581 25307 24639 25313
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25276 15531 25279
rect 18138 25276 18144 25288
rect 15519 25248 18144 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 18138 25236 18144 25248
rect 18196 25236 18202 25288
rect 26142 25276 26148 25288
rect 19076 25248 26148 25276
rect 14461 25211 14519 25217
rect 14461 25177 14473 25211
rect 14507 25208 14519 25211
rect 19076 25208 19104 25248
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 14507 25180 19104 25208
rect 20165 25211 20223 25217
rect 14507 25177 14519 25180
rect 14461 25171 14519 25177
rect 20165 25177 20177 25211
rect 20211 25208 20223 25211
rect 23474 25208 23480 25220
rect 20211 25180 23480 25208
rect 20211 25177 20223 25180
rect 20165 25171 20223 25177
rect 23474 25168 23480 25180
rect 23532 25168 23538 25220
rect 24762 25140 24768 25152
rect 24723 25112 24768 25140
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 20625 24939 20683 24945
rect 20625 24905 20637 24939
rect 20671 24936 20683 24939
rect 21358 24936 21364 24948
rect 20671 24908 21364 24936
rect 20671 24905 20683 24908
rect 20625 24899 20683 24905
rect 21358 24896 21364 24908
rect 21416 24896 21422 24948
rect 16022 24828 16028 24880
rect 16080 24868 16086 24880
rect 16482 24868 16488 24880
rect 16080 24840 16488 24868
rect 16080 24828 16086 24840
rect 16482 24828 16488 24840
rect 16540 24868 16546 24880
rect 16540 24840 16896 24868
rect 16540 24828 16546 24840
rect 16868 24809 16896 24840
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 13541 24735 13599 24741
rect 13541 24732 13553 24735
rect 13464 24704 13553 24732
rect 13464 24608 13492 24704
rect 13541 24701 13553 24704
rect 13587 24701 13599 24735
rect 13541 24695 13599 24701
rect 14550 24692 14556 24744
rect 14608 24732 14614 24744
rect 14645 24735 14703 24741
rect 14645 24732 14657 24735
rect 14608 24704 14657 24732
rect 14608 24692 14614 24704
rect 14645 24701 14657 24704
rect 14691 24732 14703 24735
rect 15381 24735 15439 24741
rect 15381 24732 15393 24735
rect 14691 24704 15393 24732
rect 14691 24701 14703 24704
rect 14645 24695 14703 24701
rect 15381 24701 15393 24704
rect 15427 24701 15439 24735
rect 15381 24695 15439 24701
rect 15933 24735 15991 24741
rect 15933 24701 15945 24735
rect 15979 24732 15991 24735
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 15979 24704 16620 24732
rect 15979 24701 15991 24704
rect 15933 24695 15991 24701
rect 14918 24664 14924 24676
rect 14879 24636 14924 24664
rect 14918 24624 14924 24636
rect 14976 24624 14982 24676
rect 13446 24596 13452 24608
rect 13407 24568 13452 24596
rect 13446 24556 13452 24568
rect 13504 24556 13510 24608
rect 13722 24596 13728 24608
rect 13683 24568 13728 24596
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 13998 24556 14004 24608
rect 14056 24596 14062 24608
rect 14277 24599 14335 24605
rect 14277 24596 14289 24599
rect 14056 24568 14289 24596
rect 14056 24556 14062 24568
rect 14277 24565 14289 24568
rect 14323 24565 14335 24599
rect 14277 24559 14335 24565
rect 16117 24599 16175 24605
rect 16117 24565 16129 24599
rect 16163 24596 16175 24599
rect 16390 24596 16396 24608
rect 16163 24568 16396 24596
rect 16163 24565 16175 24568
rect 16117 24559 16175 24565
rect 16390 24556 16396 24568
rect 16448 24556 16454 24608
rect 16592 24605 16620 24704
rect 17788 24704 18061 24732
rect 16577 24599 16635 24605
rect 16577 24565 16589 24599
rect 16623 24596 16635 24599
rect 17310 24596 17316 24608
rect 16623 24568 17316 24596
rect 16623 24565 16635 24568
rect 16577 24559 16635 24565
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 17402 24556 17408 24608
rect 17460 24596 17466 24608
rect 17788 24605 17816 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 19337 24735 19395 24741
rect 19337 24701 19349 24735
rect 19383 24732 19395 24735
rect 19426 24732 19432 24744
rect 19383 24704 19432 24732
rect 19383 24701 19395 24704
rect 19337 24695 19395 24701
rect 19426 24692 19432 24704
rect 19484 24692 19490 24744
rect 20162 24692 20168 24744
rect 20220 24732 20226 24744
rect 20441 24735 20499 24741
rect 20441 24732 20453 24735
rect 20220 24704 20453 24732
rect 20220 24692 20226 24704
rect 20441 24701 20453 24704
rect 20487 24732 20499 24735
rect 20993 24735 21051 24741
rect 20993 24732 21005 24735
rect 20487 24704 21005 24732
rect 20487 24701 20499 24704
rect 20441 24695 20499 24701
rect 20993 24701 21005 24704
rect 21039 24701 21051 24735
rect 20993 24695 21051 24701
rect 21545 24735 21603 24741
rect 21545 24701 21557 24735
rect 21591 24732 21603 24735
rect 22186 24732 22192 24744
rect 21591 24704 22192 24732
rect 21591 24701 21603 24704
rect 21545 24695 21603 24701
rect 22186 24692 22192 24704
rect 22244 24692 22250 24744
rect 24578 24732 24584 24744
rect 24539 24704 24584 24732
rect 24578 24692 24584 24704
rect 24636 24732 24642 24744
rect 25133 24735 25191 24741
rect 25133 24732 25145 24735
rect 24636 24704 25145 24732
rect 24636 24692 24642 24704
rect 25133 24701 25145 24704
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 20070 24664 20076 24676
rect 19536 24636 20076 24664
rect 17773 24599 17831 24605
rect 17773 24596 17785 24599
rect 17460 24568 17785 24596
rect 17460 24556 17466 24568
rect 17773 24565 17785 24568
rect 17819 24565 17831 24599
rect 17773 24559 17831 24565
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 18012 24568 18245 24596
rect 18012 24556 18018 24568
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 18233 24559 18291 24565
rect 18969 24599 19027 24605
rect 18969 24565 18981 24599
rect 19015 24596 19027 24599
rect 19242 24596 19248 24608
rect 19015 24568 19248 24596
rect 19015 24565 19027 24568
rect 18969 24559 19027 24565
rect 19242 24556 19248 24568
rect 19300 24556 19306 24608
rect 19536 24605 19564 24636
rect 20070 24624 20076 24636
rect 20128 24624 20134 24676
rect 19521 24599 19579 24605
rect 19521 24565 19533 24599
rect 19567 24565 19579 24599
rect 19978 24596 19984 24608
rect 19939 24568 19984 24596
rect 19521 24559 19579 24565
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 21729 24599 21787 24605
rect 21729 24565 21741 24599
rect 21775 24596 21787 24599
rect 22002 24596 22008 24608
rect 21775 24568 22008 24596
rect 21775 24565 21787 24568
rect 21729 24559 21787 24565
rect 22002 24556 22008 24568
rect 22060 24556 22066 24608
rect 22554 24596 22560 24608
rect 22467 24568 22560 24596
rect 22554 24556 22560 24568
rect 22612 24596 22618 24608
rect 23106 24596 23112 24608
rect 22612 24568 23112 24596
rect 22612 24556 22618 24568
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 24210 24556 24216 24608
rect 24268 24596 24274 24608
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 24268 24568 24409 24596
rect 24268 24556 24274 24568
rect 24397 24565 24409 24568
rect 24443 24565 24455 24599
rect 24762 24596 24768 24608
rect 24723 24568 24768 24596
rect 24397 24559 24455 24565
rect 24762 24556 24768 24568
rect 24820 24556 24826 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 12802 24392 12808 24404
rect 12763 24364 12808 24392
rect 12802 24352 12808 24364
rect 12860 24352 12866 24404
rect 14001 24395 14059 24401
rect 14001 24361 14013 24395
rect 14047 24392 14059 24395
rect 15102 24392 15108 24404
rect 14047 24364 15108 24392
rect 14047 24361 14059 24364
rect 14001 24355 14059 24361
rect 15102 24352 15108 24364
rect 15160 24352 15166 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 15930 24392 15936 24404
rect 15519 24364 15936 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 16206 24392 16212 24404
rect 16167 24364 16212 24392
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 18138 24392 18144 24404
rect 18099 24364 18144 24392
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 18690 24352 18696 24404
rect 18748 24392 18754 24404
rect 18877 24395 18935 24401
rect 18877 24392 18889 24395
rect 18748 24364 18889 24392
rect 18748 24352 18754 24364
rect 18877 24361 18889 24364
rect 18923 24361 18935 24395
rect 18877 24355 18935 24361
rect 20714 24352 20720 24404
rect 20772 24392 20778 24404
rect 21085 24395 21143 24401
rect 21085 24392 21097 24395
rect 20772 24364 21097 24392
rect 20772 24352 20778 24364
rect 21085 24361 21097 24364
rect 21131 24361 21143 24395
rect 21085 24355 21143 24361
rect 22557 24395 22615 24401
rect 22557 24361 22569 24395
rect 22603 24392 22615 24395
rect 23382 24392 23388 24404
rect 22603 24364 23388 24392
rect 22603 24361 22615 24364
rect 22557 24355 22615 24361
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 23658 24392 23664 24404
rect 23619 24364 23664 24392
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 16666 24284 16672 24336
rect 16724 24333 16730 24336
rect 16724 24327 16788 24333
rect 16724 24293 16742 24327
rect 16776 24293 16788 24327
rect 16724 24287 16788 24293
rect 16724 24284 16730 24287
rect 12158 24216 12164 24268
rect 12216 24256 12222 24268
rect 12618 24256 12624 24268
rect 12216 24228 12624 24256
rect 12216 24216 12222 24228
rect 12618 24216 12624 24228
rect 12676 24216 12682 24268
rect 13262 24216 13268 24268
rect 13320 24256 13326 24268
rect 13817 24259 13875 24265
rect 13817 24256 13829 24259
rect 13320 24228 13829 24256
rect 13320 24216 13326 24228
rect 13817 24225 13829 24228
rect 13863 24256 13875 24259
rect 14369 24259 14427 24265
rect 14369 24256 14381 24259
rect 13863 24228 14381 24256
rect 13863 24225 13875 24228
rect 13817 24219 13875 24225
rect 14369 24225 14381 24228
rect 14415 24225 14427 24259
rect 14369 24219 14427 24225
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 15746 24256 15752 24268
rect 15335 24228 15752 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15746 24216 15752 24228
rect 15804 24216 15810 24268
rect 18690 24256 18696 24268
rect 18651 24228 18696 24256
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 20898 24256 20904 24268
rect 20859 24228 20904 24256
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 22370 24256 22376 24268
rect 22331 24228 22376 24256
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 23474 24256 23480 24268
rect 23435 24228 23480 24256
rect 23474 24216 23480 24228
rect 23532 24216 23538 24268
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24176 24228 24593 24256
rect 24176 24216 24182 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 14826 24188 14832 24200
rect 14739 24160 14832 24188
rect 14826 24148 14832 24160
rect 14884 24188 14890 24200
rect 16485 24191 16543 24197
rect 16485 24188 16497 24191
rect 14884 24160 16497 24188
rect 14884 24148 14890 24160
rect 16485 24157 16497 24160
rect 16531 24157 16543 24191
rect 16485 24151 16543 24157
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24188 19855 24191
rect 20622 24188 20628 24200
rect 19843 24160 20628 24188
rect 19843 24157 19855 24160
rect 19797 24151 19855 24157
rect 20622 24148 20628 24160
rect 20680 24148 20686 24200
rect 17862 24120 17868 24132
rect 17775 24092 17868 24120
rect 17862 24080 17868 24092
rect 17920 24120 17926 24132
rect 17920 24092 18644 24120
rect 17920 24080 17926 24092
rect 18616 24064 18644 24092
rect 12529 24055 12587 24061
rect 12529 24021 12541 24055
rect 12575 24052 12587 24055
rect 12986 24052 12992 24064
rect 12575 24024 12992 24052
rect 12575 24021 12587 24024
rect 12529 24015 12587 24021
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 15746 24012 15752 24064
rect 15804 24052 15810 24064
rect 15841 24055 15899 24061
rect 15841 24052 15853 24055
rect 15804 24024 15853 24052
rect 15804 24012 15810 24024
rect 15841 24021 15853 24024
rect 15887 24021 15899 24055
rect 18598 24052 18604 24064
rect 18559 24024 18604 24052
rect 15841 24015 15899 24021
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 19426 24052 19432 24064
rect 19339 24024 19432 24052
rect 19426 24012 19432 24024
rect 19484 24052 19490 24064
rect 20530 24052 20536 24064
rect 19484 24024 20536 24052
rect 19484 24012 19490 24024
rect 20530 24012 20536 24024
rect 20588 24012 20594 24064
rect 24670 24012 24676 24064
rect 24728 24052 24734 24064
rect 24765 24055 24823 24061
rect 24765 24052 24777 24055
rect 24728 24024 24777 24052
rect 24728 24012 24734 24024
rect 24765 24021 24777 24024
rect 24811 24021 24823 24055
rect 24765 24015 24823 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 12066 23808 12072 23860
rect 12124 23848 12130 23860
rect 12161 23851 12219 23857
rect 12161 23848 12173 23851
rect 12124 23820 12173 23848
rect 12124 23808 12130 23820
rect 12161 23817 12173 23820
rect 12207 23817 12219 23851
rect 12161 23811 12219 23817
rect 12618 23808 12624 23860
rect 12676 23848 12682 23860
rect 13449 23851 13507 23857
rect 13449 23848 13461 23851
rect 12676 23820 13461 23848
rect 12676 23808 12682 23820
rect 13449 23817 13461 23820
rect 13495 23817 13507 23851
rect 13449 23811 13507 23817
rect 15930 23808 15936 23860
rect 15988 23848 15994 23860
rect 16025 23851 16083 23857
rect 16025 23848 16037 23851
rect 15988 23820 16037 23848
rect 15988 23808 15994 23820
rect 16025 23817 16037 23820
rect 16071 23817 16083 23851
rect 16025 23811 16083 23817
rect 19334 23808 19340 23860
rect 19392 23848 19398 23860
rect 19797 23851 19855 23857
rect 19797 23848 19809 23851
rect 19392 23820 19809 23848
rect 19392 23808 19398 23820
rect 19797 23817 19809 23820
rect 19843 23817 19855 23851
rect 21542 23848 21548 23860
rect 21503 23820 21548 23848
rect 19797 23811 19855 23817
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23290 23848 23296 23860
rect 22695 23820 23296 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 23474 23848 23480 23860
rect 23435 23820 23480 23848
rect 23474 23808 23480 23820
rect 23532 23808 23538 23860
rect 12986 23712 12992 23724
rect 12947 23684 12992 23712
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23712 15807 23715
rect 16666 23712 16672 23724
rect 15795 23684 16672 23712
rect 15795 23681 15807 23684
rect 15749 23675 15807 23681
rect 16666 23672 16672 23684
rect 16724 23712 16730 23724
rect 16761 23715 16819 23721
rect 16761 23712 16773 23715
rect 16724 23684 16773 23712
rect 16724 23672 16730 23684
rect 16761 23681 16773 23684
rect 16807 23712 16819 23715
rect 17221 23715 17279 23721
rect 17221 23712 17233 23715
rect 16807 23684 17233 23712
rect 16807 23681 16819 23684
rect 16761 23675 16819 23681
rect 17221 23681 17233 23684
rect 17267 23681 17279 23715
rect 18598 23712 18604 23724
rect 18559 23684 18604 23712
rect 17221 23675 17279 23681
rect 18598 23672 18604 23684
rect 18656 23672 18662 23724
rect 20898 23712 20904 23724
rect 20859 23684 20904 23712
rect 20898 23672 20904 23684
rect 20956 23672 20962 23724
rect 23492 23712 23520 23808
rect 23845 23715 23903 23721
rect 23845 23712 23857 23715
rect 23492 23684 23857 23712
rect 23845 23681 23857 23684
rect 23891 23681 23903 23715
rect 23845 23675 23903 23681
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12492 23616 12817 23644
rect 12492 23604 12498 23616
rect 12805 23613 12817 23616
rect 12851 23613 12863 23647
rect 12805 23607 12863 23613
rect 14001 23647 14059 23653
rect 14001 23613 14013 23647
rect 14047 23644 14059 23647
rect 14826 23644 14832 23656
rect 14047 23616 14832 23644
rect 14047 23613 14059 23616
rect 14001 23607 14059 23613
rect 14826 23604 14832 23616
rect 14884 23604 14890 23656
rect 16206 23604 16212 23656
rect 16264 23644 16270 23656
rect 16577 23647 16635 23653
rect 16577 23644 16589 23647
rect 16264 23616 16589 23644
rect 16264 23604 16270 23616
rect 16577 23613 16589 23616
rect 16623 23613 16635 23647
rect 16577 23607 16635 23613
rect 18138 23604 18144 23656
rect 18196 23644 18202 23656
rect 18417 23647 18475 23653
rect 18417 23644 18429 23647
rect 18196 23616 18429 23644
rect 18196 23604 18202 23616
rect 18417 23613 18429 23616
rect 18463 23613 18475 23647
rect 18417 23607 18475 23613
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 19613 23647 19671 23653
rect 19613 23644 19625 23647
rect 19484 23616 19625 23644
rect 19484 23604 19490 23616
rect 19613 23613 19625 23616
rect 19659 23644 19671 23647
rect 20165 23647 20223 23653
rect 20165 23644 20177 23647
rect 19659 23616 20177 23644
rect 19659 23613 19671 23616
rect 19613 23607 19671 23613
rect 20165 23613 20177 23616
rect 20211 23613 20223 23647
rect 20165 23607 20223 23613
rect 20806 23604 20812 23656
rect 20864 23644 20870 23656
rect 21361 23647 21419 23653
rect 21361 23644 21373 23647
rect 20864 23616 21373 23644
rect 20864 23604 20870 23616
rect 21361 23613 21373 23616
rect 21407 23644 21419 23647
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21407 23616 21925 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 21913 23607 21971 23613
rect 22465 23647 22523 23653
rect 22465 23613 22477 23647
rect 22511 23613 22523 23647
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 22465 23607 22523 23613
rect 23032 23616 23673 23644
rect 12066 23536 12072 23588
rect 12124 23576 12130 23588
rect 12526 23576 12532 23588
rect 12124 23548 12532 23576
rect 12124 23536 12130 23548
rect 12526 23536 12532 23548
rect 12584 23576 12590 23588
rect 12897 23579 12955 23585
rect 12897 23576 12909 23579
rect 12584 23548 12909 23576
rect 12584 23536 12590 23548
rect 12897 23545 12909 23548
rect 12943 23545 12955 23579
rect 12897 23539 12955 23545
rect 13909 23579 13967 23585
rect 13909 23545 13921 23579
rect 13955 23576 13967 23579
rect 14268 23579 14326 23585
rect 14268 23576 14280 23579
rect 13955 23548 14280 23576
rect 13955 23545 13967 23548
rect 13909 23539 13967 23545
rect 14268 23545 14280 23548
rect 14314 23576 14326 23579
rect 14366 23576 14372 23588
rect 14314 23548 14372 23576
rect 14314 23545 14326 23548
rect 14268 23539 14326 23545
rect 14366 23536 14372 23548
rect 14424 23536 14430 23588
rect 15930 23536 15936 23588
rect 15988 23576 15994 23588
rect 16114 23576 16120 23588
rect 15988 23548 16120 23576
rect 15988 23536 15994 23548
rect 16114 23536 16120 23548
rect 16172 23576 16178 23588
rect 16669 23579 16727 23585
rect 16669 23576 16681 23579
rect 16172 23548 16681 23576
rect 16172 23536 16178 23548
rect 16669 23545 16681 23548
rect 16715 23545 16727 23579
rect 18509 23579 18567 23585
rect 18509 23576 18521 23579
rect 16669 23539 16727 23545
rect 17788 23548 18521 23576
rect 17788 23520 17816 23548
rect 18509 23545 18521 23548
rect 18555 23576 18567 23579
rect 19978 23576 19984 23588
rect 18555 23548 19984 23576
rect 18555 23545 18567 23548
rect 18509 23539 18567 23545
rect 19978 23536 19984 23548
rect 20036 23536 20042 23588
rect 22480 23520 22508 23607
rect 8386 23468 8392 23520
rect 8444 23508 8450 23520
rect 9674 23508 9680 23520
rect 8444 23480 9680 23508
rect 8444 23468 8450 23480
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 12437 23511 12495 23517
rect 12437 23477 12449 23511
rect 12483 23508 12495 23511
rect 12802 23508 12808 23520
rect 12483 23480 12808 23508
rect 12483 23477 12495 23480
rect 12437 23471 12495 23477
rect 12802 23468 12808 23480
rect 12860 23468 12866 23520
rect 15381 23511 15439 23517
rect 15381 23477 15393 23511
rect 15427 23508 15439 23511
rect 15562 23508 15568 23520
rect 15427 23480 15568 23508
rect 15427 23477 15439 23480
rect 15381 23471 15439 23477
rect 15562 23468 15568 23480
rect 15620 23468 15626 23520
rect 16209 23511 16267 23517
rect 16209 23477 16221 23511
rect 16255 23508 16267 23511
rect 16482 23508 16488 23520
rect 16255 23480 16488 23508
rect 16255 23477 16267 23480
rect 16209 23471 16267 23477
rect 16482 23468 16488 23480
rect 16540 23468 16546 23520
rect 17770 23508 17776 23520
rect 17731 23480 17776 23508
rect 17770 23468 17776 23480
rect 17828 23468 17834 23520
rect 18046 23508 18052 23520
rect 18007 23480 18052 23508
rect 18046 23468 18052 23480
rect 18104 23468 18110 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 19061 23511 19119 23517
rect 19061 23508 19073 23511
rect 18748 23480 19073 23508
rect 18748 23468 18754 23480
rect 19061 23477 19073 23480
rect 19107 23477 19119 23511
rect 19518 23508 19524 23520
rect 19479 23480 19524 23508
rect 19061 23471 19119 23477
rect 19518 23468 19524 23480
rect 19576 23468 19582 23520
rect 22373 23511 22431 23517
rect 22373 23477 22385 23511
rect 22419 23508 22431 23511
rect 22462 23508 22468 23520
rect 22419 23480 22468 23508
rect 22419 23477 22431 23480
rect 22373 23471 22431 23477
rect 22462 23468 22468 23480
rect 22520 23468 22526 23520
rect 22646 23468 22652 23520
rect 22704 23508 22710 23520
rect 23032 23517 23060 23616
rect 23661 23613 23673 23616
rect 23707 23613 23719 23647
rect 23661 23607 23719 23613
rect 24949 23647 25007 23653
rect 24949 23613 24961 23647
rect 24995 23644 25007 23647
rect 24995 23616 25452 23644
rect 24995 23613 25007 23616
rect 24949 23607 25007 23613
rect 25424 23520 25452 23616
rect 23017 23511 23075 23517
rect 23017 23508 23029 23511
rect 22704 23480 23029 23508
rect 22704 23468 22710 23480
rect 23017 23477 23029 23480
rect 23063 23477 23075 23511
rect 23017 23471 23075 23477
rect 24118 23468 24124 23520
rect 24176 23508 24182 23520
rect 24581 23511 24639 23517
rect 24581 23508 24593 23511
rect 24176 23480 24593 23508
rect 24176 23468 24182 23480
rect 24581 23477 24593 23480
rect 24627 23477 24639 23511
rect 24581 23471 24639 23477
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 25133 23511 25191 23517
rect 25133 23508 25145 23511
rect 24912 23480 25145 23508
rect 24912 23468 24918 23480
rect 25133 23477 25145 23480
rect 25179 23477 25191 23511
rect 25133 23471 25191 23477
rect 25406 23468 25412 23520
rect 25464 23508 25470 23520
rect 25501 23511 25559 23517
rect 25501 23508 25513 23511
rect 25464 23480 25513 23508
rect 25464 23468 25470 23480
rect 25501 23477 25513 23480
rect 25547 23477 25559 23511
rect 25501 23471 25559 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 12897 23307 12955 23313
rect 12492 23276 12537 23304
rect 12492 23264 12498 23276
rect 12897 23273 12909 23307
rect 12943 23304 12955 23307
rect 14090 23304 14096 23316
rect 12943 23276 14096 23304
rect 12943 23273 12955 23276
rect 12897 23267 12955 23273
rect 11974 23100 11980 23112
rect 11935 23072 11980 23100
rect 11974 23060 11980 23072
rect 12032 23060 12038 23112
rect 12434 23060 12440 23112
rect 12492 23100 12498 23112
rect 12919 23100 12947 23267
rect 14090 23264 14096 23276
rect 14148 23304 14154 23316
rect 14826 23304 14832 23316
rect 14148 23276 14832 23304
rect 14148 23264 14154 23276
rect 14826 23264 14832 23276
rect 14884 23304 14890 23316
rect 15013 23307 15071 23313
rect 15013 23304 15025 23307
rect 14884 23276 15025 23304
rect 14884 23264 14890 23276
rect 15013 23273 15025 23276
rect 15059 23273 15071 23307
rect 15013 23267 15071 23273
rect 12986 23196 12992 23248
rect 13044 23236 13050 23248
rect 13234 23239 13292 23245
rect 13234 23236 13246 23239
rect 13044 23208 13246 23236
rect 13044 23196 13050 23208
rect 13234 23205 13246 23208
rect 13280 23205 13292 23239
rect 13234 23199 13292 23205
rect 15028 23168 15056 23267
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 16945 23307 17003 23313
rect 16945 23304 16957 23307
rect 16632 23276 16957 23304
rect 16632 23264 16638 23276
rect 16945 23273 16957 23276
rect 16991 23273 17003 23307
rect 16945 23267 17003 23273
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 21269 23307 21327 23313
rect 21269 23304 21281 23307
rect 20772 23276 21281 23304
rect 20772 23264 20778 23276
rect 21269 23273 21281 23276
rect 21315 23273 21327 23307
rect 21269 23267 21327 23273
rect 22741 23307 22799 23313
rect 22741 23273 22753 23307
rect 22787 23304 22799 23307
rect 23382 23304 23388 23316
rect 22787 23276 23388 23304
rect 22787 23273 22799 23276
rect 22741 23267 22799 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 17862 23245 17868 23248
rect 17313 23239 17371 23245
rect 17313 23236 17325 23239
rect 15304 23208 17325 23236
rect 15304 23177 15332 23208
rect 17313 23205 17325 23208
rect 17359 23205 17371 23239
rect 17856 23236 17868 23245
rect 17823 23208 17868 23236
rect 17313 23199 17371 23205
rect 17856 23199 17868 23208
rect 17862 23196 17868 23199
rect 17920 23196 17926 23248
rect 25222 23236 25228 23248
rect 25183 23208 25228 23236
rect 25222 23196 25228 23208
rect 25280 23196 25286 23248
rect 15562 23177 15568 23180
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 15028 23140 15301 23168
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15556 23168 15568 23177
rect 15523 23140 15568 23168
rect 15289 23131 15347 23137
rect 15556 23131 15568 23140
rect 15562 23128 15568 23131
rect 15620 23128 15626 23180
rect 17589 23171 17647 23177
rect 17589 23137 17601 23171
rect 17635 23168 17647 23171
rect 19337 23171 19395 23177
rect 19337 23168 19349 23171
rect 17635 23140 19349 23168
rect 17635 23137 17647 23140
rect 17589 23131 17647 23137
rect 19337 23137 19349 23140
rect 19383 23168 19395 23171
rect 19518 23168 19524 23180
rect 19383 23140 19524 23168
rect 19383 23137 19395 23140
rect 19337 23131 19395 23137
rect 19518 23128 19524 23140
rect 19576 23168 19582 23180
rect 19705 23171 19763 23177
rect 19705 23168 19717 23171
rect 19576 23140 19717 23168
rect 19576 23128 19582 23140
rect 19705 23137 19717 23140
rect 19751 23168 19763 23171
rect 20349 23171 20407 23177
rect 20349 23168 20361 23171
rect 19751 23140 20361 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 20349 23137 20361 23140
rect 20395 23168 20407 23171
rect 21266 23168 21272 23180
rect 20395 23140 21272 23168
rect 20395 23137 20407 23140
rect 20349 23131 20407 23137
rect 21266 23128 21272 23140
rect 21324 23128 21330 23180
rect 22557 23171 22615 23177
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 22830 23168 22836 23180
rect 22603 23140 22836 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 22830 23128 22836 23140
rect 22888 23128 22894 23180
rect 23661 23171 23719 23177
rect 23661 23137 23673 23171
rect 23707 23168 23719 23171
rect 23934 23168 23940 23180
rect 23707 23140 23940 23168
rect 23707 23137 23719 23140
rect 23661 23131 23719 23137
rect 23934 23128 23940 23140
rect 23992 23128 23998 23180
rect 24949 23171 25007 23177
rect 24949 23137 24961 23171
rect 24995 23168 25007 23171
rect 25038 23168 25044 23180
rect 24995 23140 25044 23168
rect 24995 23137 25007 23140
rect 24949 23131 25007 23137
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 12989 23103 13047 23109
rect 12989 23100 13001 23103
rect 12492 23072 13001 23100
rect 12492 23060 12498 23072
rect 12989 23069 13001 23072
rect 13035 23069 13047 23103
rect 12989 23063 13047 23069
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23100 19855 23103
rect 20622 23100 20628 23112
rect 19843 23072 20628 23100
rect 19843 23069 19855 23072
rect 19797 23063 19855 23069
rect 20622 23060 20628 23072
rect 20680 23060 20686 23112
rect 21358 23100 21364 23112
rect 21319 23072 21364 23100
rect 21358 23060 21364 23072
rect 21416 23060 21422 23112
rect 21453 23103 21511 23109
rect 21453 23069 21465 23103
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 16666 23032 16672 23044
rect 16627 23004 16672 23032
rect 16666 22992 16672 23004
rect 16724 22992 16730 23044
rect 21468 23032 21496 23063
rect 22370 23060 22376 23112
rect 22428 23100 22434 23112
rect 22465 23103 22523 23109
rect 22465 23100 22477 23103
rect 22428 23072 22477 23100
rect 22428 23060 22434 23072
rect 22465 23069 22477 23072
rect 22511 23100 22523 23103
rect 23845 23103 23903 23109
rect 23845 23100 23857 23103
rect 22511 23072 23857 23100
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 23845 23069 23857 23072
rect 23891 23069 23903 23103
rect 23845 23063 23903 23069
rect 21913 23035 21971 23041
rect 21913 23032 21925 23035
rect 20640 23004 21925 23032
rect 14366 22964 14372 22976
rect 14327 22936 14372 22964
rect 14366 22924 14372 22936
rect 14424 22924 14430 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 18969 22967 19027 22973
rect 18969 22964 18981 22967
rect 18932 22936 18981 22964
rect 18932 22924 18938 22936
rect 18969 22933 18981 22936
rect 19015 22933 19027 22967
rect 18969 22927 19027 22933
rect 20438 22924 20444 22976
rect 20496 22964 20502 22976
rect 20640 22973 20668 23004
rect 21913 23001 21925 23004
rect 21959 23001 21971 23035
rect 21913 22995 21971 23001
rect 20625 22967 20683 22973
rect 20625 22964 20637 22967
rect 20496 22936 20637 22964
rect 20496 22924 20502 22936
rect 20625 22933 20637 22936
rect 20671 22933 20683 22967
rect 20898 22964 20904 22976
rect 20859 22936 20904 22964
rect 20625 22927 20683 22933
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 14550 22720 14556 22772
rect 14608 22760 14614 22772
rect 14645 22763 14703 22769
rect 14645 22760 14657 22763
rect 14608 22732 14657 22760
rect 14608 22720 14614 22732
rect 14645 22729 14657 22732
rect 14691 22729 14703 22763
rect 14645 22723 14703 22729
rect 17681 22763 17739 22769
rect 17681 22729 17693 22763
rect 17727 22760 17739 22763
rect 17862 22760 17868 22772
rect 17727 22732 17868 22760
rect 17727 22729 17739 22732
rect 17681 22723 17739 22729
rect 10870 22584 10876 22636
rect 10928 22624 10934 22636
rect 11885 22627 11943 22633
rect 11885 22624 11897 22627
rect 10928 22596 11897 22624
rect 10928 22584 10934 22596
rect 11885 22593 11897 22596
rect 11931 22624 11943 22627
rect 12434 22624 12440 22636
rect 11931 22596 12440 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22624 14611 22627
rect 15197 22627 15255 22633
rect 15197 22624 15209 22627
rect 14599 22596 15209 22624
rect 14599 22593 14611 22596
rect 14553 22587 14611 22593
rect 15197 22593 15209 22596
rect 15243 22624 15255 22627
rect 15562 22624 15568 22636
rect 15243 22596 15568 22624
rect 15243 22593 15255 22596
rect 15197 22587 15255 22593
rect 15562 22584 15568 22596
rect 15620 22624 15626 22636
rect 15657 22627 15715 22633
rect 15657 22624 15669 22627
rect 15620 22596 15669 22624
rect 15620 22584 15626 22596
rect 15657 22593 15669 22596
rect 15703 22593 15715 22627
rect 15657 22587 15715 22593
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16632 22596 16865 22624
rect 16632 22584 16638 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 17034 22624 17040 22636
rect 16947 22596 17040 22624
rect 16853 22587 16911 22593
rect 17034 22584 17040 22596
rect 17092 22624 17098 22636
rect 17696 22624 17724 22723
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 20993 22763 21051 22769
rect 20993 22729 21005 22763
rect 21039 22760 21051 22763
rect 21082 22760 21088 22772
rect 21039 22732 21088 22760
rect 21039 22729 21051 22732
rect 20993 22723 21051 22729
rect 21082 22720 21088 22732
rect 21140 22760 21146 22772
rect 21358 22760 21364 22772
rect 21140 22732 21364 22760
rect 21140 22720 21146 22732
rect 21358 22720 21364 22732
rect 21416 22720 21422 22772
rect 24857 22763 24915 22769
rect 24857 22729 24869 22763
rect 24903 22760 24915 22763
rect 25038 22760 25044 22772
rect 24903 22732 25044 22760
rect 24903 22729 24915 22732
rect 24857 22723 24915 22729
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 17092 22596 17724 22624
rect 18325 22627 18383 22633
rect 17092 22584 17098 22596
rect 18325 22593 18337 22627
rect 18371 22624 18383 22627
rect 23937 22627 23995 22633
rect 18371 22596 19012 22624
rect 18371 22593 18383 22596
rect 18325 22587 18383 22593
rect 18230 22516 18236 22568
rect 18288 22556 18294 22568
rect 18984 22565 19012 22596
rect 23937 22593 23949 22627
rect 23983 22624 23995 22627
rect 24210 22624 24216 22636
rect 23983 22596 24216 22624
rect 23983 22593 23995 22596
rect 23937 22587 23995 22593
rect 24210 22584 24216 22596
rect 24268 22584 24274 22636
rect 18785 22559 18843 22565
rect 18785 22556 18797 22559
rect 18288 22528 18797 22556
rect 18288 22516 18294 22528
rect 18785 22525 18797 22528
rect 18831 22525 18843 22559
rect 18785 22519 18843 22525
rect 18969 22559 19027 22565
rect 18969 22525 18981 22559
rect 19015 22556 19027 22559
rect 19518 22556 19524 22568
rect 19015 22528 19524 22556
rect 19015 22525 19027 22528
rect 18969 22519 19027 22525
rect 12682 22491 12740 22497
rect 12682 22488 12694 22491
rect 12268 22460 12694 22488
rect 12268 22432 12296 22460
rect 12682 22457 12694 22460
rect 12728 22457 12740 22491
rect 14182 22488 14188 22500
rect 14095 22460 14188 22488
rect 12682 22451 12740 22457
rect 14182 22448 14188 22460
rect 14240 22488 14246 22500
rect 15013 22491 15071 22497
rect 15013 22488 15025 22491
rect 14240 22460 15025 22488
rect 14240 22448 14246 22460
rect 15013 22457 15025 22460
rect 15059 22457 15071 22491
rect 15013 22451 15071 22457
rect 16301 22491 16359 22497
rect 16301 22457 16313 22491
rect 16347 22488 16359 22491
rect 16761 22491 16819 22497
rect 16761 22488 16773 22491
rect 16347 22460 16773 22488
rect 16347 22457 16359 22460
rect 16301 22451 16359 22457
rect 16761 22457 16773 22460
rect 16807 22488 16819 22491
rect 16850 22488 16856 22500
rect 16807 22460 16856 22488
rect 16807 22457 16819 22460
rect 16761 22451 16819 22457
rect 16850 22448 16856 22460
rect 16908 22448 16914 22500
rect 18800 22488 18828 22519
rect 19518 22516 19524 22528
rect 19576 22516 19582 22568
rect 21177 22559 21235 22565
rect 21177 22525 21189 22559
rect 21223 22556 21235 22559
rect 21266 22556 21272 22568
rect 21223 22528 21272 22556
rect 21223 22525 21235 22528
rect 21177 22519 21235 22525
rect 21266 22516 21272 22528
rect 21324 22516 21330 22568
rect 22830 22556 22836 22568
rect 22791 22528 22836 22556
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 23661 22559 23719 22565
rect 23661 22525 23673 22559
rect 23707 22556 23719 22559
rect 24949 22559 25007 22565
rect 23707 22528 24440 22556
rect 23707 22525 23719 22528
rect 23661 22519 23719 22525
rect 18874 22488 18880 22500
rect 18787 22460 18880 22488
rect 18874 22448 18880 22460
rect 18932 22488 18938 22500
rect 19214 22491 19272 22497
rect 19214 22488 19226 22491
rect 18932 22460 19226 22488
rect 18932 22448 18938 22460
rect 19214 22457 19226 22460
rect 19260 22457 19272 22491
rect 21422 22491 21480 22497
rect 21422 22488 21434 22491
rect 19214 22451 19272 22457
rect 20456 22460 21434 22488
rect 20456 22432 20484 22460
rect 21422 22457 21434 22460
rect 21468 22457 21480 22491
rect 21422 22451 21480 22457
rect 24412 22432 24440 22528
rect 24949 22525 24961 22559
rect 24995 22556 25007 22559
rect 25038 22556 25044 22568
rect 24995 22528 25044 22556
rect 24995 22525 25007 22528
rect 24949 22519 25007 22525
rect 25038 22516 25044 22528
rect 25096 22556 25102 22568
rect 25501 22559 25559 22565
rect 25501 22556 25513 22559
rect 25096 22528 25513 22556
rect 25096 22516 25102 22528
rect 25501 22525 25513 22528
rect 25547 22525 25559 22559
rect 25501 22519 25559 22525
rect 12250 22420 12256 22432
rect 12211 22392 12256 22420
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 12986 22380 12992 22432
rect 13044 22420 13050 22432
rect 13817 22423 13875 22429
rect 13817 22420 13829 22423
rect 13044 22392 13829 22420
rect 13044 22380 13050 22392
rect 13817 22389 13829 22392
rect 13863 22389 13875 22423
rect 15102 22420 15108 22432
rect 15063 22392 15108 22420
rect 13817 22383 13875 22389
rect 15102 22380 15108 22392
rect 15160 22380 15166 22432
rect 16393 22423 16451 22429
rect 16393 22389 16405 22423
rect 16439 22420 16451 22423
rect 16482 22420 16488 22432
rect 16439 22392 16488 22420
rect 16439 22389 16451 22392
rect 16393 22383 16451 22389
rect 16482 22380 16488 22392
rect 16540 22380 16546 22432
rect 19518 22380 19524 22432
rect 19576 22420 19582 22432
rect 20349 22423 20407 22429
rect 20349 22420 20361 22423
rect 19576 22392 20361 22420
rect 19576 22380 19582 22392
rect 20349 22389 20361 22392
rect 20395 22420 20407 22423
rect 20438 22420 20444 22432
rect 20395 22392 20444 22420
rect 20395 22389 20407 22392
rect 20349 22383 20407 22389
rect 20438 22380 20444 22392
rect 20496 22380 20502 22432
rect 22554 22420 22560 22432
rect 22515 22392 22560 22420
rect 22554 22380 22560 22392
rect 22612 22380 22618 22432
rect 23477 22423 23535 22429
rect 23477 22389 23489 22423
rect 23523 22420 23535 22423
rect 23842 22420 23848 22432
rect 23523 22392 23848 22420
rect 23523 22389 23535 22392
rect 23477 22383 23535 22389
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 24394 22420 24400 22432
rect 24355 22392 24400 22420
rect 24394 22380 24400 22392
rect 24452 22380 24458 22432
rect 24854 22380 24860 22432
rect 24912 22420 24918 22432
rect 25133 22423 25191 22429
rect 25133 22420 25145 22423
rect 24912 22392 25145 22420
rect 24912 22380 24918 22392
rect 25133 22389 25145 22392
rect 25179 22389 25191 22423
rect 25133 22383 25191 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 10870 22216 10876 22228
rect 10831 22188 10876 22216
rect 10870 22176 10876 22188
rect 10928 22176 10934 22228
rect 12250 22176 12256 22228
rect 12308 22216 12314 22228
rect 12345 22219 12403 22225
rect 12345 22216 12357 22219
rect 12308 22188 12357 22216
rect 12308 22176 12314 22188
rect 12345 22185 12357 22188
rect 12391 22185 12403 22219
rect 12986 22216 12992 22228
rect 12947 22188 12992 22216
rect 12345 22179 12403 22185
rect 12986 22176 12992 22188
rect 13044 22176 13050 22228
rect 13633 22219 13691 22225
rect 13633 22185 13645 22219
rect 13679 22216 13691 22219
rect 14642 22216 14648 22228
rect 13679 22188 14648 22216
rect 13679 22185 13691 22188
rect 13633 22179 13691 22185
rect 14642 22176 14648 22188
rect 14700 22216 14706 22228
rect 15102 22216 15108 22228
rect 14700 22188 15108 22216
rect 14700 22176 14706 22188
rect 15102 22176 15108 22188
rect 15160 22176 15166 22228
rect 16761 22219 16819 22225
rect 16761 22185 16773 22219
rect 16807 22216 16819 22219
rect 17034 22216 17040 22228
rect 16807 22188 17040 22216
rect 16807 22185 16819 22188
rect 16761 22179 16819 22185
rect 17034 22176 17040 22188
rect 17092 22176 17098 22228
rect 18046 22216 18052 22228
rect 18007 22188 18052 22216
rect 18046 22176 18052 22188
rect 18104 22176 18110 22228
rect 20714 22216 20720 22228
rect 20675 22188 20720 22216
rect 20714 22176 20720 22188
rect 20772 22176 20778 22228
rect 24946 22176 24952 22228
rect 25004 22216 25010 22228
rect 25130 22216 25136 22228
rect 25004 22188 25136 22216
rect 25004 22176 25010 22188
rect 25130 22176 25136 22188
rect 25188 22176 25194 22228
rect 1394 22040 1400 22092
rect 1452 22080 1458 22092
rect 2314 22080 2320 22092
rect 1452 22052 2320 22080
rect 1452 22040 1458 22052
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 10888 22080 10916 22176
rect 14001 22151 14059 22157
rect 14001 22148 14013 22151
rect 13740 22120 14013 22148
rect 11238 22089 11244 22092
rect 10965 22083 11023 22089
rect 10965 22080 10977 22083
rect 10888 22052 10977 22080
rect 10965 22049 10977 22052
rect 11011 22049 11023 22083
rect 10965 22043 11023 22049
rect 11232 22043 11244 22089
rect 11296 22080 11302 22092
rect 11296 22052 11332 22080
rect 11238 22040 11244 22043
rect 11296 22040 11302 22052
rect 12802 22040 12808 22092
rect 12860 22080 12866 22092
rect 13449 22083 13507 22089
rect 13449 22080 13461 22083
rect 12860 22052 13461 22080
rect 12860 22040 12866 22052
rect 13449 22049 13461 22052
rect 13495 22049 13507 22083
rect 13449 22043 13507 22049
rect 13464 22012 13492 22043
rect 13538 22040 13544 22092
rect 13596 22080 13602 22092
rect 13740 22080 13768 22120
rect 14001 22117 14013 22120
rect 14047 22117 14059 22151
rect 18064 22148 18092 22176
rect 22554 22148 22560 22160
rect 14001 22111 14059 22117
rect 17880 22120 18092 22148
rect 22112 22120 22560 22148
rect 14642 22080 14648 22092
rect 13596 22052 13768 22080
rect 14603 22052 14648 22080
rect 13596 22040 13602 22052
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 16025 22083 16083 22089
rect 16025 22080 16037 22083
rect 15344 22052 16037 22080
rect 15344 22040 15350 22052
rect 16025 22049 16037 22052
rect 16071 22049 16083 22083
rect 16025 22043 16083 22049
rect 17589 22083 17647 22089
rect 17589 22049 17601 22083
rect 17635 22080 17647 22083
rect 17880 22080 17908 22120
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 17635 22052 17908 22080
rect 17972 22052 18153 22080
rect 17635 22049 17647 22052
rect 17589 22043 17647 22049
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13464 21984 14105 22012
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14277 22015 14335 22021
rect 14277 21981 14289 22015
rect 14323 22012 14335 22015
rect 14366 22012 14372 22024
rect 14323 21984 14372 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 14366 21972 14372 21984
rect 14424 22012 14430 22024
rect 14734 22012 14740 22024
rect 14424 21984 14740 22012
rect 14424 21972 14430 21984
rect 14734 21972 14740 21984
rect 14792 21972 14798 22024
rect 15562 21972 15568 22024
rect 15620 22012 15626 22024
rect 16117 22015 16175 22021
rect 16117 22012 16129 22015
rect 15620 21984 16129 22012
rect 15620 21972 15626 21984
rect 16117 21981 16129 21984
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 22012 16359 22015
rect 16482 22012 16488 22024
rect 16347 21984 16488 22012
rect 16347 21981 16359 21984
rect 16301 21975 16359 21981
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 17770 22012 17776 22024
rect 16632 21984 17776 22012
rect 16632 21972 16638 21984
rect 17770 21972 17776 21984
rect 17828 22012 17834 22024
rect 17972 22012 18000 22052
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 19610 22080 19616 22092
rect 19571 22052 19616 22080
rect 18141 22043 18199 22049
rect 19610 22040 19616 22052
rect 19668 22040 19674 22092
rect 20349 22083 20407 22089
rect 20349 22049 20361 22083
rect 20395 22080 20407 22083
rect 20898 22080 20904 22092
rect 20395 22052 20904 22080
rect 20395 22049 20407 22052
rect 20349 22043 20407 22049
rect 20898 22040 20904 22052
rect 20956 22040 20962 22092
rect 21174 22040 21180 22092
rect 21232 22080 21238 22092
rect 21352 22083 21410 22089
rect 21352 22080 21364 22083
rect 21232 22052 21364 22080
rect 21232 22040 21238 22052
rect 21352 22049 21364 22052
rect 21398 22080 21410 22083
rect 22112 22080 22140 22120
rect 22554 22108 22560 22120
rect 22612 22108 22618 22160
rect 23842 22080 23848 22092
rect 21398 22052 22140 22080
rect 23803 22052 23848 22080
rect 21398 22049 21410 22052
rect 21352 22043 21410 22049
rect 23842 22040 23848 22052
rect 23900 22040 23906 22092
rect 24121 22083 24179 22089
rect 24121 22049 24133 22083
rect 24167 22080 24179 22083
rect 24762 22080 24768 22092
rect 24167 22052 24768 22080
rect 24167 22049 24179 22052
rect 24121 22043 24179 22049
rect 24762 22040 24768 22052
rect 24820 22040 24826 22092
rect 25130 22080 25136 22092
rect 25091 22052 25136 22080
rect 25130 22040 25136 22052
rect 25188 22040 25194 22092
rect 25406 22080 25412 22092
rect 25367 22052 25412 22080
rect 25406 22040 25412 22052
rect 25464 22040 25470 22092
rect 18230 22012 18236 22024
rect 17828 21984 18000 22012
rect 18191 21984 18236 22012
rect 17828 21972 17834 21984
rect 18230 21972 18236 21984
rect 18288 21972 18294 22024
rect 19702 22012 19708 22024
rect 19663 21984 19708 22012
rect 19702 21972 19708 21984
rect 19760 21972 19766 22024
rect 19797 22015 19855 22021
rect 19797 21981 19809 22015
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 21085 22015 21143 22021
rect 21085 21981 21097 22015
rect 21131 21981 21143 22015
rect 21085 21975 21143 21981
rect 15105 21947 15163 21953
rect 15105 21913 15117 21947
rect 15151 21944 15163 21947
rect 17678 21944 17684 21956
rect 15151 21916 16344 21944
rect 17639 21916 17684 21944
rect 15151 21913 15163 21916
rect 15105 21907 15163 21913
rect 16316 21888 16344 21916
rect 17678 21904 17684 21916
rect 17736 21904 17742 21956
rect 19334 21904 19340 21956
rect 19392 21944 19398 21956
rect 19518 21944 19524 21956
rect 19392 21916 19524 21944
rect 19392 21904 19398 21916
rect 19518 21904 19524 21916
rect 19576 21944 19582 21956
rect 19812 21944 19840 21975
rect 19576 21916 19840 21944
rect 19576 21904 19582 21916
rect 10321 21879 10379 21885
rect 10321 21845 10333 21879
rect 10367 21876 10379 21879
rect 10686 21876 10692 21888
rect 10367 21848 10692 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 15565 21879 15623 21885
rect 15565 21845 15577 21879
rect 15611 21876 15623 21879
rect 15654 21876 15660 21888
rect 15611 21848 15660 21876
rect 15611 21845 15623 21848
rect 15565 21839 15623 21845
rect 15654 21836 15660 21848
rect 15712 21836 15718 21888
rect 16298 21836 16304 21888
rect 16356 21836 16362 21888
rect 18598 21836 18604 21888
rect 18656 21876 18662 21888
rect 18693 21879 18751 21885
rect 18693 21876 18705 21879
rect 18656 21848 18705 21876
rect 18656 21836 18662 21848
rect 18693 21845 18705 21848
rect 18739 21845 18751 21879
rect 18693 21839 18751 21845
rect 18874 21836 18880 21888
rect 18932 21876 18938 21888
rect 19061 21879 19119 21885
rect 19061 21876 19073 21879
rect 18932 21848 19073 21876
rect 18932 21836 18938 21848
rect 19061 21845 19073 21848
rect 19107 21845 19119 21879
rect 19061 21839 19119 21845
rect 19245 21879 19303 21885
rect 19245 21845 19257 21879
rect 19291 21876 19303 21879
rect 20346 21876 20352 21888
rect 19291 21848 20352 21876
rect 19291 21845 19303 21848
rect 19245 21839 19303 21845
rect 20346 21836 20352 21848
rect 20404 21836 20410 21888
rect 21100 21876 21128 21975
rect 24578 21904 24584 21956
rect 24636 21904 24642 21956
rect 21266 21876 21272 21888
rect 21100 21848 21272 21876
rect 21266 21836 21272 21848
rect 21324 21836 21330 21888
rect 22465 21879 22523 21885
rect 22465 21845 22477 21879
rect 22511 21876 22523 21879
rect 22554 21876 22560 21888
rect 22511 21848 22560 21876
rect 22511 21845 22523 21848
rect 22465 21839 22523 21845
rect 22554 21836 22560 21848
rect 22612 21836 22618 21888
rect 22738 21876 22744 21888
rect 22699 21848 22744 21876
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 24596 21876 24624 21904
rect 24670 21876 24676 21888
rect 24596 21848 24676 21876
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 10045 21675 10103 21681
rect 10045 21672 10057 21675
rect 9732 21644 10057 21672
rect 9732 21632 9738 21644
rect 10045 21641 10057 21644
rect 10091 21672 10103 21675
rect 11238 21672 11244 21684
rect 10091 21644 10640 21672
rect 11199 21644 11244 21672
rect 10091 21641 10103 21644
rect 10045 21635 10103 21641
rect 10226 21604 10232 21616
rect 10187 21576 10232 21604
rect 10226 21564 10232 21576
rect 10284 21564 10290 21616
rect 10612 21477 10640 21644
rect 11238 21632 11244 21644
rect 11296 21632 11302 21684
rect 14182 21672 14188 21684
rect 14143 21644 14188 21672
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 15286 21672 15292 21684
rect 15247 21644 15292 21672
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 15562 21632 15568 21684
rect 15620 21672 15626 21684
rect 15657 21675 15715 21681
rect 15657 21672 15669 21675
rect 15620 21644 15669 21672
rect 15620 21632 15626 21644
rect 15657 21641 15669 21644
rect 15703 21641 15715 21675
rect 15657 21635 15715 21641
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 18230 21672 18236 21684
rect 17543 21644 18236 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 18230 21632 18236 21644
rect 18288 21632 18294 21684
rect 19610 21632 19616 21684
rect 19668 21672 19674 21684
rect 19705 21675 19763 21681
rect 19705 21672 19717 21675
rect 19668 21644 19717 21672
rect 19668 21632 19674 21644
rect 19705 21641 19717 21644
rect 19751 21641 19763 21675
rect 23842 21672 23848 21684
rect 23803 21644 23848 21672
rect 19705 21635 19763 21641
rect 23842 21632 23848 21644
rect 23900 21632 23906 21684
rect 20438 21604 20444 21616
rect 20399 21576 20444 21604
rect 20438 21564 20444 21576
rect 20496 21564 20502 21616
rect 20622 21564 20628 21616
rect 20680 21604 20686 21616
rect 21453 21607 21511 21613
rect 21453 21604 21465 21607
rect 20680 21576 21465 21604
rect 20680 21564 20686 21576
rect 21453 21573 21465 21576
rect 21499 21604 21511 21607
rect 22002 21604 22008 21616
rect 21499 21576 22008 21604
rect 21499 21573 21511 21576
rect 21453 21567 21511 21573
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 25130 21604 25136 21616
rect 25091 21576 25136 21604
rect 25130 21564 25136 21576
rect 25188 21564 25194 21616
rect 10686 21496 10692 21548
rect 10744 21536 10750 21548
rect 10781 21539 10839 21545
rect 10781 21536 10793 21539
rect 10744 21508 10793 21536
rect 10744 21496 10750 21508
rect 10781 21505 10793 21508
rect 10827 21505 10839 21539
rect 12250 21536 12256 21548
rect 12211 21508 12256 21536
rect 10781 21499 10839 21505
rect 12250 21496 12256 21508
rect 12308 21536 12314 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12308 21508 13001 21536
rect 12308 21496 12314 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 14734 21536 14740 21548
rect 14695 21508 14740 21536
rect 12989 21499 13047 21505
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 15654 21496 15660 21548
rect 15712 21536 15718 21548
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 15712 21508 16313 21536
rect 15712 21496 15718 21508
rect 16301 21505 16313 21508
rect 16347 21505 16359 21539
rect 16301 21499 16359 21505
rect 16485 21539 16543 21545
rect 16485 21505 16497 21539
rect 16531 21536 16543 21539
rect 18874 21536 18880 21548
rect 16531 21508 16988 21536
rect 18835 21508 18880 21536
rect 16531 21505 16543 21508
rect 16485 21499 16543 21505
rect 10597 21471 10655 21477
rect 10597 21437 10609 21471
rect 10643 21437 10655 21471
rect 10597 21431 10655 21437
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 14642 21468 14648 21480
rect 14599 21440 14648 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 14642 21428 14648 21440
rect 14700 21428 14706 21480
rect 12805 21403 12863 21409
rect 12805 21400 12817 21403
rect 11808 21372 12817 21400
rect 10134 21292 10140 21344
rect 10192 21332 10198 21344
rect 10689 21335 10747 21341
rect 10689 21332 10701 21335
rect 10192 21304 10701 21332
rect 10192 21292 10198 21304
rect 10689 21301 10701 21304
rect 10735 21332 10747 21335
rect 10778 21332 10784 21344
rect 10735 21304 10784 21332
rect 10735 21301 10747 21304
rect 10689 21295 10747 21301
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11808 21341 11836 21372
rect 12805 21369 12817 21372
rect 12851 21369 12863 21403
rect 12805 21363 12863 21369
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11112 21304 11805 21332
rect 11112 21292 11118 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 12492 21304 12537 21332
rect 12492 21292 12498 21304
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 12897 21335 12955 21341
rect 12897 21332 12909 21335
rect 12768 21304 12909 21332
rect 12768 21292 12774 21304
rect 12897 21301 12909 21304
rect 12943 21301 12955 21335
rect 12897 21295 12955 21301
rect 13538 21292 13544 21344
rect 13596 21332 13602 21344
rect 13633 21335 13691 21341
rect 13633 21332 13645 21335
rect 13596 21304 13645 21332
rect 13596 21292 13602 21304
rect 13633 21301 13645 21304
rect 13679 21301 13691 21335
rect 13633 21295 13691 21301
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 14001 21335 14059 21341
rect 14001 21332 14013 21335
rect 13872 21304 14013 21332
rect 13872 21292 13878 21304
rect 14001 21301 14013 21304
rect 14047 21332 14059 21335
rect 14645 21335 14703 21341
rect 14645 21332 14657 21335
rect 14047 21304 14657 21332
rect 14047 21301 14059 21304
rect 14001 21295 14059 21301
rect 14645 21301 14657 21304
rect 14691 21332 14703 21335
rect 14826 21332 14832 21344
rect 14691 21304 14832 21332
rect 14691 21301 14703 21304
rect 14645 21295 14703 21301
rect 14826 21292 14832 21304
rect 14884 21292 14890 21344
rect 15838 21332 15844 21344
rect 15799 21304 15844 21332
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 16209 21335 16267 21341
rect 16209 21301 16221 21335
rect 16255 21332 16267 21335
rect 16298 21332 16304 21344
rect 16255 21304 16304 21332
rect 16255 21301 16267 21304
rect 16209 21295 16267 21301
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 16960 21341 16988 21508
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21536 19487 21539
rect 19518 21536 19524 21548
rect 19475 21508 19524 21536
rect 19475 21505 19487 21508
rect 19429 21499 19487 21505
rect 19518 21496 19524 21508
rect 19576 21536 19582 21548
rect 19702 21536 19708 21548
rect 19576 21508 19708 21536
rect 19576 21496 19582 21508
rect 19702 21496 19708 21508
rect 19760 21496 19766 21548
rect 20349 21539 20407 21545
rect 20349 21505 20361 21539
rect 20395 21536 20407 21539
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20395 21508 21097 21536
rect 20395 21505 20407 21508
rect 20349 21499 20407 21505
rect 21085 21505 21097 21508
rect 21131 21536 21143 21539
rect 21174 21536 21180 21548
rect 21131 21508 21180 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 21174 21496 21180 21508
rect 21232 21496 21238 21548
rect 22554 21536 22560 21548
rect 22515 21508 22560 21536
rect 22554 21496 22560 21508
rect 22612 21536 22618 21548
rect 23017 21539 23075 21545
rect 23017 21536 23029 21539
rect 22612 21508 23029 21536
rect 22612 21496 22618 21508
rect 23017 21505 23029 21508
rect 23063 21505 23075 21539
rect 23017 21499 23075 21505
rect 20809 21471 20867 21477
rect 20809 21437 20821 21471
rect 20855 21468 20867 21471
rect 20898 21468 20904 21480
rect 20855 21440 20904 21468
rect 20855 21437 20867 21440
rect 20809 21431 20867 21437
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 23934 21468 23940 21480
rect 23523 21440 23940 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 23934 21428 23940 21440
rect 23992 21468 23998 21480
rect 24213 21471 24271 21477
rect 24213 21468 24225 21471
rect 23992 21440 24225 21468
rect 23992 21428 23998 21440
rect 24213 21437 24225 21440
rect 24259 21437 24271 21471
rect 25498 21468 25504 21480
rect 25459 21440 25504 21468
rect 24213 21431 24271 21437
rect 25498 21428 25504 21440
rect 25556 21468 25562 21480
rect 26053 21471 26111 21477
rect 26053 21468 26065 21471
rect 25556 21440 26065 21468
rect 25556 21428 25562 21440
rect 26053 21437 26065 21440
rect 26099 21437 26111 21471
rect 26053 21431 26111 21437
rect 17865 21403 17923 21409
rect 17865 21369 17877 21403
rect 17911 21400 17923 21403
rect 18230 21400 18236 21412
rect 17911 21372 18236 21400
rect 17911 21369 17923 21372
rect 17865 21363 17923 21369
rect 18230 21360 18236 21372
rect 18288 21400 18294 21412
rect 18785 21403 18843 21409
rect 18785 21400 18797 21403
rect 18288 21372 18797 21400
rect 18288 21360 18294 21372
rect 18785 21369 18797 21372
rect 18831 21369 18843 21403
rect 18785 21363 18843 21369
rect 20990 21360 20996 21412
rect 21048 21400 21054 21412
rect 21821 21403 21879 21409
rect 21821 21400 21833 21403
rect 21048 21372 21833 21400
rect 21048 21360 21054 21372
rect 21821 21369 21833 21372
rect 21867 21400 21879 21403
rect 22465 21403 22523 21409
rect 22465 21400 22477 21403
rect 21867 21372 22477 21400
rect 21867 21369 21879 21372
rect 21821 21363 21879 21369
rect 22465 21369 22477 21372
rect 22511 21369 22523 21403
rect 24486 21400 24492 21412
rect 24447 21372 24492 21400
rect 22465 21363 22523 21369
rect 24486 21360 24492 21372
rect 24544 21360 24550 21412
rect 16945 21335 17003 21341
rect 16945 21301 16957 21335
rect 16991 21332 17003 21335
rect 17218 21332 17224 21344
rect 16991 21304 17224 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 18322 21332 18328 21344
rect 18283 21304 18328 21332
rect 18322 21292 18328 21304
rect 18380 21292 18386 21344
rect 18598 21292 18604 21344
rect 18656 21332 18662 21344
rect 18693 21335 18751 21341
rect 18693 21332 18705 21335
rect 18656 21304 18705 21332
rect 18656 21292 18662 21304
rect 18693 21301 18705 21304
rect 18739 21301 18751 21335
rect 18693 21295 18751 21301
rect 20346 21292 20352 21344
rect 20404 21332 20410 21344
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20404 21304 20913 21332
rect 20404 21292 20410 21304
rect 20901 21301 20913 21304
rect 20947 21301 20959 21335
rect 22002 21332 22008 21344
rect 21963 21304 22008 21332
rect 20901 21295 20959 21301
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 22373 21335 22431 21341
rect 22373 21332 22385 21335
rect 22152 21304 22385 21332
rect 22152 21292 22158 21304
rect 22373 21301 22385 21304
rect 22419 21301 22431 21335
rect 25682 21332 25688 21344
rect 25643 21304 25688 21332
rect 22373 21295 22431 21301
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 10870 21128 10876 21140
rect 10520 21100 10876 21128
rect 10520 21001 10548 21100
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 11238 21088 11244 21140
rect 11296 21128 11302 21140
rect 11885 21131 11943 21137
rect 11885 21128 11897 21131
rect 11296 21100 11897 21128
rect 11296 21088 11302 21100
rect 11885 21097 11897 21100
rect 11931 21097 11943 21131
rect 11885 21091 11943 21097
rect 12529 21131 12587 21137
rect 12529 21097 12541 21131
rect 12575 21128 12587 21131
rect 12710 21128 12716 21140
rect 12575 21100 12716 21128
rect 12575 21097 12587 21100
rect 12529 21091 12587 21097
rect 12710 21088 12716 21100
rect 12768 21088 12774 21140
rect 13170 21128 13176 21140
rect 13131 21100 13176 21128
rect 13170 21088 13176 21100
rect 13228 21088 13234 21140
rect 13817 21131 13875 21137
rect 13817 21097 13829 21131
rect 13863 21128 13875 21131
rect 14734 21128 14740 21140
rect 13863 21100 14740 21128
rect 13863 21097 13875 21100
rect 13817 21091 13875 21097
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 17770 21128 17776 21140
rect 17731 21100 17776 21128
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 19334 21128 19340 21140
rect 19295 21100 19340 21128
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 19889 21131 19947 21137
rect 19889 21097 19901 21131
rect 19935 21128 19947 21131
rect 20070 21128 20076 21140
rect 19935 21100 20076 21128
rect 19935 21097 19947 21100
rect 19889 21091 19947 21097
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 20346 21088 20352 21140
rect 20404 21128 20410 21140
rect 20441 21131 20499 21137
rect 20441 21128 20453 21131
rect 20404 21100 20453 21128
rect 20404 21088 20410 21100
rect 20441 21097 20453 21100
rect 20487 21097 20499 21131
rect 21174 21128 21180 21140
rect 21135 21100 21180 21128
rect 20441 21091 20499 21097
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 24026 21128 24032 21140
rect 23987 21100 24032 21128
rect 24026 21088 24032 21100
rect 24084 21088 24090 21140
rect 10686 21020 10692 21072
rect 10744 21069 10750 21072
rect 10744 21063 10808 21069
rect 10744 21029 10762 21063
rect 10796 21060 10808 21063
rect 11054 21060 11060 21072
rect 10796 21032 11060 21060
rect 10796 21029 10808 21032
rect 10744 21023 10808 21029
rect 10744 21020 10750 21023
rect 11054 21020 11060 21032
rect 11112 21020 11118 21072
rect 13998 21020 14004 21072
rect 14056 21060 14062 21072
rect 14642 21060 14648 21072
rect 14056 21032 14648 21060
rect 14056 21020 14062 21032
rect 14642 21020 14648 21032
rect 14700 21020 14706 21072
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20961 10563 20995
rect 13078 20992 13084 21004
rect 13039 20964 13084 20992
rect 10505 20955 10563 20961
rect 13078 20952 13084 20964
rect 13136 20952 13142 21004
rect 14458 20992 14464 21004
rect 14419 20964 14464 20992
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 15749 20995 15807 21001
rect 15749 20961 15761 20995
rect 15795 20992 15807 20995
rect 16108 20995 16166 21001
rect 16108 20992 16120 20995
rect 15795 20964 16120 20992
rect 15795 20961 15807 20964
rect 15749 20955 15807 20961
rect 16108 20961 16120 20964
rect 16154 20992 16166 20995
rect 16482 20992 16488 21004
rect 16154 20964 16488 20992
rect 16154 20961 16166 20964
rect 16108 20955 16166 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18417 20995 18475 21001
rect 18417 20992 18429 20995
rect 18012 20964 18429 20992
rect 18012 20952 18018 20964
rect 18417 20961 18429 20964
rect 18463 20961 18475 20995
rect 19426 20992 19432 21004
rect 18417 20955 18475 20961
rect 18524 20964 19432 20992
rect 13262 20924 13268 20936
rect 13223 20896 13268 20924
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 13630 20816 13636 20868
rect 13688 20856 13694 20868
rect 14182 20856 14188 20868
rect 13688 20828 14188 20856
rect 13688 20816 13694 20828
rect 14182 20816 14188 20828
rect 14240 20856 14246 20868
rect 14277 20859 14335 20865
rect 14277 20856 14289 20859
rect 14240 20828 14289 20856
rect 14240 20816 14246 20828
rect 14277 20825 14289 20828
rect 14323 20856 14335 20859
rect 15562 20856 15568 20868
rect 14323 20828 15568 20856
rect 14323 20825 14335 20828
rect 14277 20819 14335 20825
rect 15562 20816 15568 20828
rect 15620 20856 15626 20868
rect 15856 20856 15884 20887
rect 18138 20884 18144 20936
rect 18196 20924 18202 20936
rect 18524 20933 18552 20964
rect 19426 20952 19432 20964
rect 19484 20952 19490 21004
rect 19702 20992 19708 21004
rect 19663 20964 19708 20992
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 21266 20952 21272 21004
rect 21324 20992 21330 21004
rect 21726 21001 21732 21004
rect 21453 20995 21511 21001
rect 21453 20992 21465 20995
rect 21324 20964 21465 20992
rect 21324 20952 21330 20964
rect 21453 20961 21465 20964
rect 21499 20961 21511 20995
rect 21720 20992 21732 21001
rect 21687 20964 21732 20992
rect 21453 20955 21511 20961
rect 21720 20955 21732 20964
rect 21726 20952 21732 20955
rect 21784 20952 21790 21004
rect 25222 20992 25228 21004
rect 25183 20964 25228 20992
rect 25222 20952 25228 20964
rect 25280 20952 25286 21004
rect 18509 20927 18567 20933
rect 18509 20924 18521 20927
rect 18196 20896 18521 20924
rect 18196 20884 18202 20896
rect 18509 20893 18521 20896
rect 18555 20893 18567 20927
rect 18509 20887 18567 20893
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20924 18751 20927
rect 18874 20924 18880 20936
rect 18739 20896 18880 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 24026 20884 24032 20936
rect 24084 20924 24090 20936
rect 24121 20927 24179 20933
rect 24121 20924 24133 20927
rect 24084 20896 24133 20924
rect 24084 20884 24090 20896
rect 24121 20893 24133 20896
rect 24167 20893 24179 20927
rect 24121 20887 24179 20893
rect 24210 20884 24216 20936
rect 24268 20924 24274 20936
rect 24268 20896 24313 20924
rect 24268 20884 24274 20896
rect 15620 20828 15884 20856
rect 22833 20859 22891 20865
rect 15620 20816 15626 20828
rect 22833 20825 22845 20859
rect 22879 20856 22891 20859
rect 23661 20859 23719 20865
rect 22879 20828 23612 20856
rect 22879 20825 22891 20828
rect 22833 20819 22891 20825
rect 10321 20791 10379 20797
rect 10321 20757 10333 20791
rect 10367 20788 10379 20791
rect 10686 20788 10692 20800
rect 10367 20760 10692 20788
rect 10367 20757 10379 20760
rect 10321 20751 10379 20757
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 14093 20791 14151 20797
rect 14093 20788 14105 20791
rect 13964 20760 14105 20788
rect 13964 20748 13970 20760
rect 14093 20757 14105 20760
rect 14139 20757 14151 20791
rect 17218 20788 17224 20800
rect 17179 20760 17224 20788
rect 14093 20751 14151 20757
rect 17218 20748 17224 20760
rect 17276 20748 17282 20800
rect 18046 20788 18052 20800
rect 18007 20760 18052 20788
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 22370 20748 22376 20800
rect 22428 20788 22434 20800
rect 22738 20788 22744 20800
rect 22428 20760 22744 20788
rect 22428 20748 22434 20760
rect 22738 20748 22744 20760
rect 22796 20788 22802 20800
rect 23109 20791 23167 20797
rect 23109 20788 23121 20791
rect 22796 20760 23121 20788
rect 22796 20748 22802 20760
rect 23109 20757 23121 20760
rect 23155 20788 23167 20791
rect 23477 20791 23535 20797
rect 23477 20788 23489 20791
rect 23155 20760 23489 20788
rect 23155 20757 23167 20760
rect 23109 20751 23167 20757
rect 23477 20757 23489 20760
rect 23523 20757 23535 20791
rect 23584 20788 23612 20828
rect 23661 20825 23673 20859
rect 23707 20856 23719 20859
rect 24946 20856 24952 20868
rect 23707 20828 24952 20856
rect 23707 20825 23719 20828
rect 23661 20819 23719 20825
rect 24946 20816 24952 20828
rect 25004 20816 25010 20868
rect 24210 20788 24216 20800
rect 23584 20760 24216 20788
rect 23477 20751 23535 20757
rect 24210 20748 24216 20760
rect 24268 20748 24274 20800
rect 24762 20748 24768 20800
rect 24820 20788 24826 20800
rect 25409 20791 25467 20797
rect 25409 20788 25421 20791
rect 24820 20760 25421 20788
rect 24820 20748 24826 20760
rect 25409 20757 25421 20760
rect 25455 20757 25467 20791
rect 25409 20751 25467 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 9398 20584 9404 20596
rect 9359 20556 9404 20584
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 10962 20584 10968 20596
rect 10827 20556 10968 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11514 20584 11520 20596
rect 11112 20556 11520 20584
rect 11112 20544 11118 20556
rect 11514 20544 11520 20556
rect 11572 20584 11578 20596
rect 11793 20587 11851 20593
rect 11793 20584 11805 20587
rect 11572 20556 11805 20584
rect 11572 20544 11578 20556
rect 11793 20553 11805 20556
rect 11839 20553 11851 20587
rect 11793 20547 11851 20553
rect 11882 20544 11888 20596
rect 11940 20584 11946 20596
rect 15286 20584 15292 20596
rect 11940 20556 15292 20584
rect 11940 20544 11946 20556
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15565 20587 15623 20593
rect 15565 20553 15577 20587
rect 15611 20584 15623 20587
rect 16482 20584 16488 20596
rect 15611 20556 16488 20584
rect 15611 20553 15623 20556
rect 15565 20547 15623 20553
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 17497 20587 17555 20593
rect 17497 20553 17509 20587
rect 17543 20584 17555 20587
rect 17862 20584 17868 20596
rect 17543 20556 17868 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 18414 20584 18420 20596
rect 18279 20556 18420 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 18414 20544 18420 20556
rect 18472 20544 18478 20596
rect 21266 20544 21272 20596
rect 21324 20584 21330 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 21324 20556 21373 20584
rect 21324 20544 21330 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 22002 20584 22008 20596
rect 21963 20556 22008 20584
rect 21361 20547 21419 20553
rect 22002 20544 22008 20556
rect 22060 20544 22066 20596
rect 25038 20584 25044 20596
rect 24999 20556 25044 20584
rect 25038 20544 25044 20556
rect 25096 20544 25102 20596
rect 25222 20544 25228 20596
rect 25280 20584 25286 20596
rect 25961 20587 26019 20593
rect 25961 20584 25973 20587
rect 25280 20556 25973 20584
rect 25280 20544 25286 20556
rect 25961 20553 25973 20556
rect 26007 20553 26019 20587
rect 25961 20547 26019 20553
rect 17037 20519 17095 20525
rect 17037 20516 17049 20519
rect 16500 20488 17049 20516
rect 9766 20448 9772 20460
rect 9727 20420 9772 20448
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 11238 20408 11244 20460
rect 11296 20448 11302 20460
rect 11333 20451 11391 20457
rect 11333 20448 11345 20451
rect 11296 20420 11345 20448
rect 11296 20408 11302 20420
rect 11333 20417 11345 20420
rect 11379 20448 11391 20451
rect 12161 20451 12219 20457
rect 12161 20448 12173 20451
rect 11379 20420 12173 20448
rect 11379 20417 11391 20420
rect 11333 20411 11391 20417
rect 12161 20417 12173 20420
rect 12207 20448 12219 20451
rect 13262 20448 13268 20460
rect 12207 20420 13268 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13630 20448 13636 20460
rect 13591 20420 13636 20448
rect 13630 20408 13636 20420
rect 13688 20408 13694 20460
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16500 20457 16528 20488
rect 17037 20485 17049 20488
rect 17083 20485 17095 20519
rect 17037 20479 17095 20485
rect 21910 20476 21916 20528
rect 21968 20516 21974 20528
rect 23477 20519 23535 20525
rect 23477 20516 23489 20519
rect 21968 20488 23489 20516
rect 21968 20476 21974 20488
rect 23477 20485 23489 20488
rect 23523 20516 23535 20519
rect 23523 20488 24164 20516
rect 23523 20485 23535 20488
rect 23477 20479 23535 20485
rect 16485 20451 16543 20457
rect 16485 20448 16497 20451
rect 15896 20420 16497 20448
rect 15896 20408 15902 20420
rect 16485 20417 16497 20420
rect 16531 20417 16543 20451
rect 16485 20411 16543 20417
rect 16577 20451 16635 20457
rect 16577 20417 16589 20451
rect 16623 20417 16635 20451
rect 16577 20411 16635 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 21177 20451 21235 20457
rect 21177 20448 21189 20451
rect 20947 20420 21189 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 21177 20417 21189 20420
rect 21223 20448 21235 20451
rect 21726 20448 21732 20460
rect 21223 20420 21732 20448
rect 21223 20417 21235 20420
rect 21177 20411 21235 20417
rect 9398 20340 9404 20392
rect 9456 20380 9462 20392
rect 13906 20389 13912 20392
rect 9493 20383 9551 20389
rect 9493 20380 9505 20383
rect 9456 20352 9505 20380
rect 9456 20340 9462 20352
rect 9493 20349 9505 20352
rect 9539 20349 9551 20383
rect 13900 20380 13912 20389
rect 13867 20352 13912 20380
rect 9493 20343 9551 20349
rect 13900 20343 13912 20352
rect 13964 20380 13970 20392
rect 15933 20383 15991 20389
rect 15933 20380 15945 20383
rect 13964 20352 15945 20380
rect 13906 20340 13912 20343
rect 13964 20340 13970 20352
rect 15933 20349 15945 20352
rect 15979 20380 15991 20383
rect 16592 20380 16620 20411
rect 21726 20408 21732 20420
rect 21784 20448 21790 20460
rect 22554 20448 22560 20460
rect 21784 20420 22560 20448
rect 21784 20408 21790 20420
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 24136 20457 24164 20488
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 24213 20451 24271 20457
rect 24213 20417 24225 20451
rect 24259 20417 24271 20451
rect 25406 20448 25412 20460
rect 25367 20420 25412 20448
rect 24213 20411 24271 20417
rect 16942 20380 16948 20392
rect 15979 20352 16948 20380
rect 15979 20349 15991 20352
rect 15933 20343 15991 20349
rect 16942 20340 16948 20352
rect 17000 20340 17006 20392
rect 18049 20383 18107 20389
rect 18049 20349 18061 20383
rect 18095 20380 18107 20383
rect 19150 20380 19156 20392
rect 18095 20352 18736 20380
rect 19111 20352 19156 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 10321 20315 10379 20321
rect 10321 20281 10333 20315
rect 10367 20312 10379 20315
rect 11149 20315 11207 20321
rect 11149 20312 11161 20315
rect 10367 20284 11161 20312
rect 10367 20281 10379 20284
rect 10321 20275 10379 20281
rect 11149 20281 11161 20284
rect 11195 20312 11207 20315
rect 12437 20315 12495 20321
rect 12437 20312 12449 20315
rect 11195 20284 12449 20312
rect 11195 20281 11207 20284
rect 11149 20275 11207 20281
rect 12437 20281 12449 20284
rect 12483 20281 12495 20315
rect 16574 20312 16580 20324
rect 12437 20275 12495 20281
rect 16040 20284 16580 20312
rect 9858 20204 9864 20256
rect 9916 20244 9922 20256
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 9916 20216 10609 20244
rect 9916 20204 9922 20216
rect 10597 20213 10609 20216
rect 10643 20244 10655 20247
rect 11238 20244 11244 20256
rect 10643 20216 11244 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 11238 20204 11244 20216
rect 11296 20204 11302 20256
rect 12989 20247 13047 20253
rect 12989 20213 13001 20247
rect 13035 20244 13047 20247
rect 13078 20244 13084 20256
rect 13035 20216 13084 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13078 20204 13084 20216
rect 13136 20244 13142 20256
rect 14734 20244 14740 20256
rect 13136 20216 14740 20244
rect 13136 20204 13142 20216
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 16040 20253 16068 20284
rect 16574 20272 16580 20284
rect 16632 20272 16638 20324
rect 15013 20247 15071 20253
rect 15013 20244 15025 20247
rect 14884 20216 15025 20244
rect 14884 20204 14890 20216
rect 15013 20213 15025 20216
rect 15059 20213 15071 20247
rect 15013 20207 15071 20213
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20213 16083 20247
rect 16390 20244 16396 20256
rect 16351 20216 16396 20244
rect 16025 20207 16083 20213
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 17773 20247 17831 20253
rect 17773 20244 17785 20247
rect 16816 20216 17785 20244
rect 16816 20204 16822 20216
rect 17773 20213 17785 20216
rect 17819 20244 17831 20247
rect 18138 20244 18144 20256
rect 17819 20216 18144 20244
rect 17819 20213 17831 20216
rect 17773 20207 17831 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18708 20253 18736 20352
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 21545 20383 21603 20389
rect 21545 20380 21557 20383
rect 20772 20352 21557 20380
rect 20772 20340 20778 20352
rect 21545 20349 21557 20352
rect 21591 20349 21603 20383
rect 21545 20343 21603 20349
rect 21637 20383 21695 20389
rect 21637 20349 21649 20383
rect 21683 20380 21695 20383
rect 22465 20383 22523 20389
rect 22465 20380 22477 20383
rect 21683 20352 22477 20380
rect 21683 20349 21695 20352
rect 21637 20343 21695 20349
rect 22465 20349 22477 20352
rect 22511 20349 22523 20383
rect 22465 20343 22523 20349
rect 23658 20340 23664 20392
rect 23716 20380 23722 20392
rect 24228 20380 24256 20411
rect 25406 20408 25412 20420
rect 25464 20408 25470 20460
rect 24578 20380 24584 20392
rect 23716 20352 24584 20380
rect 23716 20340 23722 20352
rect 24578 20340 24584 20352
rect 24636 20380 24642 20392
rect 24673 20383 24731 20389
rect 24673 20380 24685 20383
rect 24636 20352 24685 20380
rect 24636 20340 24642 20352
rect 24673 20349 24685 20352
rect 24719 20349 24731 20383
rect 24673 20343 24731 20349
rect 24946 20340 24952 20392
rect 25004 20380 25010 20392
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 25004 20352 25237 20380
rect 25004 20340 25010 20352
rect 25225 20349 25237 20352
rect 25271 20349 25283 20383
rect 25225 20343 25283 20349
rect 19058 20312 19064 20324
rect 18971 20284 19064 20312
rect 19058 20272 19064 20284
rect 19116 20312 19122 20324
rect 19398 20315 19456 20321
rect 19398 20312 19410 20315
rect 19116 20284 19410 20312
rect 19116 20272 19122 20284
rect 19398 20281 19410 20284
rect 19444 20281 19456 20315
rect 19398 20275 19456 20281
rect 21266 20272 21272 20324
rect 21324 20312 21330 20324
rect 22278 20312 22284 20324
rect 21324 20284 22284 20312
rect 21324 20272 21330 20284
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 24029 20315 24087 20321
rect 24029 20312 24041 20315
rect 23032 20284 24041 20312
rect 23032 20256 23060 20284
rect 24029 20281 24041 20284
rect 24075 20281 24087 20315
rect 24029 20275 24087 20281
rect 18693 20247 18751 20253
rect 18693 20213 18705 20247
rect 18739 20244 18751 20247
rect 18782 20244 18788 20256
rect 18739 20216 18788 20244
rect 18739 20213 18751 20216
rect 18693 20207 18751 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 20533 20247 20591 20253
rect 20533 20244 20545 20247
rect 18932 20216 20545 20244
rect 18932 20204 18938 20216
rect 20533 20213 20545 20216
rect 20579 20213 20591 20247
rect 20533 20207 20591 20213
rect 21082 20204 21088 20256
rect 21140 20244 21146 20256
rect 21637 20247 21695 20253
rect 21637 20244 21649 20247
rect 21140 20216 21649 20244
rect 21140 20204 21146 20216
rect 21637 20213 21649 20216
rect 21683 20244 21695 20247
rect 21821 20247 21879 20253
rect 21821 20244 21833 20247
rect 21683 20216 21833 20244
rect 21683 20213 21695 20216
rect 21637 20207 21695 20213
rect 21821 20213 21833 20216
rect 21867 20213 21879 20247
rect 21821 20207 21879 20213
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 22373 20247 22431 20253
rect 22373 20244 22385 20247
rect 22152 20216 22385 20244
rect 22152 20204 22158 20216
rect 22373 20213 22385 20216
rect 22419 20213 22431 20247
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 22373 20207 22431 20213
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 23658 20244 23664 20256
rect 23619 20216 23664 20244
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 11514 20040 11520 20052
rect 11475 20012 11520 20040
rect 11514 20000 11520 20012
rect 11572 20000 11578 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13170 20040 13176 20052
rect 12851 20012 13176 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 14458 20000 14464 20052
rect 14516 20040 14522 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 14516 20012 15025 20040
rect 14516 20000 14522 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 16390 20000 16396 20052
rect 16448 20040 16454 20052
rect 17221 20043 17279 20049
rect 17221 20040 17233 20043
rect 16448 20012 17233 20040
rect 16448 20000 16454 20012
rect 17221 20009 17233 20012
rect 17267 20040 17279 20043
rect 17773 20043 17831 20049
rect 17773 20040 17785 20043
rect 17267 20012 17785 20040
rect 17267 20009 17279 20012
rect 17221 20003 17279 20009
rect 17773 20009 17785 20012
rect 17819 20009 17831 20043
rect 17773 20003 17831 20009
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18141 20043 18199 20049
rect 18141 20040 18153 20043
rect 18104 20012 18153 20040
rect 18104 20000 18110 20012
rect 18141 20009 18153 20012
rect 18187 20009 18199 20043
rect 18141 20003 18199 20009
rect 18233 20043 18291 20049
rect 18233 20009 18245 20043
rect 18279 20040 18291 20043
rect 18322 20040 18328 20052
rect 18279 20012 18328 20040
rect 18279 20009 18291 20012
rect 18233 20003 18291 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18874 20040 18880 20052
rect 18835 20012 18880 20040
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 20070 20040 20076 20052
rect 19935 20012 20076 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 20346 20040 20352 20052
rect 20307 20012 20352 20040
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20714 20040 20720 20052
rect 20675 20012 20720 20040
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 23661 20043 23719 20049
rect 23661 20009 23673 20043
rect 23707 20040 23719 20043
rect 24026 20040 24032 20052
rect 23707 20012 24032 20040
rect 23707 20009 23719 20012
rect 23661 20003 23719 20009
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 24305 20043 24363 20049
rect 24305 20040 24317 20043
rect 24176 20012 24317 20040
rect 24176 20000 24182 20012
rect 24305 20009 24317 20012
rect 24351 20009 24363 20043
rect 24305 20003 24363 20009
rect 24946 20000 24952 20052
rect 25004 20040 25010 20052
rect 25501 20043 25559 20049
rect 25501 20040 25513 20043
rect 25004 20012 25513 20040
rect 25004 20000 25010 20012
rect 25501 20009 25513 20012
rect 25547 20009 25559 20043
rect 25501 20003 25559 20009
rect 10045 19975 10103 19981
rect 10045 19941 10057 19975
rect 10091 19972 10103 19975
rect 10870 19972 10876 19984
rect 10091 19944 10876 19972
rect 10091 19941 10103 19944
rect 10045 19935 10103 19941
rect 10152 19913 10180 19944
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 12069 19975 12127 19981
rect 12069 19941 12081 19975
rect 12115 19972 12127 19975
rect 12437 19975 12495 19981
rect 12437 19972 12449 19975
rect 12115 19944 12449 19972
rect 12115 19941 12127 19944
rect 12069 19935 12127 19941
rect 12437 19941 12449 19944
rect 12483 19972 12495 19975
rect 13630 19972 13636 19984
rect 12483 19944 13636 19972
rect 12483 19941 12495 19944
rect 12437 19935 12495 19941
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 10226 19864 10232 19916
rect 10284 19904 10290 19916
rect 10393 19907 10451 19913
rect 10393 19904 10405 19907
rect 10284 19876 10405 19904
rect 10284 19864 10290 19876
rect 10393 19873 10405 19876
rect 10439 19873 10451 19907
rect 10393 19867 10451 19873
rect 12728 19836 12756 19944
rect 13630 19932 13636 19944
rect 13688 19932 13694 19984
rect 17589 19975 17647 19981
rect 17589 19972 17601 19975
rect 15571 19944 17601 19972
rect 15571 19916 15599 19944
rect 17589 19941 17601 19944
rect 17635 19941 17647 19975
rect 17589 19935 17647 19941
rect 24857 19975 24915 19981
rect 24857 19941 24869 19975
rect 24903 19972 24915 19975
rect 25314 19972 25320 19984
rect 24903 19944 25320 19972
rect 24903 19941 24915 19944
rect 24857 19935 24915 19941
rect 25314 19932 25320 19944
rect 25372 19932 25378 19984
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 13153 19907 13211 19913
rect 13153 19904 13165 19907
rect 12860 19876 13165 19904
rect 12860 19864 12866 19876
rect 13153 19873 13165 19876
rect 13199 19904 13211 19907
rect 14826 19904 14832 19916
rect 13199 19876 14832 19904
rect 13199 19873 13211 19876
rect 13153 19867 13211 19873
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 15562 19904 15568 19916
rect 15523 19876 15568 19904
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 15821 19907 15879 19913
rect 15821 19904 15833 19907
rect 15712 19876 15833 19904
rect 15712 19864 15718 19876
rect 15821 19873 15833 19876
rect 15867 19873 15879 19907
rect 19702 19904 19708 19916
rect 19663 19876 19708 19904
rect 15821 19867 15879 19873
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 21177 19907 21235 19913
rect 21177 19873 21189 19907
rect 21223 19904 21235 19907
rect 21266 19904 21272 19916
rect 21223 19876 21272 19904
rect 21223 19873 21235 19876
rect 21177 19867 21235 19873
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 22370 19864 22376 19916
rect 22428 19904 22434 19916
rect 22548 19907 22606 19913
rect 22548 19904 22560 19907
rect 22428 19876 22560 19904
rect 22428 19864 22434 19876
rect 22548 19873 22560 19876
rect 22594 19904 22606 19907
rect 24029 19907 24087 19913
rect 24029 19904 24041 19907
rect 22594 19876 24041 19904
rect 22594 19873 22606 19876
rect 22548 19867 22606 19873
rect 24029 19873 24041 19876
rect 24075 19904 24087 19907
rect 24210 19904 24216 19916
rect 24075 19876 24216 19904
rect 24075 19873 24087 19876
rect 24029 19867 24087 19873
rect 24210 19864 24216 19876
rect 24268 19864 24274 19916
rect 24946 19904 24952 19916
rect 24907 19876 24952 19904
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 12897 19839 12955 19845
rect 12897 19836 12909 19839
rect 12728 19808 12909 19836
rect 12897 19805 12909 19808
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 18138 19796 18144 19848
rect 18196 19836 18202 19848
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 18196 19808 18337 19836
rect 18196 19796 18202 19808
rect 18325 19805 18337 19808
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 19208 19808 19625 19836
rect 19208 19796 19214 19808
rect 19613 19805 19625 19808
rect 19659 19836 19671 19839
rect 22278 19836 22284 19848
rect 19659 19808 22284 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 24578 19796 24584 19848
rect 24636 19836 24642 19848
rect 25041 19839 25099 19845
rect 25041 19836 25053 19839
rect 24636 19808 25053 19836
rect 24636 19796 24642 19808
rect 25041 19805 25053 19808
rect 25087 19836 25099 19839
rect 25958 19836 25964 19848
rect 25087 19808 25964 19836
rect 25087 19805 25099 19808
rect 25041 19799 25099 19805
rect 25958 19796 25964 19808
rect 26016 19796 26022 19848
rect 13906 19728 13912 19780
rect 13964 19768 13970 19780
rect 14645 19771 14703 19777
rect 14645 19768 14657 19771
rect 13964 19740 14657 19768
rect 13964 19728 13970 19740
rect 14645 19737 14657 19740
rect 14691 19737 14703 19771
rect 16942 19768 16948 19780
rect 16903 19740 16948 19768
rect 14645 19731 14703 19737
rect 16942 19728 16948 19740
rect 17000 19728 17006 19780
rect 23474 19728 23480 19780
rect 23532 19768 23538 19780
rect 24489 19771 24547 19777
rect 24489 19768 24501 19771
rect 23532 19740 24501 19768
rect 23532 19728 23538 19740
rect 24489 19737 24501 19740
rect 24535 19737 24547 19771
rect 24489 19731 24547 19737
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 14240 19672 14289 19700
rect 14240 19660 14246 19672
rect 14277 19669 14289 19672
rect 14323 19669 14335 19703
rect 14277 19663 14335 19669
rect 19245 19703 19303 19709
rect 19245 19669 19257 19703
rect 19291 19700 19303 19703
rect 19334 19700 19340 19712
rect 19291 19672 19340 19700
rect 19291 19669 19303 19672
rect 19245 19663 19303 19669
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 22152 19672 22197 19700
rect 22152 19660 22158 19672
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 10597 19499 10655 19505
rect 10597 19465 10609 19499
rect 10643 19496 10655 19499
rect 10870 19496 10876 19508
rect 10643 19468 10876 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 10870 19456 10876 19468
rect 10928 19496 10934 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 10928 19468 11805 19496
rect 10928 19456 10934 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 11793 19459 11851 19465
rect 12253 19499 12311 19505
rect 12253 19465 12265 19499
rect 12299 19496 12311 19499
rect 12802 19496 12808 19508
rect 12299 19468 12808 19496
rect 12299 19465 12311 19468
rect 12253 19459 12311 19465
rect 290 19320 296 19372
rect 348 19360 354 19372
rect 382 19360 388 19372
rect 348 19332 388 19360
rect 348 19320 354 19332
rect 382 19320 388 19332
rect 440 19320 446 19372
rect 11808 19360 11836 19459
rect 12802 19456 12808 19468
rect 12860 19496 12866 19508
rect 14093 19499 14151 19505
rect 14093 19496 14105 19499
rect 12860 19468 14105 19496
rect 12860 19456 12866 19468
rect 14093 19465 14105 19468
rect 14139 19465 14151 19499
rect 15286 19496 15292 19508
rect 14093 19459 14151 19465
rect 14384 19468 15292 19496
rect 14277 19431 14335 19437
rect 14277 19397 14289 19431
rect 14323 19428 14335 19431
rect 14384 19428 14412 19468
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 17126 19456 17132 19508
rect 17184 19496 17190 19508
rect 17402 19496 17408 19508
rect 17184 19468 17408 19496
rect 17184 19456 17190 19468
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 18322 19456 18328 19508
rect 18380 19496 18386 19508
rect 18509 19499 18567 19505
rect 18509 19496 18521 19499
rect 18380 19468 18521 19496
rect 18380 19456 18386 19468
rect 18509 19465 18521 19468
rect 18555 19465 18567 19499
rect 18509 19459 18567 19465
rect 21913 19499 21971 19505
rect 21913 19465 21925 19499
rect 21959 19496 21971 19499
rect 22370 19496 22376 19508
rect 21959 19468 22376 19496
rect 21959 19465 21971 19468
rect 21913 19459 21971 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 24670 19456 24676 19508
rect 24728 19496 24734 19508
rect 24765 19499 24823 19505
rect 24765 19496 24777 19499
rect 24728 19468 24777 19496
rect 24728 19456 24734 19468
rect 24765 19465 24777 19468
rect 24811 19496 24823 19499
rect 24946 19496 24952 19508
rect 24811 19468 24952 19496
rect 24811 19465 24823 19468
rect 24765 19459 24823 19465
rect 24946 19456 24952 19468
rect 25004 19456 25010 19508
rect 25958 19496 25964 19508
rect 25919 19468 25964 19496
rect 25958 19456 25964 19468
rect 26016 19456 26022 19508
rect 14323 19400 14412 19428
rect 14323 19397 14335 19400
rect 14277 19391 14335 19397
rect 14734 19388 14740 19440
rect 14792 19428 14798 19440
rect 17497 19431 17555 19437
rect 14792 19400 15332 19428
rect 14792 19388 14798 19400
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 11808 19332 12449 19360
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 15197 19363 15255 19369
rect 15197 19360 15209 19363
rect 14884 19332 15209 19360
rect 14884 19320 14890 19332
rect 15197 19329 15209 19332
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 10226 19292 10232 19304
rect 10187 19264 10232 19292
rect 10226 19252 10232 19264
rect 10284 19252 10290 19304
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 14332 19264 14473 19292
rect 14332 19252 14338 19264
rect 14461 19261 14473 19264
rect 14507 19292 14519 19295
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14507 19264 15117 19292
rect 14507 19261 14519 19264
rect 14461 19255 14519 19261
rect 15105 19261 15117 19264
rect 15151 19261 15163 19295
rect 15105 19255 15163 19261
rect 12618 19184 12624 19236
rect 12676 19233 12682 19236
rect 12676 19227 12740 19233
rect 12676 19193 12694 19227
rect 12728 19193 12740 19227
rect 12676 19187 12740 19193
rect 12676 19184 12682 19187
rect 13906 19184 13912 19236
rect 13964 19224 13970 19236
rect 15013 19227 15071 19233
rect 15013 19224 15025 19227
rect 13964 19196 15025 19224
rect 13964 19184 13970 19196
rect 15013 19193 15025 19196
rect 15059 19193 15071 19227
rect 15013 19187 15071 19193
rect 11330 19156 11336 19168
rect 11291 19128 11336 19156
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 13814 19156 13820 19168
rect 13775 19128 13820 19156
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14274 19156 14280 19168
rect 14235 19128 14280 19156
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 14642 19156 14648 19168
rect 14603 19128 14648 19156
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 15304 19156 15332 19400
rect 17497 19397 17509 19431
rect 17543 19428 17555 19431
rect 18874 19428 18880 19440
rect 17543 19400 18880 19428
rect 17543 19397 17555 19400
rect 17497 19391 17555 19397
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16540 19332 17049 19360
rect 16540 19320 16546 19332
rect 17037 19329 17049 19332
rect 17083 19360 17095 19363
rect 17512 19360 17540 19391
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 23661 19431 23719 19437
rect 23661 19397 23673 19431
rect 23707 19397 23719 19431
rect 23661 19391 23719 19397
rect 17083 19332 17540 19360
rect 17083 19329 17095 19332
rect 17037 19323 17095 19329
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 17828 19332 17908 19360
rect 17828 19320 17834 19332
rect 15933 19295 15991 19301
rect 15933 19261 15945 19295
rect 15979 19292 15991 19295
rect 16761 19295 16819 19301
rect 16761 19292 16773 19295
rect 15979 19264 16773 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 16761 19261 16773 19264
rect 16807 19292 16819 19295
rect 16850 19292 16856 19304
rect 16807 19264 16856 19292
rect 16807 19261 16819 19264
rect 16761 19255 16819 19261
rect 16850 19252 16856 19264
rect 16908 19292 16914 19304
rect 17402 19292 17408 19304
rect 16908 19264 17408 19292
rect 16908 19252 16914 19264
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 17880 19292 17908 19332
rect 18138 19320 18144 19372
rect 18196 19320 18202 19372
rect 19150 19360 19156 19372
rect 19111 19332 19156 19360
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 22554 19360 22560 19372
rect 22515 19332 22560 19360
rect 22554 19320 22560 19332
rect 22612 19320 22618 19372
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 22830 19360 22836 19372
rect 22704 19332 22836 19360
rect 22704 19320 22710 19332
rect 22830 19320 22836 19332
rect 22888 19320 22894 19372
rect 23676 19360 23704 19391
rect 23400 19332 23704 19360
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17880 19264 18061 19292
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 15654 19184 15660 19236
rect 15712 19224 15718 19236
rect 17218 19224 17224 19236
rect 15712 19196 17224 19224
rect 15712 19184 15718 19196
rect 17218 19184 17224 19196
rect 17276 19224 17282 19236
rect 17773 19227 17831 19233
rect 17773 19224 17785 19227
rect 17276 19196 17785 19224
rect 17276 19184 17282 19196
rect 17773 19193 17785 19196
rect 17819 19224 17831 19227
rect 18156 19224 18184 19320
rect 19702 19292 19708 19304
rect 17819 19196 18184 19224
rect 18984 19264 19708 19292
rect 17819 19193 17831 19196
rect 17773 19187 17831 19193
rect 16206 19156 16212 19168
rect 15304 19128 16212 19156
rect 16206 19116 16212 19128
rect 16264 19116 16270 19168
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 16393 19159 16451 19165
rect 16393 19156 16405 19159
rect 16356 19128 16405 19156
rect 16356 19116 16362 19128
rect 16393 19125 16405 19128
rect 16439 19125 16451 19159
rect 16393 19119 16451 19125
rect 16482 19116 16488 19168
rect 16540 19156 16546 19168
rect 16853 19159 16911 19165
rect 16853 19156 16865 19159
rect 16540 19128 16865 19156
rect 16540 19116 16546 19128
rect 16853 19125 16865 19128
rect 16899 19156 16911 19159
rect 17310 19156 17316 19168
rect 16899 19128 17316 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 18984 19165 19012 19264
rect 19702 19252 19708 19264
rect 19760 19252 19766 19304
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19292 20959 19295
rect 22738 19292 22744 19304
rect 20947 19264 22744 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 19334 19184 19340 19236
rect 19392 19233 19398 19236
rect 19392 19227 19456 19233
rect 19392 19193 19410 19227
rect 19444 19193 19456 19227
rect 19392 19187 19456 19193
rect 19392 19184 19398 19187
rect 22094 19184 22100 19236
rect 22152 19224 22158 19236
rect 22373 19227 22431 19233
rect 22373 19224 22385 19227
rect 22152 19196 22385 19224
rect 22152 19184 22158 19196
rect 22373 19193 22385 19196
rect 22419 19224 22431 19227
rect 23400 19224 23428 19332
rect 24026 19320 24032 19372
rect 24084 19360 24090 19372
rect 24213 19363 24271 19369
rect 24213 19360 24225 19363
rect 24084 19332 24225 19360
rect 24084 19320 24090 19332
rect 24213 19329 24225 19332
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 23477 19295 23535 19301
rect 23477 19261 23489 19295
rect 23523 19292 23535 19295
rect 23658 19292 23664 19304
rect 23523 19264 23664 19292
rect 23523 19261 23535 19264
rect 23477 19255 23535 19261
rect 23658 19252 23664 19264
rect 23716 19292 23722 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 23716 19264 24133 19292
rect 23716 19252 23722 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 25222 19292 25228 19304
rect 25183 19264 25228 19292
rect 24121 19255 24179 19261
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 25498 19224 25504 19236
rect 22419 19196 23428 19224
rect 25459 19196 25504 19224
rect 22419 19193 22431 19196
rect 22373 19187 22431 19193
rect 25498 19184 25504 19196
rect 25556 19184 25562 19236
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18932 19128 18981 19156
rect 18932 19116 18938 19128
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 18969 19119 19027 19125
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 19116 19128 20545 19156
rect 19116 19116 19122 19128
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 20533 19119 20591 19125
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 22002 19156 22008 19168
rect 21963 19128 22008 19156
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 22465 19159 22523 19165
rect 22465 19125 22477 19159
rect 22511 19156 22523 19159
rect 22738 19156 22744 19168
rect 22511 19128 22744 19156
rect 22511 19125 22523 19128
rect 22465 19119 22523 19125
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 23109 19159 23167 19165
rect 23109 19125 23121 19159
rect 23155 19156 23167 19159
rect 24029 19159 24087 19165
rect 24029 19156 24041 19159
rect 23155 19128 24041 19156
rect 23155 19125 23167 19128
rect 23109 19119 23167 19125
rect 24029 19125 24041 19128
rect 24075 19156 24087 19159
rect 24118 19156 24124 19168
rect 24075 19128 24124 19156
rect 24075 19125 24087 19128
rect 24029 19119 24087 19125
rect 24118 19116 24124 19128
rect 24176 19116 24182 19168
rect 25133 19159 25191 19165
rect 25133 19125 25145 19159
rect 25179 19156 25191 19159
rect 25314 19156 25320 19168
rect 25179 19128 25320 19156
rect 25179 19125 25191 19128
rect 25133 19119 25191 19125
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 14369 18955 14427 18961
rect 14369 18952 14381 18955
rect 13688 18924 14381 18952
rect 13688 18912 13694 18924
rect 14369 18921 14381 18924
rect 14415 18921 14427 18955
rect 14369 18915 14427 18921
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 14553 18955 14611 18961
rect 14553 18952 14565 18955
rect 14516 18924 14565 18952
rect 14516 18912 14522 18924
rect 14553 18921 14565 18924
rect 14599 18921 14611 18955
rect 15654 18952 15660 18964
rect 15615 18924 15660 18952
rect 14553 18915 14611 18921
rect 15654 18912 15660 18924
rect 15712 18912 15718 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 17129 18955 17187 18961
rect 17129 18952 17141 18955
rect 16632 18924 17141 18952
rect 16632 18912 16638 18924
rect 17129 18921 17141 18924
rect 17175 18921 17187 18955
rect 17862 18952 17868 18964
rect 17823 18924 17868 18952
rect 17129 18915 17187 18921
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19392 18924 19809 18952
rect 19392 18912 19398 18924
rect 19797 18921 19809 18924
rect 19843 18952 19855 18955
rect 19978 18952 19984 18964
rect 19843 18924 19984 18952
rect 19843 18921 19855 18924
rect 19797 18915 19855 18921
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20714 18952 20720 18964
rect 20675 18924 20720 18952
rect 20714 18912 20720 18924
rect 20772 18912 20778 18964
rect 21361 18955 21419 18961
rect 21361 18921 21373 18955
rect 21407 18952 21419 18955
rect 21450 18952 21456 18964
rect 21407 18924 21456 18952
rect 21407 18921 21419 18924
rect 21361 18915 21419 18921
rect 21450 18912 21456 18924
rect 21508 18912 21514 18964
rect 22097 18955 22155 18961
rect 22097 18921 22109 18955
rect 22143 18952 22155 18955
rect 22554 18952 22560 18964
rect 22143 18924 22560 18952
rect 22143 18921 22155 18924
rect 22097 18915 22155 18921
rect 22554 18912 22560 18924
rect 22612 18952 22618 18964
rect 23198 18952 23204 18964
rect 22612 18924 23204 18952
rect 22612 18912 22618 18924
rect 23198 18912 23204 18924
rect 23256 18952 23262 18964
rect 23661 18955 23719 18961
rect 23661 18952 23673 18955
rect 23256 18924 23673 18952
rect 23256 18912 23262 18924
rect 23661 18921 23673 18924
rect 23707 18921 23719 18955
rect 23661 18915 23719 18921
rect 25222 18912 25228 18964
rect 25280 18952 25286 18964
rect 25501 18955 25559 18961
rect 25501 18952 25513 18955
rect 25280 18924 25513 18952
rect 25280 18912 25286 18924
rect 25501 18921 25513 18924
rect 25547 18921 25559 18955
rect 25501 18915 25559 18921
rect 13449 18887 13507 18893
rect 13449 18853 13461 18887
rect 13495 18884 13507 18887
rect 13998 18884 14004 18896
rect 13495 18856 14004 18884
rect 13495 18853 13507 18856
rect 13449 18847 13507 18853
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 19150 18884 19156 18896
rect 18432 18856 19156 18884
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11756 18788 11805 18816
rect 11756 18776 11762 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11793 18779 11851 18785
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13357 18819 13415 18825
rect 13357 18816 13369 18819
rect 12768 18788 13369 18816
rect 12768 18776 12774 18788
rect 13357 18785 13369 18788
rect 13403 18785 13415 18819
rect 14734 18816 14740 18828
rect 14695 18788 14740 18816
rect 13357 18779 13415 18785
rect 14734 18776 14740 18788
rect 14792 18776 14798 18828
rect 16390 18776 16396 18828
rect 16448 18816 16454 18828
rect 18432 18825 18460 18856
rect 19150 18844 19156 18856
rect 19208 18844 19214 18896
rect 24857 18887 24915 18893
rect 24857 18853 24869 18887
rect 24903 18884 24915 18887
rect 25038 18884 25044 18896
rect 24903 18856 25044 18884
rect 24903 18853 24915 18856
rect 24857 18847 24915 18853
rect 25038 18844 25044 18856
rect 25096 18844 25102 18896
rect 16485 18819 16543 18825
rect 16485 18816 16497 18819
rect 16448 18788 16497 18816
rect 16448 18776 16454 18788
rect 16485 18785 16497 18788
rect 16531 18785 16543 18819
rect 16485 18779 16543 18785
rect 18417 18819 18475 18825
rect 18417 18785 18429 18819
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 18506 18776 18512 18828
rect 18564 18816 18570 18828
rect 18673 18819 18731 18825
rect 18673 18816 18685 18819
rect 18564 18788 18685 18816
rect 18564 18776 18570 18788
rect 18673 18785 18685 18788
rect 18719 18785 18731 18819
rect 21174 18816 21180 18828
rect 21135 18788 21180 18816
rect 18673 18779 18731 18785
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 22370 18776 22376 18828
rect 22428 18816 22434 18828
rect 22537 18819 22595 18825
rect 22537 18816 22549 18819
rect 22428 18788 22549 18816
rect 22428 18776 22434 18788
rect 22537 18785 22549 18788
rect 22583 18816 22595 18819
rect 23937 18819 23995 18825
rect 23937 18816 23949 18819
rect 22583 18788 23949 18816
rect 22583 18785 22595 18788
rect 22537 18779 22595 18785
rect 23937 18785 23949 18788
rect 23983 18816 23995 18819
rect 24026 18816 24032 18828
rect 23983 18788 24032 18816
rect 23983 18785 23995 18788
rect 23937 18779 23995 18785
rect 24026 18776 24032 18788
rect 24084 18816 24090 18828
rect 24305 18819 24363 18825
rect 24305 18816 24317 18819
rect 24084 18788 24317 18816
rect 24084 18776 24090 18788
rect 24305 18785 24317 18788
rect 24351 18785 24363 18819
rect 24305 18779 24363 18785
rect 11514 18708 11520 18760
rect 11572 18748 11578 18760
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11572 18720 11897 18748
rect 11572 18708 11578 18720
rect 11885 18717 11897 18720
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12250 18748 12256 18760
rect 12115 18720 12256 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18748 13691 18751
rect 14182 18748 14188 18760
rect 13679 18720 14188 18748
rect 13679 18717 13691 18720
rect 13633 18711 13691 18717
rect 11422 18680 11428 18692
rect 11383 18652 11428 18680
rect 11422 18640 11428 18652
rect 11480 18640 11486 18692
rect 12529 18683 12587 18689
rect 12529 18649 12541 18683
rect 12575 18680 12587 18683
rect 12618 18680 12624 18692
rect 12575 18652 12624 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 12618 18640 12624 18652
rect 12676 18680 12682 18692
rect 13648 18680 13676 18711
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 16577 18751 16635 18757
rect 16577 18748 16589 18751
rect 16264 18720 16589 18748
rect 16264 18708 16270 18720
rect 16577 18717 16589 18720
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 16669 18751 16727 18757
rect 16669 18717 16681 18751
rect 16715 18717 16727 18751
rect 22278 18748 22284 18760
rect 22239 18720 22284 18748
rect 16669 18711 16727 18717
rect 12676 18652 13676 18680
rect 12676 18640 12682 18652
rect 16482 18640 16488 18692
rect 16540 18680 16546 18692
rect 16684 18680 16712 18711
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 24946 18748 24952 18760
rect 24907 18720 24952 18748
rect 24946 18708 24952 18720
rect 25004 18708 25010 18760
rect 25130 18748 25136 18760
rect 25091 18720 25136 18748
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 16540 18652 16712 18680
rect 16540 18640 16546 18652
rect 24210 18640 24216 18692
rect 24268 18680 24274 18692
rect 24489 18683 24547 18689
rect 24489 18680 24501 18683
rect 24268 18652 24501 18680
rect 24268 18640 24274 18652
rect 24489 18649 24501 18652
rect 24535 18649 24547 18683
rect 24489 18643 24547 18649
rect 12894 18612 12900 18624
rect 12855 18584 12900 18612
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 12989 18615 13047 18621
rect 12989 18581 13001 18615
rect 13035 18612 13047 18615
rect 13170 18612 13176 18624
rect 13035 18584 13176 18612
rect 13035 18581 13047 18584
rect 12989 18575 13047 18581
rect 13170 18572 13176 18584
rect 13228 18612 13234 18624
rect 14001 18615 14059 18621
rect 14001 18612 14013 18615
rect 13228 18584 14013 18612
rect 13228 18572 13234 18584
rect 14001 18581 14013 18584
rect 14047 18581 14059 18615
rect 14001 18575 14059 18581
rect 15105 18615 15163 18621
rect 15105 18581 15117 18615
rect 15151 18612 15163 18615
rect 15562 18612 15568 18624
rect 15151 18584 15568 18612
rect 15151 18581 15163 18584
rect 15105 18575 15163 18581
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 15933 18615 15991 18621
rect 15933 18612 15945 18615
rect 15712 18584 15945 18612
rect 15712 18572 15718 18584
rect 15933 18581 15945 18584
rect 15979 18581 15991 18615
rect 16114 18612 16120 18624
rect 16075 18584 16120 18612
rect 15933 18575 15991 18581
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 18141 18615 18199 18621
rect 18141 18612 18153 18615
rect 18012 18584 18153 18612
rect 18012 18572 18018 18584
rect 18141 18581 18153 18584
rect 18187 18581 18199 18615
rect 20070 18612 20076 18624
rect 20031 18584 20076 18612
rect 18141 18575 18199 18581
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 11330 18368 11336 18420
rect 11388 18408 11394 18420
rect 12710 18408 12716 18420
rect 11388 18380 12716 18408
rect 11388 18368 11394 18380
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 13909 18411 13967 18417
rect 13909 18377 13921 18411
rect 13955 18408 13967 18411
rect 13998 18408 14004 18420
rect 13955 18380 14004 18408
rect 13955 18377 13967 18380
rect 13909 18371 13967 18377
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 14182 18408 14188 18420
rect 14143 18380 14188 18408
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 14550 18368 14556 18420
rect 14608 18408 14614 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 14608 18380 14841 18408
rect 14608 18368 14614 18380
rect 14829 18377 14841 18380
rect 14875 18408 14887 18411
rect 19058 18408 19064 18420
rect 14875 18380 15516 18408
rect 19019 18380 19064 18408
rect 14875 18377 14887 18380
rect 14829 18371 14887 18377
rect 11514 18300 11520 18352
rect 11572 18340 11578 18352
rect 11698 18340 11704 18352
rect 11572 18312 11704 18340
rect 11572 18300 11578 18312
rect 11698 18300 11704 18312
rect 11756 18340 11762 18352
rect 11793 18343 11851 18349
rect 11793 18340 11805 18343
rect 11756 18312 11805 18340
rect 11756 18300 11762 18312
rect 11793 18309 11805 18312
rect 11839 18309 11851 18343
rect 11793 18303 11851 18309
rect 12434 18300 12440 18352
rect 12492 18340 12498 18352
rect 12805 18343 12863 18349
rect 12805 18340 12817 18343
rect 12492 18312 12817 18340
rect 12492 18300 12498 18312
rect 12805 18309 12817 18312
rect 12851 18309 12863 18343
rect 14016 18340 14044 18368
rect 14274 18340 14280 18352
rect 14016 18312 14280 18340
rect 12805 18303 12863 18309
rect 14274 18300 14280 18312
rect 14332 18300 14338 18352
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 13265 18275 13323 18281
rect 13265 18272 13277 18275
rect 12952 18244 13277 18272
rect 12952 18232 12958 18244
rect 13265 18241 13277 18244
rect 13311 18241 13323 18275
rect 13446 18272 13452 18284
rect 13359 18244 13452 18272
rect 13265 18235 13323 18241
rect 13446 18232 13452 18244
rect 13504 18272 13510 18284
rect 13814 18272 13820 18284
rect 13504 18244 13820 18272
rect 13504 18232 13510 18244
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 15488 18281 15516 18380
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20625 18411 20683 18417
rect 20625 18408 20637 18411
rect 20036 18380 20637 18408
rect 20036 18368 20042 18380
rect 20625 18377 20637 18380
rect 20671 18408 20683 18411
rect 22370 18408 22376 18420
rect 20671 18380 20944 18408
rect 22331 18380 22376 18408
rect 20671 18377 20683 18380
rect 20625 18371 20683 18377
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15562 18232 15568 18284
rect 15620 18272 15626 18284
rect 15620 18244 15665 18272
rect 15620 18232 15626 18244
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 17313 18275 17371 18281
rect 17313 18272 17325 18275
rect 16448 18244 17325 18272
rect 16448 18232 16454 18244
rect 17313 18241 17325 18244
rect 17359 18241 17371 18275
rect 19076 18272 19104 18368
rect 19245 18343 19303 18349
rect 19245 18309 19257 18343
rect 19291 18340 19303 18343
rect 19426 18340 19432 18352
rect 19291 18312 19432 18340
rect 19291 18309 19303 18312
rect 19245 18303 19303 18309
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 20070 18300 20076 18352
rect 20128 18340 20134 18352
rect 20809 18343 20867 18349
rect 20809 18340 20821 18343
rect 20128 18312 20821 18340
rect 20128 18300 20134 18312
rect 20809 18309 20821 18312
rect 20855 18309 20867 18343
rect 20809 18303 20867 18309
rect 19797 18275 19855 18281
rect 19797 18272 19809 18275
rect 19076 18244 19809 18272
rect 17313 18235 17371 18241
rect 19797 18241 19809 18244
rect 19843 18241 19855 18275
rect 20254 18272 20260 18284
rect 20215 18244 20260 18272
rect 19797 18235 19855 18241
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 20916 18272 20944 18380
rect 22370 18368 22376 18380
rect 22428 18368 22434 18420
rect 22646 18408 22652 18420
rect 22607 18380 22652 18408
rect 22646 18368 22652 18380
rect 22704 18368 22710 18420
rect 22738 18368 22744 18420
rect 22796 18408 22802 18420
rect 23661 18411 23719 18417
rect 23661 18408 23673 18411
rect 22796 18380 23673 18408
rect 22796 18368 22802 18380
rect 23661 18377 23673 18380
rect 23707 18377 23719 18411
rect 23661 18371 23719 18377
rect 24118 18368 24124 18420
rect 24176 18408 24182 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 24176 18380 24685 18408
rect 24176 18368 24182 18380
rect 24673 18377 24685 18380
rect 24719 18408 24731 18411
rect 24946 18408 24952 18420
rect 24719 18380 24952 18408
rect 24719 18377 24731 18380
rect 24673 18371 24731 18377
rect 24946 18368 24952 18380
rect 25004 18368 25010 18420
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 20916 18244 21373 18272
rect 21361 18241 21373 18244
rect 21407 18241 21419 18275
rect 21818 18272 21824 18284
rect 21779 18244 21824 18272
rect 21361 18235 21419 18241
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 24026 18232 24032 18284
rect 24084 18272 24090 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 24084 18244 24225 18272
rect 24084 18232 24090 18244
rect 24213 18241 24225 18244
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 11422 18204 11428 18216
rect 11383 18176 11428 18204
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 13170 18204 13176 18216
rect 13131 18176 13176 18204
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 16574 18204 16580 18216
rect 16535 18176 16580 18204
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 20070 18204 20076 18216
rect 19751 18176 20076 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 15194 18096 15200 18148
rect 15252 18136 15258 18148
rect 15381 18139 15439 18145
rect 15381 18136 15393 18139
rect 15252 18108 15393 18136
rect 15252 18096 15258 18108
rect 15381 18105 15393 18108
rect 15427 18136 15439 18139
rect 15838 18136 15844 18148
rect 15427 18108 15844 18136
rect 15427 18105 15439 18108
rect 15381 18099 15439 18105
rect 15838 18096 15844 18108
rect 15896 18096 15902 18148
rect 16850 18136 16856 18148
rect 16811 18108 16856 18136
rect 16850 18096 16856 18108
rect 16908 18096 16914 18148
rect 17954 18096 17960 18148
rect 18012 18136 18018 18148
rect 18506 18136 18512 18148
rect 18012 18108 18512 18136
rect 18012 18096 18018 18108
rect 18506 18096 18512 18108
rect 18564 18136 18570 18148
rect 18693 18139 18751 18145
rect 18693 18136 18705 18139
rect 18564 18108 18705 18136
rect 18564 18096 18570 18108
rect 18693 18105 18705 18108
rect 18739 18105 18751 18139
rect 20272 18136 20300 18232
rect 20714 18164 20720 18216
rect 20772 18204 20778 18216
rect 21177 18207 21235 18213
rect 21177 18204 21189 18207
rect 20772 18176 21189 18204
rect 20772 18164 20778 18176
rect 21177 18173 21189 18176
rect 21223 18173 21235 18207
rect 22462 18204 22468 18216
rect 22423 18176 22468 18204
rect 21177 18167 21235 18173
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 22738 18164 22744 18216
rect 22796 18204 22802 18216
rect 23014 18204 23020 18216
rect 22796 18176 23020 18204
rect 22796 18164 22802 18176
rect 23014 18164 23020 18176
rect 23072 18204 23078 18216
rect 25222 18204 25228 18216
rect 23072 18176 24072 18204
rect 25183 18176 25228 18204
rect 23072 18164 23078 18176
rect 24044 18145 24072 18176
rect 25222 18164 25228 18176
rect 25280 18204 25286 18216
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25280 18176 25789 18204
rect 25280 18164 25286 18176
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 21269 18139 21327 18145
rect 21269 18136 21281 18139
rect 20272 18108 21281 18136
rect 18693 18099 18751 18105
rect 21269 18105 21281 18108
rect 21315 18105 21327 18139
rect 21269 18099 21327 18105
rect 24029 18139 24087 18145
rect 24029 18105 24041 18139
rect 24075 18105 24087 18139
rect 24029 18099 24087 18105
rect 12250 18068 12256 18080
rect 12211 18040 12256 18068
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 15013 18071 15071 18077
rect 15013 18037 15025 18071
rect 15059 18068 15071 18071
rect 15102 18068 15108 18080
rect 15059 18040 15108 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 16209 18071 16267 18077
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 16482 18068 16488 18080
rect 16255 18040 16488 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 18046 18068 18052 18080
rect 17911 18040 18052 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18230 18068 18236 18080
rect 18191 18040 18236 18068
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19392 18040 19625 18068
rect 19392 18028 19398 18040
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 19613 18031 19671 18037
rect 23014 18028 23020 18080
rect 23072 18068 23078 18080
rect 23385 18071 23443 18077
rect 23385 18068 23397 18071
rect 23072 18040 23397 18068
rect 23072 18028 23078 18040
rect 23385 18037 23397 18040
rect 23431 18068 23443 18071
rect 24121 18071 24179 18077
rect 24121 18068 24133 18071
rect 23431 18040 24133 18068
rect 23431 18037 23443 18040
rect 23385 18031 23443 18037
rect 24121 18037 24133 18040
rect 24167 18037 24179 18071
rect 25038 18068 25044 18080
rect 24999 18040 25044 18068
rect 24121 18031 24179 18037
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 25406 18068 25412 18080
rect 25367 18040 25412 18068
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12952 17836 13001 17864
rect 12952 17824 12958 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 14093 17867 14151 17873
rect 14093 17864 14105 17867
rect 13495 17836 14105 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 14093 17833 14105 17836
rect 14139 17864 14151 17867
rect 14642 17864 14648 17876
rect 14139 17836 14648 17864
rect 14139 17833 14151 17836
rect 14093 17827 14151 17833
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 15010 17864 15016 17876
rect 14971 17836 15016 17864
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 16206 17864 16212 17876
rect 16167 17836 16212 17864
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 17954 17864 17960 17876
rect 17915 17836 17960 17864
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 18877 17867 18935 17873
rect 18877 17833 18889 17867
rect 18923 17864 18935 17867
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 18923 17836 19625 17864
rect 18923 17833 18935 17836
rect 18877 17827 18935 17833
rect 19613 17833 19625 17836
rect 19659 17864 19671 17867
rect 20901 17867 20959 17873
rect 20901 17864 20913 17867
rect 19659 17836 20913 17864
rect 19659 17833 19671 17836
rect 19613 17827 19671 17833
rect 20901 17833 20913 17836
rect 20947 17833 20959 17867
rect 20901 17827 20959 17833
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22152 17836 22197 17864
rect 22152 17824 22158 17836
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24305 17867 24363 17873
rect 24305 17864 24317 17867
rect 24084 17836 24317 17864
rect 24084 17824 24090 17836
rect 24305 17833 24317 17836
rect 24351 17864 24363 17867
rect 24673 17867 24731 17873
rect 24673 17864 24685 17867
rect 24351 17836 24685 17864
rect 24351 17833 24363 17836
rect 24305 17827 24363 17833
rect 24673 17833 24685 17836
rect 24719 17864 24731 17867
rect 25130 17864 25136 17876
rect 24719 17836 25136 17864
rect 24719 17833 24731 17836
rect 24673 17827 24731 17833
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 14553 17799 14611 17805
rect 14553 17765 14565 17799
rect 14599 17796 14611 17799
rect 14734 17796 14740 17808
rect 14599 17768 14740 17796
rect 14599 17765 14611 17768
rect 14553 17759 14611 17765
rect 14734 17756 14740 17768
rect 14792 17756 14798 17808
rect 16574 17756 16580 17808
rect 16632 17796 16638 17808
rect 16844 17799 16902 17805
rect 16844 17796 16856 17799
rect 16632 17768 16856 17796
rect 16632 17756 16638 17768
rect 16844 17765 16856 17768
rect 16890 17796 16902 17799
rect 16942 17796 16948 17808
rect 16890 17768 16948 17796
rect 16890 17765 16902 17768
rect 16844 17759 16902 17765
rect 16942 17756 16948 17768
rect 17000 17756 17006 17808
rect 18506 17756 18512 17808
rect 18564 17796 18570 17808
rect 18564 17768 19288 17796
rect 18564 17756 18570 17768
rect 11698 17728 11704 17740
rect 11659 17700 11704 17728
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 12342 17728 12348 17740
rect 11756 17700 12348 17728
rect 11756 17688 11762 17700
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17728 13415 17731
rect 13538 17728 13544 17740
rect 13403 17700 13544 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 14366 17688 14372 17740
rect 14424 17728 14430 17740
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 14424 17700 15301 17728
rect 14424 17688 14430 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 17770 17728 17776 17740
rect 15289 17691 15347 17697
rect 16592 17700 17776 17728
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12897 17663 12955 17669
rect 12897 17629 12909 17663
rect 12943 17660 12955 17663
rect 13446 17660 13452 17672
rect 12943 17632 13452 17660
rect 12943 17629 12955 17632
rect 12897 17623 12955 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 13633 17663 13691 17669
rect 13633 17629 13645 17663
rect 13679 17660 13691 17663
rect 14182 17660 14188 17672
rect 13679 17632 14188 17660
rect 13679 17629 13691 17632
rect 13633 17623 13691 17629
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 15565 17663 15623 17669
rect 15565 17629 15577 17663
rect 15611 17660 15623 17663
rect 15930 17660 15936 17672
rect 15611 17632 15936 17660
rect 15611 17629 15623 17632
rect 15565 17623 15623 17629
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 16592 17669 16620 17700
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18322 17728 18328 17740
rect 18012 17700 18328 17728
rect 18012 17688 18018 17700
rect 18322 17688 18328 17700
rect 18380 17728 18386 17740
rect 19153 17731 19211 17737
rect 19153 17728 19165 17731
rect 18380 17700 19165 17728
rect 18380 17688 18386 17700
rect 19153 17697 19165 17700
rect 19199 17697 19211 17731
rect 19260 17728 19288 17768
rect 19334 17756 19340 17808
rect 19392 17796 19398 17808
rect 19705 17799 19763 17805
rect 19705 17796 19717 17799
rect 19392 17768 19717 17796
rect 19392 17756 19398 17768
rect 19705 17765 19717 17768
rect 19751 17796 19763 17799
rect 20162 17796 20168 17808
rect 19751 17768 20168 17796
rect 19751 17765 19763 17768
rect 19705 17759 19763 17765
rect 20162 17756 20168 17768
rect 20220 17756 20226 17808
rect 23198 17805 23204 17808
rect 23192 17796 23204 17805
rect 23159 17768 23204 17796
rect 23192 17759 23204 17768
rect 23198 17756 23204 17759
rect 23256 17756 23262 17808
rect 20717 17731 20775 17737
rect 20717 17728 20729 17731
rect 19260 17700 20729 17728
rect 19153 17691 19211 17697
rect 20717 17697 20729 17700
rect 20763 17697 20775 17731
rect 21266 17728 21272 17740
rect 21227 17700 21272 17728
rect 20717 17691 20775 17697
rect 16577 17663 16635 17669
rect 16577 17629 16589 17663
rect 16623 17629 16635 17663
rect 19168 17660 19196 17691
rect 19889 17663 19947 17669
rect 19168 17632 19380 17660
rect 16577 17623 16635 17629
rect 12529 17595 12587 17601
rect 12529 17561 12541 17595
rect 12575 17592 12587 17595
rect 12618 17592 12624 17604
rect 12575 17564 12624 17592
rect 12575 17561 12587 17564
rect 12529 17555 12587 17561
rect 12618 17552 12624 17564
rect 12676 17552 12682 17604
rect 18046 17552 18052 17604
rect 18104 17592 18110 17604
rect 19242 17592 19248 17604
rect 18104 17564 19248 17592
rect 18104 17552 18110 17564
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 19352 17592 19380 17632
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 19978 17660 19984 17672
rect 19935 17632 19984 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20257 17595 20315 17601
rect 20257 17592 20269 17595
rect 19352 17564 20269 17592
rect 20257 17561 20269 17564
rect 20303 17561 20315 17595
rect 20732 17592 20760 17691
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17728 25191 17731
rect 25222 17728 25228 17740
rect 25179 17700 25228 17728
rect 25179 17697 25191 17700
rect 25133 17691 25191 17697
rect 25222 17688 25228 17700
rect 25280 17688 25286 17740
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20956 17632 21373 17660
rect 20956 17620 20962 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 21453 17663 21511 17669
rect 21453 17629 21465 17663
rect 21499 17660 21511 17663
rect 21542 17660 21548 17672
rect 21499 17632 21548 17660
rect 21499 17629 21511 17632
rect 21453 17623 21511 17629
rect 21468 17592 21496 17623
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 22922 17660 22928 17672
rect 22883 17632 22928 17660
rect 22922 17620 22928 17632
rect 22980 17620 22986 17672
rect 20732 17564 21496 17592
rect 20257 17555 20315 17561
rect 11609 17527 11667 17533
rect 11609 17493 11621 17527
rect 11655 17524 11667 17527
rect 11882 17524 11888 17536
rect 11655 17496 11888 17524
rect 11655 17493 11667 17496
rect 11609 17487 11667 17493
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 18230 17524 18236 17536
rect 18191 17496 18236 17524
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18966 17524 18972 17536
rect 18927 17496 18972 17524
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 22462 17524 22468 17536
rect 22423 17496 22468 17524
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 25314 17524 25320 17536
rect 25275 17496 25320 17524
rect 25314 17484 25320 17496
rect 25372 17484 25378 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 10965 17323 11023 17329
rect 10965 17289 10977 17323
rect 11011 17320 11023 17323
rect 11698 17320 11704 17332
rect 11011 17292 11704 17320
rect 11011 17289 11023 17292
rect 10965 17283 11023 17289
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 14182 17320 14188 17332
rect 14143 17292 14188 17320
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 19337 17323 19395 17329
rect 19337 17289 19349 17323
rect 19383 17320 19395 17323
rect 19978 17320 19984 17332
rect 19383 17292 19984 17320
rect 19383 17289 19395 17292
rect 19337 17283 19395 17289
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 22373 17323 22431 17329
rect 22373 17320 22385 17323
rect 21324 17292 22385 17320
rect 21324 17280 21330 17292
rect 22373 17289 22385 17292
rect 22419 17289 22431 17323
rect 22373 17283 22431 17289
rect 23109 17323 23167 17329
rect 23109 17289 23121 17323
rect 23155 17320 23167 17323
rect 23198 17320 23204 17332
rect 23155 17292 23204 17320
rect 23155 17289 23167 17292
rect 23109 17283 23167 17289
rect 23198 17280 23204 17292
rect 23256 17280 23262 17332
rect 14642 17252 14648 17264
rect 13464 17224 14648 17252
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 11606 17184 11612 17196
rect 11379 17156 11612 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 11057 17119 11115 17125
rect 11057 17085 11069 17119
rect 11103 17116 11115 17119
rect 11103 17088 11928 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11900 17057 11928 17088
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12032 17088 12449 17116
rect 12032 17076 12038 17088
rect 12437 17085 12449 17088
rect 12483 17116 12495 17119
rect 13464 17116 13492 17224
rect 14642 17212 14648 17224
rect 14700 17252 14706 17264
rect 14700 17224 15608 17252
rect 14700 17212 14706 17224
rect 12483 17088 13492 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 14826 17116 14832 17128
rect 14516 17088 14832 17116
rect 14516 17076 14522 17088
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 15580 17125 15608 17224
rect 21910 17212 21916 17264
rect 21968 17252 21974 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21968 17224 22017 17252
rect 21968 17212 21974 17224
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 25314 17252 25320 17264
rect 25275 17224 25320 17252
rect 22005 17215 22063 17221
rect 25314 17212 25320 17224
rect 25372 17212 25378 17264
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 18288 17156 18613 17184
rect 18288 17144 18294 17156
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 19978 17184 19984 17196
rect 19939 17156 19984 17184
rect 18601 17147 18659 17153
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 20772 17156 21557 17184
rect 20772 17144 20778 17156
rect 21545 17153 21557 17156
rect 21591 17153 21603 17187
rect 21545 17147 21603 17153
rect 15565 17119 15623 17125
rect 15565 17085 15577 17119
rect 15611 17116 15623 17119
rect 15654 17116 15660 17128
rect 15611 17088 15660 17116
rect 15611 17085 15623 17088
rect 15565 17079 15623 17085
rect 15654 17076 15660 17088
rect 15712 17076 15718 17128
rect 17310 17076 17316 17128
rect 17368 17116 17374 17128
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17368 17088 17877 17116
rect 17368 17076 17374 17088
rect 17865 17085 17877 17088
rect 17911 17116 17923 17119
rect 17911 17088 18552 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 12342 17048 12348 17060
rect 11931 17020 12348 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 12342 17008 12348 17020
rect 12400 17008 12406 17060
rect 12704 17051 12762 17057
rect 12704 17017 12716 17051
rect 12750 17048 12762 17051
rect 12802 17048 12808 17060
rect 12750 17020 12808 17048
rect 12750 17017 12762 17020
rect 12704 17011 12762 17017
rect 12802 17008 12808 17020
rect 12860 17008 12866 17060
rect 13170 17008 13176 17060
rect 13228 17048 13234 17060
rect 14366 17048 14372 17060
rect 13228 17020 14372 17048
rect 13228 17008 13234 17020
rect 14366 17008 14372 17020
rect 14424 17048 14430 17060
rect 14553 17051 14611 17057
rect 14553 17048 14565 17051
rect 14424 17020 14565 17048
rect 14424 17008 14430 17020
rect 14553 17017 14565 17020
rect 14599 17017 14611 17051
rect 14553 17011 14611 17017
rect 15473 17051 15531 17057
rect 15473 17017 15485 17051
rect 15519 17048 15531 17051
rect 15810 17051 15868 17057
rect 15810 17048 15822 17051
rect 15519 17020 15822 17048
rect 15519 17017 15531 17020
rect 15473 17011 15531 17017
rect 15810 17017 15822 17020
rect 15856 17048 15868 17051
rect 16574 17048 16580 17060
rect 15856 17020 16580 17048
rect 15856 17017 15868 17020
rect 15810 17011 15868 17017
rect 16574 17008 16580 17020
rect 16632 17008 16638 17060
rect 18417 17051 18475 17057
rect 18417 17048 18429 17051
rect 17420 17020 18429 17048
rect 17420 16992 17448 17020
rect 18417 17017 18429 17020
rect 18463 17017 18475 17051
rect 18417 17011 18475 17017
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11296 16952 12173 16980
rect 11296 16940 11302 16952
rect 12161 16949 12173 16952
rect 12207 16980 12219 16983
rect 13446 16980 13452 16992
rect 12207 16952 13452 16980
rect 12207 16949 12219 16952
rect 12161 16943 12219 16949
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 13596 16952 13829 16980
rect 13596 16940 13602 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 13817 16943 13875 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17402 16980 17408 16992
rect 17363 16952 17408 16980
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18524 16989 18552 17088
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19484 17088 19717 17116
rect 19484 17076 19490 17088
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 21361 17119 21419 17125
rect 20671 17088 21312 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 18690 17008 18696 17060
rect 18748 17048 18754 17060
rect 20809 17051 20867 17057
rect 20809 17048 20821 17051
rect 18748 17020 20821 17048
rect 18748 17008 18754 17020
rect 20809 17017 20821 17020
rect 20855 17048 20867 17051
rect 20898 17048 20904 17060
rect 20855 17020 20904 17048
rect 20855 17017 20867 17020
rect 20809 17011 20867 17017
rect 20898 17008 20904 17020
rect 20956 17008 20962 17060
rect 21284 17048 21312 17088
rect 21361 17085 21373 17119
rect 21407 17116 21419 17119
rect 21928 17116 21956 17212
rect 22554 17184 22560 17196
rect 22515 17156 22560 17184
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 22094 17116 22100 17128
rect 21407 17088 22100 17116
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 22094 17076 22100 17088
rect 22152 17076 22158 17128
rect 22186 17076 22192 17128
rect 22244 17116 22250 17128
rect 22922 17116 22928 17128
rect 22244 17088 22928 17116
rect 22244 17076 22250 17088
rect 22922 17076 22928 17088
rect 22980 17116 22986 17128
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 22980 17088 23673 17116
rect 22980 17076 22986 17088
rect 23661 17085 23673 17088
rect 23707 17116 23719 17119
rect 23707 17088 24164 17116
rect 23707 17085 23719 17088
rect 23661 17079 23719 17085
rect 24136 17060 24164 17088
rect 21450 17048 21456 17060
rect 21284 17020 21456 17048
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 23477 17051 23535 17057
rect 23477 17017 23489 17051
rect 23523 17048 23535 17051
rect 23928 17051 23986 17057
rect 23928 17048 23940 17051
rect 23523 17020 23940 17048
rect 23523 17017 23535 17020
rect 23477 17011 23535 17017
rect 23928 17017 23940 17020
rect 23974 17048 23986 17051
rect 24026 17048 24032 17060
rect 23974 17020 24032 17048
rect 23974 17017 23986 17020
rect 23928 17011 23986 17017
rect 24026 17008 24032 17020
rect 24084 17008 24090 17060
rect 24118 17008 24124 17060
rect 24176 17008 24182 17060
rect 18049 16983 18107 16989
rect 18049 16980 18061 16983
rect 18012 16952 18061 16980
rect 18012 16940 18018 16952
rect 18049 16949 18061 16952
rect 18095 16949 18107 16983
rect 18049 16943 18107 16949
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16980 18567 16983
rect 18598 16980 18604 16992
rect 18555 16952 18604 16980
rect 18555 16949 18567 16952
rect 18509 16943 18567 16949
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 19300 16952 20453 16980
rect 19300 16940 19306 16952
rect 20441 16949 20453 16952
rect 20487 16980 20499 16983
rect 20625 16983 20683 16989
rect 20625 16980 20637 16983
rect 20487 16952 20637 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 20625 16949 20637 16952
rect 20671 16949 20683 16983
rect 20990 16980 20996 16992
rect 20951 16952 20996 16980
rect 20625 16943 20683 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 23290 16980 23296 16992
rect 22152 16952 23296 16980
rect 22152 16940 22158 16952
rect 23290 16940 23296 16952
rect 23348 16940 23354 16992
rect 25038 16980 25044 16992
rect 24999 16952 25044 16980
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 10870 16776 10876 16788
rect 10831 16748 10876 16776
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 14458 16776 14464 16788
rect 14419 16748 14464 16776
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 14826 16776 14832 16788
rect 14787 16748 14832 16776
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16632 16748 16681 16776
rect 16632 16736 16638 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16942 16776 16948 16788
rect 16903 16748 16948 16776
rect 16669 16739 16727 16745
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 17770 16736 17776 16788
rect 17828 16776 17834 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 17828 16748 17877 16776
rect 17828 16736 17834 16748
rect 17865 16745 17877 16748
rect 17911 16745 17923 16779
rect 17865 16739 17923 16745
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 18141 16779 18199 16785
rect 18141 16776 18153 16779
rect 18104 16748 18153 16776
rect 18104 16736 18110 16748
rect 18141 16745 18153 16748
rect 18187 16745 18199 16779
rect 18506 16776 18512 16788
rect 18419 16748 18512 16776
rect 18141 16739 18199 16745
rect 18506 16736 18512 16748
rect 18564 16776 18570 16788
rect 19334 16776 19340 16788
rect 18564 16748 19196 16776
rect 19295 16748 19340 16776
rect 18564 16736 18570 16748
rect 11977 16711 12035 16717
rect 11977 16677 11989 16711
rect 12023 16708 12035 16711
rect 12526 16708 12532 16720
rect 12023 16680 12532 16708
rect 12023 16677 12035 16680
rect 11977 16671 12035 16677
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 15562 16717 15568 16720
rect 15556 16708 15568 16717
rect 15523 16680 15568 16708
rect 15556 16671 15568 16680
rect 15562 16668 15568 16671
rect 15620 16668 15626 16720
rect 15654 16668 15660 16720
rect 15712 16668 15718 16720
rect 17405 16711 17463 16717
rect 17405 16677 17417 16711
rect 17451 16708 17463 16711
rect 18966 16708 18972 16720
rect 17451 16680 18972 16708
rect 17451 16677 17463 16680
rect 17405 16671 17463 16677
rect 11238 16640 11244 16652
rect 11199 16612 11244 16640
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16640 11391 16643
rect 11606 16640 11612 16652
rect 11379 16612 11612 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 12704 16643 12762 16649
rect 12704 16640 12716 16643
rect 12360 16612 12716 16640
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16572 11575 16575
rect 11698 16572 11704 16584
rect 11563 16544 11704 16572
rect 11563 16541 11575 16544
rect 11517 16535 11575 16541
rect 11698 16532 11704 16544
rect 11756 16572 11762 16584
rect 12360 16572 12388 16612
rect 12704 16609 12716 16612
rect 12750 16640 12762 16643
rect 13538 16640 13544 16652
rect 12750 16612 13544 16640
rect 12750 16609 12762 16612
rect 12704 16603 12762 16609
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15672 16640 15700 16668
rect 17678 16640 17684 16652
rect 15335 16612 15700 16640
rect 17639 16612 17684 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 17678 16600 17684 16612
rect 17736 16600 17742 16652
rect 18064 16649 18092 16680
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 19168 16708 19196 16748
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 20257 16779 20315 16785
rect 20257 16776 20269 16779
rect 19484 16748 20269 16776
rect 19484 16736 19490 16748
rect 20257 16745 20269 16748
rect 20303 16745 20315 16779
rect 20714 16776 20720 16788
rect 20675 16748 20720 16776
rect 20257 16739 20315 16745
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 22278 16776 22284 16788
rect 22239 16748 22284 16776
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 23934 16776 23940 16788
rect 23895 16748 23940 16776
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 24210 16736 24216 16788
rect 24268 16776 24274 16788
rect 24305 16779 24363 16785
rect 24305 16776 24317 16779
rect 24268 16748 24317 16776
rect 24268 16736 24274 16748
rect 24305 16745 24317 16748
rect 24351 16776 24363 16779
rect 24946 16776 24952 16788
rect 24351 16748 24952 16776
rect 24351 16745 24363 16748
rect 24305 16739 24363 16745
rect 24946 16736 24952 16748
rect 25004 16736 25010 16788
rect 21726 16708 21732 16720
rect 19168 16680 21732 16708
rect 21726 16668 21732 16680
rect 21784 16668 21790 16720
rect 23845 16711 23903 16717
rect 23845 16677 23857 16711
rect 23891 16708 23903 16711
rect 24118 16708 24124 16720
rect 23891 16680 24124 16708
rect 23891 16677 23903 16680
rect 23845 16671 23903 16677
rect 24118 16668 24124 16680
rect 24176 16708 24182 16720
rect 24857 16711 24915 16717
rect 24857 16708 24869 16711
rect 24176 16680 24869 16708
rect 24176 16668 24182 16680
rect 24857 16677 24869 16680
rect 24903 16677 24915 16711
rect 24857 16671 24915 16677
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16609 18107 16643
rect 18049 16603 18107 16609
rect 18601 16643 18659 16649
rect 18601 16609 18613 16643
rect 18647 16640 18659 16643
rect 19150 16640 19156 16652
rect 18647 16612 19156 16640
rect 18647 16609 18659 16612
rect 18601 16603 18659 16609
rect 11756 16544 12388 16572
rect 12437 16575 12495 16581
rect 11756 16532 11762 16544
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 11974 16464 11980 16516
rect 12032 16504 12038 16516
rect 12452 16504 12480 16535
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 18616 16572 18644 16603
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 19978 16640 19984 16652
rect 19751 16612 19984 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 21174 16600 21180 16652
rect 21232 16640 21238 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 21232 16612 21281 16640
rect 21232 16600 21238 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 22646 16640 22652 16652
rect 22607 16612 22652 16640
rect 21269 16603 21327 16609
rect 22646 16600 22652 16612
rect 22704 16640 22710 16652
rect 23385 16643 23443 16649
rect 23385 16640 23397 16643
rect 22704 16612 23397 16640
rect 22704 16600 22710 16612
rect 23385 16609 23397 16612
rect 23431 16609 23443 16643
rect 25038 16640 25044 16652
rect 23385 16603 23443 16609
rect 24780 16612 25044 16640
rect 18472 16544 18644 16572
rect 18693 16575 18751 16581
rect 18472 16532 18478 16544
rect 18693 16541 18705 16575
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 12032 16476 12480 16504
rect 12032 16464 12038 16476
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 18708 16504 18736 16535
rect 18288 16476 18736 16504
rect 18288 16464 18294 16476
rect 21266 16464 21272 16516
rect 21324 16504 21330 16516
rect 21376 16504 21404 16535
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 22922 16572 22928 16584
rect 21508 16544 21553 16572
rect 22883 16544 22928 16572
rect 21508 16532 21514 16544
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 24210 16532 24216 16584
rect 24268 16572 24274 16584
rect 24397 16575 24455 16581
rect 24397 16572 24409 16575
rect 24268 16544 24409 16572
rect 24268 16532 24274 16544
rect 24397 16541 24409 16544
rect 24443 16541 24455 16575
rect 24397 16535 24455 16541
rect 24489 16575 24547 16581
rect 24489 16541 24501 16575
rect 24535 16572 24547 16575
rect 24780 16572 24808 16612
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 24535 16544 24808 16572
rect 24535 16541 24547 16544
rect 24489 16535 24547 16541
rect 21324 16476 21404 16504
rect 21324 16464 21330 16476
rect 23566 16464 23572 16516
rect 23624 16504 23630 16516
rect 24504 16504 24532 16535
rect 23624 16476 24532 16504
rect 23624 16464 23630 16476
rect 12345 16439 12403 16445
rect 12345 16405 12357 16439
rect 12391 16436 12403 16439
rect 12802 16436 12808 16448
rect 12391 16408 12808 16436
rect 12391 16405 12403 16408
rect 12345 16399 12403 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 13814 16436 13820 16448
rect 13775 16408 13820 16436
rect 13814 16396 13820 16408
rect 13872 16436 13878 16448
rect 14093 16439 14151 16445
rect 14093 16436 14105 16439
rect 13872 16408 14105 16436
rect 13872 16396 13878 16408
rect 14093 16405 14105 16408
rect 14139 16405 14151 16439
rect 19886 16436 19892 16448
rect 19847 16408 19892 16436
rect 14093 16399 14151 16405
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 20898 16436 20904 16448
rect 20859 16408 20904 16436
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 22002 16436 22008 16448
rect 21963 16408 22008 16436
rect 22002 16396 22008 16408
rect 22060 16436 22066 16448
rect 22186 16436 22192 16448
rect 22060 16408 22192 16436
rect 22060 16396 22066 16408
rect 22186 16396 22192 16408
rect 22244 16396 22250 16448
rect 24857 16439 24915 16445
rect 24857 16405 24869 16439
rect 24903 16436 24915 16439
rect 25038 16436 25044 16448
rect 24903 16408 25044 16436
rect 24903 16405 24915 16408
rect 24857 16399 24915 16405
rect 25038 16396 25044 16408
rect 25096 16396 25102 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 11238 16232 11244 16244
rect 11199 16204 11244 16232
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 11698 16232 11704 16244
rect 11659 16204 11704 16232
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 13538 16232 13544 16244
rect 12492 16204 12537 16232
rect 13499 16204 13544 16232
rect 12492 16192 12498 16204
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 15562 16232 15568 16244
rect 15427 16204 15568 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 15749 16235 15807 16241
rect 15749 16201 15761 16235
rect 15795 16232 15807 16235
rect 16206 16232 16212 16244
rect 15795 16204 16212 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 16206 16192 16212 16204
rect 16264 16192 16270 16244
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 18288 16204 19441 16232
rect 18288 16192 18294 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 22922 16192 22928 16244
rect 22980 16232 22986 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22980 16204 23029 16232
rect 22980 16192 22986 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 23017 16195 23075 16201
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 23566 16232 23572 16244
rect 23523 16204 23572 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 24029 16235 24087 16241
rect 24029 16201 24041 16235
rect 24075 16232 24087 16235
rect 24210 16232 24216 16244
rect 24075 16204 24216 16232
rect 24075 16201 24087 16204
rect 24029 16195 24087 16201
rect 24210 16192 24216 16204
rect 24268 16232 24274 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 24268 16204 25053 16232
rect 24268 16192 24274 16204
rect 25041 16201 25053 16204
rect 25087 16201 25099 16235
rect 25041 16195 25099 16201
rect 14001 16167 14059 16173
rect 14001 16164 14013 16167
rect 12912 16136 14013 16164
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 12912 16105 12940 16136
rect 14001 16133 14013 16136
rect 14047 16133 14059 16167
rect 16761 16167 16819 16173
rect 16761 16164 16773 16167
rect 14001 16127 14059 16133
rect 16224 16136 16773 16164
rect 12897 16099 12955 16105
rect 12897 16096 12909 16099
rect 12860 16068 12909 16096
rect 12860 16056 12866 16068
rect 12897 16065 12909 16068
rect 12943 16065 12955 16099
rect 13078 16096 13084 16108
rect 13039 16068 13084 16096
rect 12897 16059 12955 16065
rect 13078 16056 13084 16068
rect 13136 16056 13142 16108
rect 14458 16096 14464 16108
rect 14419 16068 14464 16096
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14568 16028 14596 16059
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 16224 16105 16252 16136
rect 16761 16133 16773 16136
rect 16807 16133 16819 16167
rect 16761 16127 16819 16133
rect 22649 16167 22707 16173
rect 22649 16133 22661 16167
rect 22695 16164 22707 16167
rect 23382 16164 23388 16176
rect 22695 16136 23388 16164
rect 22695 16133 22707 16136
rect 22649 16127 22707 16133
rect 23382 16124 23388 16136
rect 23440 16124 23446 16176
rect 24946 16124 24952 16176
rect 25004 16164 25010 16176
rect 25409 16167 25467 16173
rect 25409 16164 25421 16167
rect 25004 16136 25421 16164
rect 25004 16124 25010 16136
rect 25409 16133 25421 16136
rect 25455 16133 25467 16167
rect 25409 16127 25467 16133
rect 16209 16099 16267 16105
rect 16209 16096 16221 16099
rect 15344 16068 16221 16096
rect 15344 16056 15350 16068
rect 16209 16065 16221 16068
rect 16255 16065 16267 16099
rect 16209 16059 16267 16065
rect 16298 16056 16304 16108
rect 16356 16096 16362 16108
rect 16393 16099 16451 16105
rect 16393 16096 16405 16099
rect 16356 16068 16405 16096
rect 16356 16056 16362 16068
rect 16393 16065 16405 16068
rect 16439 16096 16451 16099
rect 16482 16096 16488 16108
rect 16439 16068 16488 16096
rect 16439 16065 16451 16068
rect 16393 16059 16451 16065
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 23198 16056 23204 16108
rect 23256 16096 23262 16108
rect 23845 16099 23903 16105
rect 23845 16096 23857 16099
rect 23256 16068 23857 16096
rect 23256 16056 23262 16068
rect 23845 16065 23857 16068
rect 23891 16065 23903 16099
rect 23845 16059 23903 16065
rect 13872 16000 14596 16028
rect 13872 15988 13878 16000
rect 17770 15988 17776 16040
rect 17828 16028 17834 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17828 16000 18061 16028
rect 17828 15988 17834 16000
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 20070 16028 20076 16040
rect 18095 16000 20076 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 20070 15988 20076 16000
rect 20128 16028 20134 16040
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 20128 16000 20269 16028
rect 20128 15988 20134 16000
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 22278 16028 22284 16040
rect 22239 16000 22284 16028
rect 20257 15991 20315 15997
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 16028 22523 16031
rect 22922 16028 22928 16040
rect 22511 16000 22928 16028
rect 22511 15997 22523 16000
rect 22465 15991 22523 15997
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 23860 16028 23888 16059
rect 24026 16056 24032 16108
rect 24084 16096 24090 16108
rect 24394 16096 24400 16108
rect 24084 16068 24400 16096
rect 24084 16056 24090 16068
rect 24394 16056 24400 16068
rect 24452 16096 24458 16108
rect 24581 16099 24639 16105
rect 24581 16096 24593 16099
rect 24452 16068 24593 16096
rect 24452 16056 24458 16068
rect 24581 16065 24593 16068
rect 24627 16065 24639 16099
rect 25590 16096 25596 16108
rect 25551 16068 25596 16096
rect 24581 16059 24639 16065
rect 25590 16056 25596 16068
rect 25648 16056 25654 16108
rect 24489 16031 24547 16037
rect 24489 16028 24501 16031
rect 23860 16000 24501 16028
rect 24489 15997 24501 16000
rect 24535 15997 24547 16031
rect 24489 15991 24547 15997
rect 11882 15920 11888 15972
rect 11940 15960 11946 15972
rect 12253 15963 12311 15969
rect 12253 15960 12265 15963
rect 11940 15932 12265 15960
rect 11940 15920 11946 15932
rect 12253 15929 12265 15932
rect 12299 15960 12311 15963
rect 13078 15960 13084 15972
rect 12299 15932 13084 15960
rect 12299 15929 12311 15932
rect 12253 15923 12311 15929
rect 13078 15920 13084 15932
rect 13136 15920 13142 15972
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 18316 15963 18374 15969
rect 18316 15960 18328 15963
rect 18196 15932 18328 15960
rect 18196 15920 18202 15932
rect 18316 15929 18328 15932
rect 18362 15960 18374 15963
rect 20524 15963 20582 15969
rect 18362 15932 20208 15960
rect 18362 15929 18374 15932
rect 18316 15923 18374 15929
rect 10965 15895 11023 15901
rect 10965 15861 10977 15895
rect 11011 15892 11023 15895
rect 11606 15892 11612 15904
rect 11011 15864 11612 15892
rect 11011 15861 11023 15864
rect 10965 15855 11023 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 12584 15864 12817 15892
rect 12584 15852 12590 15864
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 12805 15855 12863 15861
rect 12894 15852 12900 15904
rect 12952 15892 12958 15904
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 12952 15864 13829 15892
rect 12952 15852 12958 15864
rect 13817 15861 13829 15864
rect 13863 15892 13875 15895
rect 14369 15895 14427 15901
rect 14369 15892 14381 15895
rect 13863 15864 14381 15892
rect 13863 15861 13875 15864
rect 13817 15855 13875 15861
rect 14369 15861 14381 15864
rect 14415 15861 14427 15895
rect 16114 15892 16120 15904
rect 16075 15864 16120 15892
rect 14369 15855 14427 15861
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 17494 15892 17500 15904
rect 17455 15864 17500 15892
rect 17494 15852 17500 15864
rect 17552 15852 17558 15904
rect 17865 15895 17923 15901
rect 17865 15861 17877 15895
rect 17911 15892 17923 15895
rect 19150 15892 19156 15904
rect 17911 15864 19156 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 19797 15895 19855 15901
rect 19797 15861 19809 15895
rect 19843 15892 19855 15895
rect 19978 15892 19984 15904
rect 19843 15864 19984 15892
rect 19843 15861 19855 15864
rect 19797 15855 19855 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20180 15901 20208 15932
rect 20524 15929 20536 15963
rect 20570 15960 20582 15963
rect 20622 15960 20628 15972
rect 20570 15932 20628 15960
rect 20570 15929 20582 15932
rect 20524 15923 20582 15929
rect 20622 15920 20628 15932
rect 20680 15920 20686 15972
rect 21266 15920 21272 15972
rect 21324 15960 21330 15972
rect 21913 15963 21971 15969
rect 21913 15960 21925 15963
rect 21324 15932 21925 15960
rect 21324 15920 21330 15932
rect 21913 15929 21925 15932
rect 21959 15929 21971 15963
rect 21913 15923 21971 15929
rect 23842 15920 23848 15972
rect 23900 15960 23906 15972
rect 24210 15960 24216 15972
rect 23900 15932 24216 15960
rect 23900 15920 23906 15932
rect 24210 15920 24216 15932
rect 24268 15920 24274 15972
rect 20165 15895 20223 15901
rect 20165 15861 20177 15895
rect 20211 15892 20223 15895
rect 21450 15892 21456 15904
rect 20211 15864 21456 15892
rect 20211 15861 20223 15864
rect 20165 15855 20223 15861
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 21542 15852 21548 15904
rect 21600 15892 21606 15904
rect 21637 15895 21695 15901
rect 21637 15892 21649 15895
rect 21600 15864 21649 15892
rect 21600 15852 21606 15864
rect 21637 15861 21649 15864
rect 21683 15861 21695 15895
rect 21637 15855 21695 15861
rect 21726 15852 21732 15904
rect 21784 15892 21790 15904
rect 24397 15895 24455 15901
rect 24397 15892 24409 15895
rect 21784 15864 24409 15892
rect 21784 15852 21790 15864
rect 24397 15861 24409 15864
rect 24443 15892 24455 15895
rect 24762 15892 24768 15904
rect 24443 15864 24768 15892
rect 24443 15861 24455 15864
rect 24397 15855 24455 15861
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 13136 15660 13277 15688
rect 13136 15648 13142 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 14001 15691 14059 15697
rect 14001 15657 14013 15691
rect 14047 15688 14059 15691
rect 14182 15688 14188 15700
rect 14047 15660 14188 15688
rect 14047 15657 14059 15660
rect 14001 15651 14059 15657
rect 14182 15648 14188 15660
rect 14240 15688 14246 15700
rect 14642 15688 14648 15700
rect 14240 15660 14648 15688
rect 14240 15648 14246 15660
rect 14642 15648 14648 15660
rect 14700 15688 14706 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 14700 15660 15025 15688
rect 14700 15648 14706 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 15013 15651 15071 15657
rect 16114 15648 16120 15700
rect 16172 15688 16178 15700
rect 16577 15691 16635 15697
rect 16577 15688 16589 15691
rect 16172 15660 16589 15688
rect 16172 15648 16178 15660
rect 16577 15657 16589 15660
rect 16623 15688 16635 15691
rect 17862 15688 17868 15700
rect 16623 15660 17868 15688
rect 16623 15657 16635 15660
rect 16577 15651 16635 15657
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 18138 15688 18144 15700
rect 18099 15660 18144 15688
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 19242 15688 19248 15700
rect 19203 15660 19248 15688
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 20438 15688 20444 15700
rect 20395 15660 20444 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 20438 15648 20444 15660
rect 20496 15688 20502 15700
rect 20622 15688 20628 15700
rect 20496 15660 20628 15688
rect 20496 15648 20502 15660
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 24394 15688 24400 15700
rect 22060 15660 22140 15688
rect 24355 15660 24400 15688
rect 22060 15648 22066 15660
rect 15657 15623 15715 15629
rect 15657 15589 15669 15623
rect 15703 15620 15715 15623
rect 16022 15620 16028 15632
rect 15703 15592 16028 15620
rect 15703 15589 15715 15592
rect 15657 15583 15715 15589
rect 16022 15580 16028 15592
rect 16080 15580 16086 15632
rect 16209 15623 16267 15629
rect 16209 15589 16221 15623
rect 16255 15620 16267 15623
rect 16298 15620 16304 15632
rect 16255 15592 16304 15620
rect 16255 15589 16267 15592
rect 16209 15583 16267 15589
rect 16298 15580 16304 15592
rect 16356 15580 16362 15632
rect 17126 15620 17132 15632
rect 17039 15592 17132 15620
rect 17126 15580 17132 15592
rect 17184 15620 17190 15632
rect 17310 15620 17316 15632
rect 17184 15592 17316 15620
rect 17184 15580 17190 15592
rect 17310 15580 17316 15592
rect 17368 15580 17374 15632
rect 19978 15580 19984 15632
rect 20036 15620 20042 15632
rect 21361 15623 21419 15629
rect 21361 15620 21373 15623
rect 20036 15592 21373 15620
rect 20036 15580 20042 15592
rect 21361 15589 21373 15592
rect 21407 15589 21419 15623
rect 21361 15583 21419 15589
rect 11974 15552 11980 15564
rect 11900 15524 11980 15552
rect 11900 15493 11928 15524
rect 11974 15512 11980 15524
rect 12032 15512 12038 15564
rect 12158 15561 12164 15564
rect 12152 15552 12164 15561
rect 12119 15524 12164 15552
rect 12152 15515 12164 15524
rect 12158 15512 12164 15515
rect 12216 15512 12222 15564
rect 15286 15512 15292 15564
rect 15344 15552 15350 15564
rect 15381 15555 15439 15561
rect 15381 15552 15393 15555
rect 15344 15524 15393 15552
rect 15344 15512 15350 15524
rect 15381 15521 15393 15524
rect 15427 15521 15439 15555
rect 15381 15515 15439 15521
rect 16482 15512 16488 15564
rect 16540 15552 16546 15564
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 16540 15524 17049 15552
rect 16540 15512 16546 15524
rect 17037 15521 17049 15524
rect 17083 15552 17095 15555
rect 18233 15555 18291 15561
rect 18233 15552 18245 15555
rect 17083 15524 18245 15552
rect 17083 15521 17095 15524
rect 17037 15515 17095 15521
rect 18233 15521 18245 15524
rect 18279 15521 18291 15555
rect 18233 15515 18291 15521
rect 19518 15512 19524 15564
rect 19576 15552 19582 15564
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 19576 15524 19625 15552
rect 19576 15512 19582 15524
rect 19613 15521 19625 15524
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 20254 15552 20260 15564
rect 19751 15524 20260 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 11885 15487 11943 15493
rect 11885 15484 11897 15487
rect 11716 15456 11897 15484
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 10962 15348 10968 15360
rect 10919 15320 10968 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11716 15357 11744 15456
rect 11885 15453 11897 15456
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13872 15456 14105 15484
rect 13872 15444 13878 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 19153 15487 19211 15493
rect 19153 15453 19165 15487
rect 19199 15484 19211 15487
rect 19720 15484 19748 15515
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 20898 15512 20904 15564
rect 20956 15552 20962 15564
rect 21085 15555 21143 15561
rect 21085 15552 21097 15555
rect 20956 15524 21097 15552
rect 20956 15512 20962 15524
rect 21085 15521 21097 15524
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 19199 15456 19748 15484
rect 19199 15453 19211 15456
rect 19153 15447 19211 15453
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 17236 15416 17264 15447
rect 19794 15444 19800 15496
rect 19852 15484 19858 15496
rect 19852 15456 19897 15484
rect 19852 15444 19858 15456
rect 20070 15444 20076 15496
rect 20128 15484 20134 15496
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 20128 15456 21833 15484
rect 20128 15444 20134 15456
rect 21821 15453 21833 15456
rect 21867 15484 21879 15487
rect 22112 15484 22140 15660
rect 24394 15648 24400 15660
rect 24452 15648 24458 15700
rect 24670 15648 24676 15700
rect 24728 15688 24734 15700
rect 25038 15688 25044 15700
rect 24728 15660 25044 15688
rect 24728 15648 24734 15660
rect 25038 15648 25044 15660
rect 25096 15688 25102 15700
rect 25593 15691 25651 15697
rect 25593 15688 25605 15691
rect 25096 15660 25605 15688
rect 25096 15648 25102 15660
rect 25593 15657 25605 15660
rect 25639 15657 25651 15691
rect 25593 15651 25651 15657
rect 22640 15555 22698 15561
rect 22640 15521 22652 15555
rect 22686 15552 22698 15555
rect 23014 15552 23020 15564
rect 22686 15524 23020 15552
rect 22686 15521 22698 15524
rect 22640 15515 22698 15521
rect 23014 15512 23020 15524
rect 23072 15512 23078 15564
rect 24946 15552 24952 15564
rect 24907 15524 24952 15552
rect 24946 15512 24952 15524
rect 25004 15552 25010 15564
rect 26142 15552 26148 15564
rect 25004 15524 26148 15552
rect 25004 15512 25010 15524
rect 26142 15512 26148 15524
rect 26200 15512 26206 15564
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 21867 15456 22293 15484
rect 21867 15453 21879 15456
rect 21821 15447 21879 15453
rect 22281 15453 22293 15456
rect 22327 15484 22339 15487
rect 22373 15487 22431 15493
rect 22373 15484 22385 15487
rect 22327 15456 22385 15484
rect 22327 15453 22339 15456
rect 22281 15447 22339 15453
rect 22373 15453 22385 15456
rect 22419 15453 22431 15487
rect 25038 15484 25044 15496
rect 24999 15456 25044 15484
rect 22373 15447 22431 15453
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 25130 15444 25136 15496
rect 25188 15484 25194 15496
rect 25188 15456 25233 15484
rect 25188 15444 25194 15456
rect 18230 15416 18236 15428
rect 15620 15388 18236 15416
rect 15620 15376 15626 15388
rect 18230 15376 18236 15388
rect 18288 15416 18294 15428
rect 18693 15419 18751 15425
rect 18693 15416 18705 15419
rect 18288 15388 18705 15416
rect 18288 15376 18294 15388
rect 18693 15385 18705 15388
rect 18739 15385 18751 15419
rect 18693 15379 18751 15385
rect 23474 15376 23480 15428
rect 23532 15416 23538 15428
rect 24581 15419 24639 15425
rect 24581 15416 24593 15419
rect 23532 15388 24593 15416
rect 23532 15376 23538 15388
rect 24581 15385 24593 15388
rect 24627 15385 24639 15419
rect 24581 15379 24639 15385
rect 11333 15351 11391 15357
rect 11333 15348 11345 15351
rect 11204 15320 11345 15348
rect 11204 15308 11210 15320
rect 11333 15317 11345 15320
rect 11379 15348 11391 15351
rect 11701 15351 11759 15357
rect 11701 15348 11713 15351
rect 11379 15320 11713 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11701 15317 11713 15320
rect 11747 15317 11759 15351
rect 13538 15348 13544 15360
rect 13499 15320 13544 15348
rect 11701 15311 11759 15317
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 16669 15351 16727 15357
rect 16669 15317 16681 15351
rect 16715 15348 16727 15351
rect 16758 15348 16764 15360
rect 16715 15320 16764 15348
rect 16715 15317 16727 15320
rect 16669 15311 16727 15317
rect 16758 15308 16764 15320
rect 16816 15348 16822 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 16816 15320 17693 15348
rect 16816 15308 16822 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 20806 15348 20812 15360
rect 20763 15320 20812 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 23290 15308 23296 15360
rect 23348 15348 23354 15360
rect 23753 15351 23811 15357
rect 23753 15348 23765 15351
rect 23348 15320 23765 15348
rect 23348 15308 23354 15320
rect 23753 15317 23765 15320
rect 23799 15317 23811 15351
rect 23753 15311 23811 15317
rect 24121 15351 24179 15357
rect 24121 15317 24133 15351
rect 24167 15348 24179 15351
rect 24762 15348 24768 15360
rect 24167 15320 24768 15348
rect 24167 15317 24179 15320
rect 24121 15311 24179 15317
rect 24762 15308 24768 15320
rect 24820 15348 24826 15360
rect 26050 15348 26056 15360
rect 24820 15320 26056 15348
rect 24820 15308 24826 15320
rect 26050 15308 26056 15320
rect 26108 15308 26114 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 12621 15147 12679 15153
rect 12621 15144 12633 15147
rect 12584 15116 12633 15144
rect 12584 15104 12590 15116
rect 12621 15113 12633 15116
rect 12667 15113 12679 15147
rect 12621 15107 12679 15113
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 15841 15147 15899 15153
rect 15841 15144 15853 15147
rect 15528 15116 15853 15144
rect 15528 15104 15534 15116
rect 15841 15113 15853 15116
rect 15887 15113 15899 15147
rect 15841 15107 15899 15113
rect 16301 15147 16359 15153
rect 16301 15113 16313 15147
rect 16347 15144 16359 15147
rect 16482 15144 16488 15156
rect 16347 15116 16488 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 18230 15104 18236 15156
rect 18288 15144 18294 15156
rect 18598 15144 18604 15156
rect 18288 15116 18604 15144
rect 18288 15104 18294 15116
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 20898 15104 20904 15156
rect 20956 15144 20962 15156
rect 21545 15147 21603 15153
rect 21545 15144 21557 15147
rect 20956 15116 21557 15144
rect 20956 15104 20962 15116
rect 21545 15113 21557 15116
rect 21591 15113 21603 15147
rect 21545 15107 21603 15113
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 23382 15144 23388 15156
rect 22235 15116 23388 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 15562 15076 15568 15088
rect 15523 15048 15568 15076
rect 15562 15036 15568 15048
rect 15620 15036 15626 15088
rect 16390 15076 16396 15088
rect 16351 15048 16396 15076
rect 16390 15036 16396 15048
rect 16448 15036 16454 15088
rect 21269 15079 21327 15085
rect 21269 15045 21281 15079
rect 21315 15076 21327 15079
rect 21450 15076 21456 15088
rect 21315 15048 21456 15076
rect 21315 15045 21327 15048
rect 21269 15039 21327 15045
rect 21450 15036 21456 15048
rect 21508 15036 21514 15088
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 15008 10747 15011
rect 11422 15008 11428 15020
rect 10735 14980 11428 15008
rect 10735 14977 10747 14980
rect 10689 14971 10747 14977
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 12158 15008 12164 15020
rect 11931 14980 12164 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12158 14968 12164 14980
rect 12216 15008 12222 15020
rect 13173 15011 13231 15017
rect 13173 15008 13185 15011
rect 12216 14980 13185 15008
rect 12216 14968 12222 14980
rect 13173 14977 13185 14980
rect 13219 15008 13231 15011
rect 13630 15008 13636 15020
rect 13219 14980 13636 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 14182 15008 14188 15020
rect 14143 14980 14188 15008
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 16298 14968 16304 15020
rect 16356 15008 16362 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16356 14980 16957 15008
rect 16356 14968 16362 14980
rect 16945 14977 16957 14980
rect 16991 14977 17003 15011
rect 18598 15008 18604 15020
rect 18559 14980 18604 15008
rect 16945 14971 17003 14977
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 11112 14912 11253 14940
rect 11112 14900 11118 14912
rect 11241 14909 11253 14912
rect 11287 14940 11299 14943
rect 12526 14940 12532 14952
rect 11287 14912 12532 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 12986 14940 12992 14952
rect 12899 14912 12992 14940
rect 12986 14900 12992 14912
rect 13044 14940 13050 14952
rect 13722 14940 13728 14952
rect 13044 14912 13728 14940
rect 13044 14900 13050 14912
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 16758 14940 16764 14952
rect 16719 14912 16764 14940
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 16850 14900 16856 14952
rect 16908 14940 16914 14952
rect 17862 14940 17868 14952
rect 16908 14912 17868 14940
rect 16908 14900 16914 14912
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 19889 14943 19947 14949
rect 19889 14909 19901 14943
rect 19935 14940 19947 14943
rect 19978 14940 19984 14952
rect 19935 14912 19984 14940
rect 19935 14909 19947 14912
rect 19889 14903 19947 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 22296 14949 22324 15116
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 25130 15144 25136 15156
rect 23952 15116 25136 15144
rect 23014 15076 23020 15088
rect 22975 15048 23020 15076
rect 23014 15036 23020 15048
rect 23072 15076 23078 15088
rect 23952 15085 23980 15116
rect 25130 15104 25136 15116
rect 25188 15144 25194 15156
rect 25501 15147 25559 15153
rect 25501 15144 25513 15147
rect 25188 15116 25513 15144
rect 25188 15104 25194 15116
rect 25501 15113 25513 15116
rect 25547 15113 25559 15147
rect 26234 15144 26240 15156
rect 26195 15116 26240 15144
rect 25501 15107 25559 15113
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 23937 15079 23995 15085
rect 23937 15076 23949 15079
rect 23072 15048 23949 15076
rect 23072 15036 23078 15048
rect 23937 15045 23949 15048
rect 23983 15045 23995 15079
rect 23937 15039 23995 15045
rect 22462 15008 22468 15020
rect 22423 14980 22468 15008
rect 22462 14968 22468 14980
rect 22520 14968 22526 15020
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 24121 14943 24179 14949
rect 24121 14909 24133 14943
rect 24167 14940 24179 14943
rect 24670 14940 24676 14952
rect 24167 14912 24676 14940
rect 24167 14909 24179 14912
rect 24121 14903 24179 14909
rect 24670 14900 24676 14912
rect 24728 14900 24734 14952
rect 10321 14875 10379 14881
rect 10321 14841 10333 14875
rect 10367 14872 10379 14875
rect 11149 14875 11207 14881
rect 11149 14872 11161 14875
rect 10367 14844 11161 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 11149 14841 11161 14844
rect 11195 14872 11207 14875
rect 12342 14872 12348 14884
rect 11195 14844 12348 14872
rect 11195 14841 11207 14844
rect 11149 14835 11207 14841
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 14093 14875 14151 14881
rect 14093 14841 14105 14875
rect 14139 14872 14151 14875
rect 14274 14872 14280 14884
rect 14139 14844 14280 14872
rect 14139 14841 14151 14844
rect 14093 14835 14151 14841
rect 14274 14832 14280 14844
rect 14332 14872 14338 14884
rect 14430 14875 14488 14881
rect 14430 14872 14442 14875
rect 14332 14844 14442 14872
rect 14332 14832 14338 14844
rect 14430 14841 14442 14844
rect 14476 14841 14488 14875
rect 18417 14875 18475 14881
rect 18417 14872 18429 14875
rect 14430 14835 14488 14841
rect 17788 14844 18429 14872
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 12299 14776 13093 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 13081 14773 13093 14776
rect 13127 14804 13139 14807
rect 13262 14804 13268 14816
rect 13127 14776 13268 14804
rect 13127 14773 13139 14776
rect 13081 14767 13139 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 17310 14764 17316 14816
rect 17368 14804 17374 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 17368 14776 17417 14804
rect 17368 14764 17374 14776
rect 17405 14773 17417 14776
rect 17451 14773 17463 14807
rect 17405 14767 17463 14773
rect 17494 14764 17500 14816
rect 17552 14804 17558 14816
rect 17788 14813 17816 14844
rect 18417 14841 18429 14844
rect 18463 14841 18475 14875
rect 18417 14835 18475 14841
rect 19705 14875 19763 14881
rect 19705 14841 19717 14875
rect 19751 14872 19763 14875
rect 19794 14872 19800 14884
rect 19751 14844 19800 14872
rect 19751 14841 19763 14844
rect 19705 14835 19763 14841
rect 19794 14832 19800 14844
rect 19852 14872 19858 14884
rect 20156 14875 20214 14881
rect 20156 14872 20168 14875
rect 19852 14844 20168 14872
rect 19852 14832 19858 14844
rect 20156 14841 20168 14844
rect 20202 14872 20214 14875
rect 21542 14872 21548 14884
rect 20202 14844 21548 14872
rect 20202 14841 20214 14844
rect 20156 14835 20214 14841
rect 21542 14832 21548 14844
rect 21600 14832 21606 14884
rect 24394 14881 24400 14884
rect 23477 14875 23535 14881
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 24388 14872 24400 14881
rect 23523 14844 24400 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 24388 14835 24400 14844
rect 24394 14832 24400 14835
rect 24452 14832 24458 14884
rect 25038 14832 25044 14884
rect 25096 14872 25102 14884
rect 25777 14875 25835 14881
rect 25777 14872 25789 14875
rect 25096 14844 25789 14872
rect 25096 14832 25102 14844
rect 25777 14841 25789 14844
rect 25823 14841 25835 14875
rect 25777 14835 25835 14841
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 17552 14776 17785 14804
rect 17552 14764 17558 14776
rect 17773 14773 17785 14776
rect 17819 14773 17831 14807
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 17773 14767 17831 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18506 14804 18512 14816
rect 18467 14776 18512 14804
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 19337 14807 19395 14813
rect 19337 14773 19349 14807
rect 19383 14804 19395 14807
rect 19518 14804 19524 14816
rect 19383 14776 19524 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 12713 14603 12771 14609
rect 12713 14569 12725 14603
rect 12759 14600 12771 14603
rect 12986 14600 12992 14612
rect 12759 14572 12992 14600
rect 12759 14569 12771 14572
rect 12713 14563 12771 14569
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 15102 14600 15108 14612
rect 13679 14572 15108 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 16298 14560 16304 14612
rect 16356 14600 16362 14612
rect 16393 14603 16451 14609
rect 16393 14600 16405 14603
rect 16356 14572 16405 14600
rect 16356 14560 16362 14572
rect 16393 14569 16405 14572
rect 16439 14569 16451 14603
rect 16393 14563 16451 14569
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 16632 14572 16681 14600
rect 16632 14560 16638 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 16669 14563 16727 14569
rect 20901 14603 20959 14609
rect 20901 14569 20913 14603
rect 20947 14600 20959 14603
rect 21266 14600 21272 14612
rect 20947 14572 21272 14600
rect 20947 14569 20959 14572
rect 20901 14563 20959 14569
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 21361 14603 21419 14609
rect 21361 14569 21373 14603
rect 21407 14600 21419 14603
rect 21634 14600 21640 14612
rect 21407 14572 21640 14600
rect 21407 14569 21419 14572
rect 21361 14563 21419 14569
rect 21634 14560 21640 14572
rect 21692 14600 21698 14612
rect 22465 14603 22523 14609
rect 22465 14600 22477 14603
rect 21692 14572 22477 14600
rect 21692 14560 21698 14572
rect 22465 14569 22477 14572
rect 22511 14569 22523 14603
rect 22465 14563 22523 14569
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 22612 14572 22845 14600
rect 22612 14560 22618 14572
rect 22833 14569 22845 14572
rect 22879 14600 22891 14603
rect 23382 14600 23388 14612
rect 22879 14572 23388 14600
rect 22879 14569 22891 14572
rect 22833 14563 22891 14569
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 24029 14603 24087 14609
rect 24029 14569 24041 14603
rect 24075 14600 24087 14603
rect 24946 14600 24952 14612
rect 24075 14572 24952 14600
rect 24075 14569 24087 14572
rect 24029 14563 24087 14569
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 11232 14535 11290 14541
rect 11232 14501 11244 14535
rect 11278 14532 11290 14535
rect 11882 14532 11888 14544
rect 11278 14504 11888 14532
rect 11278 14501 11290 14504
rect 11232 14495 11290 14501
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 13998 14532 14004 14544
rect 13959 14504 14004 14532
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 15746 14532 15752 14544
rect 15611 14504 15752 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 16117 14535 16175 14541
rect 16117 14501 16129 14535
rect 16163 14532 16175 14535
rect 16850 14532 16856 14544
rect 16163 14504 16856 14532
rect 16163 14501 16175 14504
rect 16117 14495 16175 14501
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 20806 14532 20812 14544
rect 19628 14504 20812 14532
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 10962 14464 10968 14476
rect 10551 14436 10968 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13228 14436 14105 14464
rect 13228 14424 13234 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 14642 14424 14648 14476
rect 14700 14464 14706 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 14700 14436 15301 14464
rect 14700 14424 14706 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 17017 14467 17075 14473
rect 17017 14464 17029 14467
rect 16632 14436 17029 14464
rect 16632 14424 16638 14436
rect 17017 14433 17029 14436
rect 17063 14433 17075 14467
rect 17017 14427 17075 14433
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19628 14473 19656 14504
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 22925 14535 22983 14541
rect 22925 14501 22937 14535
rect 22971 14532 22983 14535
rect 23014 14532 23020 14544
rect 22971 14504 23020 14532
rect 22971 14501 22983 14504
rect 22925 14495 22983 14501
rect 23014 14492 23020 14504
rect 23072 14492 23078 14544
rect 23750 14492 23756 14544
rect 23808 14532 23814 14544
rect 24489 14535 24547 14541
rect 24489 14532 24501 14535
rect 23808 14504 24501 14532
rect 23808 14492 23814 14504
rect 24489 14501 24501 14504
rect 24535 14501 24547 14535
rect 24489 14495 24547 14501
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 19484 14436 19625 14464
rect 19484 14424 19490 14436
rect 19613 14433 19625 14436
rect 19659 14433 19671 14467
rect 19613 14427 19671 14433
rect 19705 14467 19763 14473
rect 19705 14433 19717 14467
rect 19751 14464 19763 14467
rect 19978 14464 19984 14476
rect 19751 14436 19984 14464
rect 19751 14433 19763 14436
rect 19705 14427 19763 14433
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 20990 14424 20996 14476
rect 21048 14464 21054 14476
rect 21269 14467 21327 14473
rect 21269 14464 21281 14467
rect 21048 14436 21281 14464
rect 21048 14424 21054 14436
rect 21269 14433 21281 14436
rect 21315 14433 21327 14467
rect 21269 14427 21327 14433
rect 23934 14424 23940 14476
rect 23992 14464 23998 14476
rect 24397 14467 24455 14473
rect 24397 14464 24409 14467
rect 23992 14436 24409 14464
rect 23992 14424 23998 14436
rect 24397 14433 24409 14436
rect 24443 14464 24455 14467
rect 25590 14464 25596 14476
rect 24443 14436 25596 14464
rect 24443 14433 24455 14436
rect 24397 14427 24455 14433
rect 25590 14424 25596 14436
rect 25648 14424 25654 14476
rect 14182 14396 14188 14408
rect 14143 14368 14188 14396
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14396 16727 14399
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 16715 14368 16773 14396
rect 16715 14365 16727 14368
rect 16669 14359 16727 14365
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14396 20775 14399
rect 21542 14396 21548 14408
rect 20763 14368 21548 14396
rect 20763 14365 20775 14368
rect 20717 14359 20775 14365
rect 19153 14331 19211 14337
rect 19153 14297 19165 14331
rect 19199 14328 19211 14331
rect 19334 14328 19340 14340
rect 19199 14300 19340 14328
rect 19199 14297 19211 14300
rect 19153 14291 19211 14297
rect 19334 14288 19340 14300
rect 19392 14328 19398 14340
rect 19812 14328 19840 14359
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 23109 14399 23167 14405
rect 23109 14365 23121 14399
rect 23155 14396 23167 14399
rect 23290 14396 23296 14408
rect 23155 14368 23296 14396
rect 23155 14365 23167 14368
rect 23109 14359 23167 14365
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 24673 14399 24731 14405
rect 24673 14365 24685 14399
rect 24719 14396 24731 14399
rect 25133 14399 25191 14405
rect 25133 14396 25145 14399
rect 24719 14368 25145 14396
rect 24719 14365 24731 14368
rect 24673 14359 24731 14365
rect 25133 14365 25145 14368
rect 25179 14396 25191 14399
rect 25222 14396 25228 14408
rect 25179 14368 25228 14396
rect 25179 14365 25191 14368
rect 25133 14359 25191 14365
rect 19392 14300 19840 14328
rect 19392 14288 19398 14300
rect 21818 14288 21824 14340
rect 21876 14328 21882 14340
rect 22738 14328 22744 14340
rect 21876 14300 22744 14328
rect 21876 14288 21882 14300
rect 22738 14288 22744 14300
rect 22796 14288 22802 14340
rect 23937 14331 23995 14337
rect 23937 14297 23949 14331
rect 23983 14328 23995 14331
rect 24394 14328 24400 14340
rect 23983 14300 24400 14328
rect 23983 14297 23995 14300
rect 23937 14291 23995 14297
rect 24394 14288 24400 14300
rect 24452 14328 24458 14340
rect 24688 14328 24716 14359
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 24452 14300 24716 14328
rect 24452 14288 24458 14300
rect 10870 14260 10876 14272
rect 10831 14232 10876 14260
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 12342 14260 12348 14272
rect 12303 14232 12348 14260
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 13170 14260 13176 14272
rect 13131 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13446 14260 13452 14272
rect 13407 14232 13452 14260
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 14734 14260 14740 14272
rect 14695 14232 14740 14260
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 15378 14220 15384 14272
rect 15436 14260 15442 14272
rect 15838 14260 15844 14272
rect 15436 14232 15844 14260
rect 15436 14220 15442 14232
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 18141 14263 18199 14269
rect 18141 14260 18153 14263
rect 18012 14232 18153 14260
rect 18012 14220 18018 14232
rect 18141 14229 18153 14232
rect 18187 14260 18199 14263
rect 18417 14263 18475 14269
rect 18417 14260 18429 14263
rect 18187 14232 18429 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 18417 14229 18429 14232
rect 18463 14260 18475 14263
rect 18598 14260 18604 14272
rect 18463 14232 18604 14260
rect 18463 14229 18475 14232
rect 18417 14223 18475 14229
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 20349 14263 20407 14269
rect 20349 14229 20361 14263
rect 20395 14260 20407 14263
rect 20806 14260 20812 14272
rect 20395 14232 20812 14260
rect 20395 14229 20407 14232
rect 20349 14223 20407 14229
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 22097 14263 22155 14269
rect 22097 14229 22109 14263
rect 22143 14260 22155 14263
rect 22554 14260 22560 14272
rect 22143 14232 22560 14260
rect 22143 14229 22155 14232
rect 22097 14223 22155 14229
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 23566 14260 23572 14272
rect 23527 14232 23572 14260
rect 23566 14220 23572 14232
rect 23624 14220 23630 14272
rect 25130 14220 25136 14272
rect 25188 14260 25194 14272
rect 25409 14263 25467 14269
rect 25409 14260 25421 14263
rect 25188 14232 25421 14260
rect 25188 14220 25194 14232
rect 25409 14229 25421 14232
rect 25455 14229 25467 14263
rect 25409 14223 25467 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 11882 14056 11888 14068
rect 11843 14028 11888 14056
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 13228 14028 13645 14056
rect 13228 14016 13234 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 14182 14016 14188 14068
rect 14240 14016 14246 14068
rect 14642 14056 14648 14068
rect 14603 14028 14648 14056
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14056 15163 14059
rect 15562 14056 15568 14068
rect 15151 14028 15568 14056
rect 15151 14025 15163 14028
rect 15105 14019 15163 14025
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 19334 14056 19340 14068
rect 17911 14028 19340 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 20070 14056 20076 14068
rect 20031 14028 20076 14056
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 20254 14056 20260 14068
rect 20215 14028 20260 14056
rect 20254 14016 20260 14028
rect 20312 14016 20318 14068
rect 21361 14059 21419 14065
rect 21361 14025 21373 14059
rect 21407 14056 21419 14059
rect 21542 14056 21548 14068
rect 21407 14028 21548 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 23382 14056 23388 14068
rect 23343 14028 23388 14056
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 23750 14016 23756 14068
rect 23808 14056 23814 14068
rect 24029 14059 24087 14065
rect 24029 14056 24041 14059
rect 23808 14028 24041 14056
rect 23808 14016 23814 14028
rect 24029 14025 24041 14028
rect 24075 14025 24087 14059
rect 24029 14019 24087 14025
rect 24581 14059 24639 14065
rect 24581 14025 24593 14059
rect 24627 14056 24639 14059
rect 25038 14056 25044 14068
rect 24627 14028 25044 14056
rect 24627 14025 24639 14028
rect 24581 14019 24639 14025
rect 25038 14016 25044 14028
rect 25096 14016 25102 14068
rect 25590 14056 25596 14068
rect 25551 14028 25596 14056
rect 25590 14016 25596 14028
rect 25648 14016 25654 14068
rect 9401 13991 9459 13997
rect 9401 13957 9413 13991
rect 9447 13988 9459 13991
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 9447 13960 10793 13988
rect 9447 13957 9459 13960
rect 9401 13951 9459 13957
rect 9508 13861 9536 13960
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 13541 13991 13599 13997
rect 13541 13957 13553 13991
rect 13587 13988 13599 13991
rect 14200 13988 14228 14016
rect 16574 13988 16580 14000
rect 13587 13960 14228 13988
rect 16535 13960 16580 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 16574 13948 16580 13960
rect 16632 13988 16638 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 16632 13960 17417 13988
rect 16632 13948 16638 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 19797 13991 19855 13997
rect 19797 13957 19809 13991
rect 19843 13988 19855 13991
rect 20438 13988 20444 14000
rect 19843 13960 20444 13988
rect 19843 13957 19855 13960
rect 19797 13951 19855 13957
rect 20438 13948 20444 13960
rect 20496 13988 20502 14000
rect 21818 13988 21824 14000
rect 20496 13960 20852 13988
rect 21779 13960 21824 13988
rect 20496 13948 20502 13960
rect 9766 13920 9772 13932
rect 9727 13892 9772 13920
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 10928 13892 11345 13920
rect 10928 13880 10934 13892
rect 11333 13889 11345 13892
rect 11379 13920 11391 13923
rect 11882 13920 11888 13932
rect 11379 13892 11888 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 13504 13892 14105 13920
rect 13504 13880 13510 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 15102 13920 15108 13932
rect 14231 13892 15108 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 10778 13852 10784 13864
rect 10367 13824 10784 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 10778 13812 10784 13824
rect 10836 13852 10842 13864
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 10836 13824 11253 13852
rect 10836 13812 10842 13824
rect 11241 13821 11253 13824
rect 11287 13821 11299 13855
rect 11241 13815 11299 13821
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 14200 13852 14228 13883
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 20824 13929 20852 13960
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 20809 13923 20867 13929
rect 20809 13889 20821 13923
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 13219 13824 14228 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 15470 13861 15476 13864
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 14424 13824 15209 13852
rect 14424 13812 14430 13824
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15464 13852 15476 13861
rect 15431 13824 15476 13852
rect 15197 13815 15255 13821
rect 15464 13815 15476 13824
rect 15470 13812 15476 13815
rect 15528 13812 15534 13864
rect 17954 13812 17960 13864
rect 18012 13812 18018 13864
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13852 18107 13855
rect 18874 13852 18880 13864
rect 18095 13824 18880 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 20824 13852 20852 13883
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 23290 13920 23296 13932
rect 22612 13892 22657 13920
rect 22848 13892 23296 13920
rect 22612 13880 22618 13892
rect 22848 13852 22876 13892
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 25222 13920 25228 13932
rect 25135 13892 25228 13920
rect 25222 13880 25228 13892
rect 25280 13920 25286 13932
rect 25590 13920 25596 13932
rect 25280 13892 25596 13920
rect 25280 13880 25286 13892
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 23014 13852 23020 13864
rect 20824 13824 22876 13852
rect 22975 13824 23020 13852
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 23934 13812 23940 13864
rect 23992 13852 23998 13864
rect 24397 13855 24455 13861
rect 24397 13852 24409 13855
rect 23992 13824 24409 13852
rect 23992 13812 23998 13824
rect 24397 13821 24409 13824
rect 24443 13852 24455 13855
rect 25038 13852 25044 13864
rect 24443 13824 24808 13852
rect 24999 13824 25044 13852
rect 24443 13821 24455 13824
rect 24397 13815 24455 13821
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 13630 13784 13636 13796
rect 12492 13756 13636 13784
rect 12492 13744 12498 13756
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 16758 13744 16764 13796
rect 16816 13784 16822 13796
rect 17972 13784 18000 13812
rect 18294 13787 18352 13793
rect 18294 13784 18306 13787
rect 16816 13756 18306 13784
rect 16816 13744 16822 13756
rect 18294 13753 18306 13756
rect 18340 13753 18352 13787
rect 18294 13747 18352 13753
rect 20070 13744 20076 13796
rect 20128 13784 20134 13796
rect 20625 13787 20683 13793
rect 20625 13784 20637 13787
rect 20128 13756 20637 13784
rect 20128 13744 20134 13756
rect 20625 13753 20637 13756
rect 20671 13753 20683 13787
rect 20625 13747 20683 13753
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22373 13787 22431 13793
rect 22373 13784 22385 13787
rect 22152 13756 22385 13784
rect 22152 13744 22158 13756
rect 22373 13753 22385 13756
rect 22419 13753 22431 13787
rect 22373 13747 22431 13753
rect 22465 13787 22523 13793
rect 22465 13753 22477 13787
rect 22511 13784 22523 13787
rect 22738 13784 22744 13796
rect 22511 13756 22744 13784
rect 22511 13753 22523 13756
rect 22465 13747 22523 13753
rect 22738 13744 22744 13756
rect 22796 13744 22802 13796
rect 24780 13784 24808 13824
rect 25038 13812 25044 13824
rect 25096 13812 25102 13864
rect 24949 13787 25007 13793
rect 24949 13784 24961 13787
rect 24780 13756 24961 13784
rect 24949 13753 24961 13756
rect 24995 13753 25007 13787
rect 24949 13747 25007 13753
rect 10686 13716 10692 13728
rect 10599 13688 10692 13716
rect 10686 13676 10692 13688
rect 10744 13716 10750 13728
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 10744 13688 11161 13716
rect 10744 13676 10750 13688
rect 11149 13685 11161 13688
rect 11195 13685 11207 13719
rect 12618 13716 12624 13728
rect 12579 13688 12624 13716
rect 11149 13679 11207 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 13998 13716 14004 13728
rect 13959 13688 14004 13716
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 17129 13719 17187 13725
rect 17129 13685 17141 13719
rect 17175 13716 17187 13719
rect 17586 13716 17592 13728
rect 17175 13688 17592 13716
rect 17175 13685 17187 13688
rect 17129 13679 17187 13685
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 18966 13676 18972 13728
rect 19024 13716 19030 13728
rect 19429 13719 19487 13725
rect 19429 13716 19441 13719
rect 19024 13688 19441 13716
rect 19024 13676 19030 13688
rect 19429 13685 19441 13688
rect 19475 13685 19487 13719
rect 19429 13679 19487 13685
rect 20717 13719 20775 13725
rect 20717 13685 20729 13719
rect 20763 13716 20775 13719
rect 20806 13716 20812 13728
rect 20763 13688 20812 13716
rect 20763 13685 20775 13688
rect 20717 13679 20775 13685
rect 20806 13676 20812 13688
rect 20864 13676 20870 13728
rect 22005 13719 22063 13725
rect 22005 13685 22017 13719
rect 22051 13716 22063 13719
rect 22554 13716 22560 13728
rect 22051 13688 22560 13716
rect 22051 13685 22063 13688
rect 22005 13679 22063 13685
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 10042 13512 10048 13524
rect 10003 13484 10048 13512
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10686 13512 10692 13524
rect 10183 13484 10692 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 11940 13484 12541 13512
rect 11940 13472 11946 13484
rect 12529 13481 12541 13484
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 13173 13515 13231 13521
rect 13173 13481 13185 13515
rect 13219 13512 13231 13515
rect 13998 13512 14004 13524
rect 13219 13484 14004 13512
rect 13219 13481 13231 13484
rect 13173 13475 13231 13481
rect 11416 13447 11474 13453
rect 11416 13413 11428 13447
rect 11462 13444 11474 13447
rect 11790 13444 11796 13456
rect 11462 13416 11796 13444
rect 11462 13413 11474 13416
rect 11416 13407 11474 13413
rect 11790 13404 11796 13416
rect 11848 13444 11854 13456
rect 12342 13444 12348 13456
rect 11848 13416 12348 13444
rect 11848 13404 11854 13416
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 13188 13444 13216 13475
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 15473 13515 15531 13521
rect 15473 13481 15485 13515
rect 15519 13512 15531 13515
rect 16482 13512 16488 13524
rect 15519 13484 16488 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 16577 13515 16635 13521
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 16758 13512 16764 13524
rect 16623 13484 16764 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 18322 13512 18328 13524
rect 16908 13484 16953 13512
rect 18283 13484 18328 13512
rect 16908 13472 16914 13484
rect 18322 13472 18328 13484
rect 18380 13512 18386 13524
rect 18690 13512 18696 13524
rect 18380 13484 18696 13512
rect 18380 13472 18386 13484
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 20717 13515 20775 13521
rect 20717 13481 20729 13515
rect 20763 13512 20775 13515
rect 20990 13512 20996 13524
rect 20763 13484 20996 13512
rect 20763 13481 20775 13484
rect 20717 13475 20775 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21634 13512 21640 13524
rect 21595 13484 21640 13512
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 23290 13512 23296 13524
rect 23251 13484 23296 13512
rect 23290 13472 23296 13484
rect 23348 13472 23354 13524
rect 12492 13416 13216 13444
rect 12492 13404 12498 13416
rect 13262 13404 13268 13456
rect 13320 13444 13326 13456
rect 14550 13444 14556 13456
rect 13320 13416 14556 13444
rect 13320 13404 13326 13416
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 15841 13447 15899 13453
rect 15841 13413 15853 13447
rect 15887 13444 15899 13447
rect 16022 13444 16028 13456
rect 15887 13416 16028 13444
rect 15887 13413 15899 13416
rect 15841 13407 15899 13413
rect 16022 13404 16028 13416
rect 16080 13444 16086 13456
rect 16206 13444 16212 13456
rect 16080 13416 16212 13444
rect 16080 13404 16086 13416
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 17034 13444 17040 13456
rect 16995 13416 17040 13444
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 18966 13404 18972 13456
rect 19024 13444 19030 13456
rect 19122 13447 19180 13453
rect 19122 13444 19134 13447
rect 19024 13416 19134 13444
rect 19024 13404 19030 13416
rect 19122 13413 19134 13416
rect 19168 13413 19180 13447
rect 19122 13407 19180 13413
rect 24026 13404 24032 13456
rect 24084 13453 24090 13456
rect 24084 13447 24148 13453
rect 24084 13413 24102 13447
rect 24136 13413 24148 13447
rect 24084 13407 24148 13413
rect 24084 13404 24090 13407
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 13998 13376 14004 13388
rect 12676 13348 14004 13376
rect 12676 13336 12682 13348
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 14093 13379 14151 13385
rect 14093 13345 14105 13379
rect 14139 13376 14151 13379
rect 15102 13376 15108 13388
rect 14139 13348 15108 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 11112 13280 11161 13308
rect 11112 13268 11118 13280
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 14108 13308 14136 13339
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 16942 13376 16948 13388
rect 15948 13348 16948 13376
rect 14274 13308 14280 13320
rect 13587 13280 14136 13308
rect 14235 13280 14280 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 15948 13317 15976 13348
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 18874 13376 18880 13388
rect 18835 13348 18880 13376
rect 18874 13336 18880 13348
rect 18932 13336 18938 13388
rect 20898 13376 20904 13388
rect 20859 13348 20904 13376
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 22554 13336 22560 13388
rect 22612 13376 22618 13388
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 22612 13348 22661 13376
rect 22612 13336 22618 13348
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 22649 13339 22707 13345
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15028 13280 15945 13308
rect 13630 13240 13636 13252
rect 13591 13212 13636 13240
rect 13630 13200 13636 13212
rect 13688 13200 13694 13252
rect 14734 13240 14740 13252
rect 14695 13212 14740 13240
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 11146 13172 11152 13184
rect 10919 13144 11152 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 15028 13181 15056 13280
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 16025 13311 16083 13317
rect 16025 13277 16037 13311
rect 16071 13308 16083 13311
rect 16574 13308 16580 13320
rect 16071 13280 16580 13308
rect 16071 13277 16083 13280
rect 16025 13271 16083 13277
rect 15378 13200 15384 13252
rect 15436 13240 15442 13252
rect 16040 13240 16068 13271
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 20772 13280 21097 13308
rect 20772 13268 20778 13280
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22741 13311 22799 13317
rect 22741 13308 22753 13311
rect 21968 13280 22753 13308
rect 21968 13268 21974 13280
rect 22741 13277 22753 13280
rect 22787 13277 22799 13311
rect 22922 13308 22928 13320
rect 22883 13280 22928 13308
rect 22741 13271 22799 13277
rect 22922 13268 22928 13280
rect 22980 13268 22986 13320
rect 23566 13268 23572 13320
rect 23624 13308 23630 13320
rect 23845 13311 23903 13317
rect 23845 13308 23857 13311
rect 23624 13280 23857 13308
rect 23624 13268 23630 13280
rect 15436 13212 16068 13240
rect 15436 13200 15442 13212
rect 20806 13200 20812 13252
rect 20864 13240 20870 13252
rect 22646 13240 22652 13252
rect 20864 13212 22652 13240
rect 20864 13200 20870 13212
rect 22646 13200 22652 13212
rect 22704 13200 22710 13252
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 12124 13144 15025 13172
rect 12124 13132 12130 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15013 13135 15071 13141
rect 18322 13132 18328 13184
rect 18380 13172 18386 13184
rect 19150 13172 19156 13184
rect 18380 13144 19156 13172
rect 18380 13132 18386 13144
rect 19150 13132 19156 13144
rect 19208 13132 19214 13184
rect 20162 13132 20168 13184
rect 20220 13172 20226 13184
rect 20257 13175 20315 13181
rect 20257 13172 20269 13175
rect 20220 13144 20269 13172
rect 20220 13132 20226 13144
rect 20257 13141 20269 13144
rect 20303 13141 20315 13175
rect 20257 13135 20315 13141
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22278 13172 22284 13184
rect 22152 13144 22197 13172
rect 22239 13144 22284 13172
rect 22152 13132 22158 13144
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 23382 13132 23388 13184
rect 23440 13172 23446 13184
rect 23676 13181 23704 13280
rect 23845 13277 23857 13280
rect 23891 13277 23903 13311
rect 23845 13271 23903 13277
rect 23661 13175 23719 13181
rect 23661 13172 23673 13175
rect 23440 13144 23673 13172
rect 23440 13132 23446 13144
rect 23661 13141 23673 13144
rect 23707 13141 23719 13175
rect 25222 13172 25228 13184
rect 25183 13144 25228 13172
rect 23661 13135 23719 13141
rect 25222 13132 25228 13144
rect 25280 13132 25286 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13998 12928 14004 12980
rect 14056 12968 14062 12980
rect 14093 12971 14151 12977
rect 14093 12968 14105 12971
rect 14056 12940 14105 12968
rect 14056 12928 14062 12940
rect 14093 12937 14105 12940
rect 14139 12937 14151 12971
rect 14093 12931 14151 12937
rect 14274 12928 14280 12980
rect 14332 12968 14338 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 14332 12940 16037 12968
rect 14332 12928 14338 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 16025 12931 16083 12937
rect 17037 12971 17095 12977
rect 17037 12937 17049 12971
rect 17083 12968 17095 12971
rect 17862 12968 17868 12980
rect 17083 12940 17868 12968
rect 17083 12937 17095 12940
rect 17037 12931 17095 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19024 12940 19441 12968
rect 19024 12928 19030 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 20530 12968 20536 12980
rect 19429 12931 19487 12937
rect 19904 12940 20536 12968
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 11425 12835 11483 12841
rect 11425 12832 11437 12835
rect 10367 12804 11437 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 11425 12801 11437 12804
rect 11471 12832 11483 12835
rect 11808 12832 11836 12928
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 11940 12872 12173 12900
rect 11940 12860 11946 12872
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 12161 12863 12219 12869
rect 18325 12903 18383 12909
rect 18325 12869 18337 12903
rect 18371 12900 18383 12903
rect 19334 12900 19340 12912
rect 18371 12872 19340 12900
rect 18371 12869 18383 12872
rect 18325 12863 18383 12869
rect 11471 12804 11836 12832
rect 12176 12832 12204 12863
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 19702 12900 19708 12912
rect 19663 12872 19708 12900
rect 19702 12860 19708 12872
rect 19760 12860 19766 12912
rect 16761 12835 16819 12841
rect 12176 12804 12572 12832
rect 11471 12801 11483 12804
rect 11425 12795 11483 12801
rect 12434 12764 12440 12776
rect 12395 12736 12440 12764
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12544 12764 12572 12804
rect 16761 12801 16773 12835
rect 16807 12832 16819 12835
rect 17494 12832 17500 12844
rect 16807 12804 17500 12832
rect 16807 12801 16819 12804
rect 16761 12795 16819 12801
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 17586 12792 17592 12844
rect 17644 12832 17650 12844
rect 18782 12832 18788 12844
rect 17644 12804 17689 12832
rect 18743 12804 18788 12832
rect 17644 12792 17650 12804
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 12693 12767 12751 12773
rect 12693 12764 12705 12767
rect 12544 12736 12705 12764
rect 12693 12733 12705 12736
rect 12739 12733 12751 12767
rect 12693 12727 12751 12733
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 13136 12736 14657 12764
rect 13136 12724 13142 12736
rect 14645 12733 14657 12736
rect 14691 12764 14703 12767
rect 14734 12764 14740 12776
rect 14691 12736 14740 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 16850 12724 16856 12776
rect 16908 12764 16914 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 16908 12736 17417 12764
rect 16908 12724 16914 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 18892 12764 18920 12795
rect 18966 12792 18972 12844
rect 19024 12832 19030 12844
rect 19904 12841 19932 12940
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 22922 12968 22928 12980
rect 22835 12940 22928 12968
rect 22922 12928 22928 12940
rect 22980 12968 22986 12980
rect 23477 12971 23535 12977
rect 23477 12968 23489 12971
rect 22980 12940 23489 12968
rect 22980 12928 22986 12940
rect 23477 12937 23489 12940
rect 23523 12968 23535 12971
rect 24026 12968 24032 12980
rect 23523 12940 24032 12968
rect 23523 12937 23535 12940
rect 23477 12931 23535 12937
rect 24026 12928 24032 12940
rect 24084 12968 24090 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 24084 12940 25053 12968
rect 24084 12928 24090 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 25041 12931 25099 12937
rect 23658 12860 23664 12912
rect 23716 12860 23722 12912
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 19024 12804 19901 12832
rect 19024 12792 19030 12804
rect 19889 12801 19901 12804
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 22373 12835 22431 12841
rect 22373 12801 22385 12835
rect 22419 12832 22431 12835
rect 23106 12832 23112 12844
rect 22419 12804 23112 12832
rect 22419 12801 22431 12804
rect 22373 12795 22431 12801
rect 23106 12792 23112 12804
rect 23164 12792 23170 12844
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 23676 12832 23704 12860
rect 23532 12804 23704 12832
rect 23532 12792 23538 12804
rect 18892 12736 19104 12764
rect 17405 12727 17463 12733
rect 10689 12699 10747 12705
rect 10689 12665 10701 12699
rect 10735 12696 10747 12699
rect 11149 12699 11207 12705
rect 11149 12696 11161 12699
rect 10735 12668 11161 12696
rect 10735 12665 10747 12668
rect 10689 12659 10747 12665
rect 11149 12665 11161 12668
rect 11195 12696 11207 12699
rect 11974 12696 11980 12708
rect 11195 12668 11980 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 11974 12656 11980 12668
rect 12032 12656 12038 12708
rect 14553 12699 14611 12705
rect 14553 12665 14565 12699
rect 14599 12696 14611 12699
rect 14826 12696 14832 12708
rect 14599 12668 14832 12696
rect 14599 12665 14611 12668
rect 14553 12659 14611 12665
rect 14826 12656 14832 12668
rect 14884 12705 14890 12708
rect 14884 12699 14948 12705
rect 14884 12665 14902 12699
rect 14936 12665 14948 12699
rect 14884 12659 14948 12665
rect 16669 12699 16727 12705
rect 16669 12665 16681 12699
rect 16715 12696 16727 12699
rect 17497 12699 17555 12705
rect 17497 12696 17509 12699
rect 16715 12668 17509 12696
rect 16715 12665 16727 12668
rect 16669 12659 16727 12665
rect 17497 12665 17509 12668
rect 17543 12696 17555 12699
rect 17678 12696 17684 12708
rect 17543 12668 17684 12696
rect 17543 12665 17555 12668
rect 17497 12659 17555 12665
rect 14884 12656 14890 12659
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 18693 12699 18751 12705
rect 18693 12665 18705 12699
rect 18739 12696 18751 12699
rect 18874 12696 18880 12708
rect 18739 12668 18880 12696
rect 18739 12665 18751 12668
rect 18693 12659 18751 12665
rect 18874 12656 18880 12668
rect 18932 12656 18938 12708
rect 11238 12628 11244 12640
rect 11199 12600 11244 12628
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 14734 12628 14740 12640
rect 13863 12600 14740 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 14734 12588 14740 12600
rect 14792 12588 14798 12640
rect 19076 12628 19104 12736
rect 19702 12724 19708 12776
rect 19760 12764 19766 12776
rect 20162 12773 20168 12776
rect 20145 12767 20168 12773
rect 20145 12764 20157 12767
rect 19760 12736 20157 12764
rect 19760 12724 19766 12736
rect 20145 12733 20157 12736
rect 20220 12764 20226 12776
rect 21542 12764 21548 12776
rect 20220 12736 20293 12764
rect 21503 12736 21548 12764
rect 20145 12727 20168 12733
rect 20162 12724 20168 12727
rect 20220 12724 20226 12736
rect 21542 12724 21548 12736
rect 21600 12724 21606 12776
rect 22097 12767 22155 12773
rect 22097 12733 22109 12767
rect 22143 12764 22155 12767
rect 22278 12764 22284 12776
rect 22143 12736 22284 12764
rect 22143 12733 22155 12736
rect 22097 12727 22155 12733
rect 22278 12724 22284 12736
rect 22336 12764 22342 12776
rect 22922 12764 22928 12776
rect 22336 12736 22928 12764
rect 22336 12724 22342 12736
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 23661 12767 23719 12773
rect 23661 12764 23673 12767
rect 23440 12736 23673 12764
rect 23440 12724 23446 12736
rect 23661 12733 23673 12736
rect 23707 12764 23719 12767
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 23707 12736 25329 12764
rect 23707 12733 23719 12736
rect 23661 12727 23719 12733
rect 25317 12733 25329 12736
rect 25363 12764 25375 12767
rect 25685 12767 25743 12773
rect 25685 12764 25697 12767
rect 25363 12736 25697 12764
rect 25363 12733 25375 12736
rect 25317 12727 25375 12733
rect 25685 12733 25697 12736
rect 25731 12733 25743 12767
rect 25685 12727 25743 12733
rect 20714 12656 20720 12708
rect 20772 12696 20778 12708
rect 21910 12696 21916 12708
rect 20772 12668 21916 12696
rect 20772 12656 20778 12668
rect 21910 12656 21916 12668
rect 21968 12656 21974 12708
rect 23750 12656 23756 12708
rect 23808 12696 23814 12708
rect 23906 12699 23964 12705
rect 23906 12696 23918 12699
rect 23808 12668 23918 12696
rect 23808 12656 23814 12668
rect 23906 12665 23918 12668
rect 23952 12665 23964 12699
rect 23906 12659 23964 12665
rect 19426 12628 19432 12640
rect 19076 12600 19432 12628
rect 19426 12588 19432 12600
rect 19484 12628 19490 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 19484 12600 21281 12628
rect 19484 12588 19490 12600
rect 21269 12597 21281 12600
rect 21315 12628 21327 12631
rect 21450 12628 21456 12640
rect 21315 12600 21456 12628
rect 21315 12597 21327 12600
rect 21269 12591 21327 12597
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 22370 12588 22376 12640
rect 22428 12628 22434 12640
rect 23566 12628 23572 12640
rect 22428 12600 23572 12628
rect 22428 12588 22434 12600
rect 23566 12588 23572 12600
rect 23624 12588 23630 12640
rect 24210 12588 24216 12640
rect 24268 12628 24274 12640
rect 24670 12628 24676 12640
rect 24268 12600 24676 12628
rect 24268 12588 24274 12600
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10505 12427 10563 12433
rect 10505 12424 10517 12427
rect 10192 12396 10517 12424
rect 10192 12384 10198 12396
rect 10505 12393 10517 12396
rect 10551 12393 10563 12427
rect 10505 12387 10563 12393
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11517 12427 11575 12433
rect 11517 12424 11529 12427
rect 11112 12396 11529 12424
rect 11112 12384 11118 12396
rect 11517 12393 11529 12396
rect 11563 12393 11575 12427
rect 11517 12387 11575 12393
rect 12069 12427 12127 12433
rect 12069 12393 12081 12427
rect 12115 12424 12127 12427
rect 12342 12424 12348 12436
rect 12115 12396 12348 12424
rect 12115 12393 12127 12396
rect 12069 12387 12127 12393
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 12584 12396 13645 12424
rect 12584 12384 12590 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 15102 12424 15108 12436
rect 13872 12396 15108 12424
rect 13872 12384 13878 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 16761 12427 16819 12433
rect 15804 12396 15976 12424
rect 15804 12384 15810 12396
rect 10873 12359 10931 12365
rect 10873 12325 10885 12359
rect 10919 12356 10931 12359
rect 10962 12356 10968 12368
rect 10919 12328 10968 12356
rect 10919 12325 10931 12328
rect 10873 12319 10931 12325
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 14737 12359 14795 12365
rect 14737 12356 14749 12359
rect 13096 12328 14749 12356
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 12308 12260 12449 12288
rect 12308 12248 12314 12260
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12189 11023 12223
rect 11146 12220 11152 12232
rect 11107 12192 11152 12220
rect 10965 12183 11023 12189
rect 10980 12152 11008 12183
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 12158 12180 12164 12232
rect 12216 12220 12222 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12216 12192 12541 12220
rect 12216 12180 12222 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12710 12220 12716 12232
rect 12623 12192 12716 12220
rect 12529 12183 12587 12189
rect 12710 12180 12716 12192
rect 12768 12220 12774 12232
rect 13096 12220 13124 12328
rect 14737 12325 14749 12328
rect 14783 12356 14795 12359
rect 15378 12356 15384 12368
rect 14783 12328 15384 12356
rect 14783 12325 14795 12328
rect 14737 12319 14795 12325
rect 15378 12316 15384 12328
rect 15436 12316 15442 12368
rect 15948 12356 15976 12396
rect 16761 12393 16773 12427
rect 16807 12424 16819 12427
rect 17034 12424 17040 12436
rect 16807 12396 17040 12424
rect 16807 12393 16819 12396
rect 16761 12387 16819 12393
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 19208 12396 19257 12424
rect 19208 12384 19214 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 20533 12427 20591 12433
rect 20533 12393 20545 12427
rect 20579 12424 20591 12427
rect 21082 12424 21088 12436
rect 20579 12396 21088 12424
rect 20579 12393 20591 12396
rect 20533 12387 20591 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 22554 12424 22560 12436
rect 22515 12396 22560 12424
rect 22554 12384 22560 12396
rect 22612 12384 22618 12436
rect 22922 12424 22928 12436
rect 22883 12396 22928 12424
rect 22922 12384 22928 12396
rect 22980 12384 22986 12436
rect 25590 12424 25596 12436
rect 25551 12396 25596 12424
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 17862 12356 17868 12368
rect 15488 12328 15884 12356
rect 15948 12328 17868 12356
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12288 13231 12291
rect 13998 12288 14004 12300
rect 13219 12260 14004 12288
rect 13219 12257 13231 12260
rect 13173 12251 13231 12257
rect 13998 12248 14004 12260
rect 14056 12248 14062 12300
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14148 12260 14872 12288
rect 14148 12248 14154 12260
rect 14274 12220 14280 12232
rect 12768 12192 13124 12220
rect 14235 12192 14280 12220
rect 12768 12180 12774 12192
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 11054 12152 11060 12164
rect 10980 12124 11060 12152
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 13446 12112 13452 12164
rect 13504 12152 13510 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 13504 12124 13553 12152
rect 13504 12112 13510 12124
rect 13541 12121 13553 12124
rect 13587 12152 13599 12155
rect 14292 12152 14320 12180
rect 13587 12124 14320 12152
rect 14844 12152 14872 12260
rect 14918 12248 14924 12300
rect 14976 12288 14982 12300
rect 15488 12288 15516 12328
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14976 12260 15516 12288
rect 15580 12260 15669 12288
rect 14976 12248 14982 12260
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15580 12220 15608 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15746 12220 15752 12232
rect 15344 12192 15608 12220
rect 15707 12192 15752 12220
rect 15344 12180 15350 12192
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15856 12229 15884 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 17954 12316 17960 12368
rect 18012 12356 18018 12368
rect 18598 12356 18604 12368
rect 18012 12328 18604 12356
rect 18012 12316 18018 12328
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 18874 12356 18880 12368
rect 18835 12328 18880 12356
rect 18874 12316 18880 12328
rect 18932 12316 18938 12368
rect 22186 12316 22192 12368
rect 22244 12356 22250 12368
rect 23290 12356 23296 12368
rect 22244 12328 23296 12356
rect 22244 12316 22250 12328
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 24480 12359 24538 12365
rect 24480 12325 24492 12359
rect 24526 12356 24538 12359
rect 24854 12356 24860 12368
rect 24526 12328 24860 12356
rect 24526 12325 24538 12328
rect 24480 12319 24538 12325
rect 24854 12316 24860 12328
rect 24912 12356 24918 12368
rect 25222 12356 25228 12368
rect 24912 12328 25228 12356
rect 24912 12316 24918 12328
rect 25222 12316 25228 12328
rect 25280 12316 25286 12368
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 16816 12260 17233 12288
rect 16816 12248 16822 12260
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 18782 12288 18788 12300
rect 18739 12260 18788 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 18782 12248 18788 12260
rect 18840 12248 18846 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19392 12260 19625 12288
rect 19392 12248 19398 12260
rect 19613 12257 19625 12260
rect 19659 12288 19671 12291
rect 20254 12288 20260 12300
rect 19659 12260 20260 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 21168 12291 21226 12297
rect 21168 12257 21180 12291
rect 21214 12288 21226 12291
rect 21450 12288 21456 12300
rect 21214 12260 21456 12288
rect 21214 12257 21226 12260
rect 21168 12251 21226 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 23106 12288 23112 12300
rect 23067 12260 23112 12288
rect 23106 12248 23112 12260
rect 23164 12248 23170 12300
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17313 12223 17371 12229
rect 17313 12220 17325 12223
rect 17184 12192 17325 12220
rect 17184 12180 17190 12192
rect 17313 12189 17325 12192
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 16853 12155 16911 12161
rect 16853 12152 16865 12155
rect 14844 12124 16865 12152
rect 13587 12121 13599 12124
rect 13541 12115 13599 12121
rect 16853 12121 16865 12124
rect 16899 12121 16911 12155
rect 17420 12152 17448 12183
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 19208 12192 19717 12220
rect 19208 12180 19214 12192
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 19886 12220 19892 12232
rect 19847 12192 19892 12220
rect 19705 12183 19763 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 20530 12180 20536 12232
rect 20588 12220 20594 12232
rect 20901 12223 20959 12229
rect 20901 12220 20913 12223
rect 20588 12192 20913 12220
rect 20588 12180 20594 12192
rect 20901 12189 20913 12192
rect 20947 12189 20959 12223
rect 20901 12183 20959 12189
rect 23382 12180 23388 12232
rect 23440 12220 23446 12232
rect 24029 12223 24087 12229
rect 24029 12220 24041 12223
rect 23440 12192 24041 12220
rect 23440 12180 23446 12192
rect 24029 12189 24041 12192
rect 24075 12220 24087 12223
rect 24213 12223 24271 12229
rect 24213 12220 24225 12223
rect 24075 12192 24225 12220
rect 24075 12189 24087 12192
rect 24029 12183 24087 12189
rect 24213 12189 24225 12192
rect 24259 12189 24271 12223
rect 24213 12183 24271 12189
rect 18138 12152 18144 12164
rect 16853 12115 16911 12121
rect 17328 12124 17448 12152
rect 18051 12124 18144 12152
rect 11977 12087 12035 12093
rect 11977 12053 11989 12087
rect 12023 12084 12035 12087
rect 12434 12084 12440 12096
rect 12023 12056 12440 12084
rect 12023 12053 12035 12056
rect 11977 12047 12035 12053
rect 12434 12044 12440 12056
rect 12492 12084 12498 12096
rect 13078 12084 13084 12096
rect 12492 12056 13084 12084
rect 12492 12044 12498 12056
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 14274 12044 14280 12096
rect 14332 12084 14338 12096
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 14332 12056 15025 12084
rect 14332 12044 14338 12056
rect 15013 12053 15025 12056
rect 15059 12084 15071 12087
rect 15746 12084 15752 12096
rect 15059 12056 15752 12084
rect 15059 12053 15071 12056
rect 15013 12047 15071 12053
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 16080 12056 16313 12084
rect 16080 12044 16086 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16301 12047 16359 12053
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 17328 12084 17356 12124
rect 18138 12112 18144 12124
rect 18196 12152 18202 12164
rect 18782 12152 18788 12164
rect 18196 12124 18788 12152
rect 18196 12112 18202 12124
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 23474 12112 23480 12164
rect 23532 12152 23538 12164
rect 24118 12152 24124 12164
rect 23532 12124 24124 12152
rect 23532 12112 23538 12124
rect 24118 12112 24124 12124
rect 24176 12112 24182 12164
rect 16632 12056 17356 12084
rect 16632 12044 16638 12056
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18417 12087 18475 12093
rect 18417 12084 18429 12087
rect 18288 12056 18429 12084
rect 18288 12044 18294 12056
rect 18417 12053 18429 12056
rect 18463 12084 18475 12087
rect 18693 12087 18751 12093
rect 18693 12084 18705 12087
rect 18463 12056 18705 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 18693 12053 18705 12056
rect 18739 12053 18751 12087
rect 18693 12047 18751 12053
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 22244 12056 22293 12084
rect 22244 12044 22250 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 23750 12084 23756 12096
rect 23711 12056 23756 12084
rect 22281 12047 22339 12053
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 10597 11883 10655 11889
rect 10597 11849 10609 11883
rect 10643 11880 10655 11883
rect 10962 11880 10968 11892
rect 10643 11852 10968 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12710 11880 12716 11892
rect 12299 11852 12716 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 13357 11883 13415 11889
rect 13357 11849 13369 11883
rect 13403 11880 13415 11883
rect 13446 11880 13452 11892
rect 13403 11852 13452 11880
rect 13403 11849 13415 11852
rect 13357 11843 13415 11849
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 16025 11883 16083 11889
rect 16025 11880 16037 11883
rect 14056 11852 16037 11880
rect 14056 11840 14062 11852
rect 16025 11849 16037 11852
rect 16071 11849 16083 11883
rect 16025 11843 16083 11849
rect 19521 11883 19579 11889
rect 19521 11849 19533 11883
rect 19567 11880 19579 11883
rect 19886 11880 19892 11892
rect 19567 11852 19892 11880
rect 19567 11849 19579 11852
rect 19521 11843 19579 11849
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 20346 11880 20352 11892
rect 20307 11852 20352 11880
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 20622 11880 20628 11892
rect 20487 11852 20628 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 21450 11880 21456 11892
rect 21411 11852 21456 11880
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 22002 11880 22008 11892
rect 21963 11852 22008 11880
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 24854 11840 24860 11892
rect 24912 11840 24918 11892
rect 10873 11815 10931 11821
rect 10873 11781 10885 11815
rect 10919 11812 10931 11815
rect 11054 11812 11060 11824
rect 10919 11784 11060 11812
rect 10919 11781 10931 11784
rect 10873 11775 10931 11781
rect 11054 11772 11060 11784
rect 11112 11812 11118 11824
rect 11112 11784 13676 11812
rect 11112 11772 11118 11784
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11744 11851 11747
rect 12250 11744 12256 11756
rect 11839 11716 12256 11744
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 13354 11744 13360 11756
rect 12851 11716 13360 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13648 11744 13676 11784
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 15197 11815 15255 11821
rect 15197 11812 15209 11815
rect 14884 11784 15209 11812
rect 14884 11772 14890 11784
rect 15197 11781 15209 11784
rect 15243 11781 15255 11815
rect 15562 11812 15568 11824
rect 15523 11784 15568 11812
rect 15197 11775 15255 11781
rect 15562 11772 15568 11784
rect 15620 11772 15626 11824
rect 24872 11812 24900 11840
rect 22664 11784 24900 11812
rect 13648 11716 13952 11744
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11676 12587 11679
rect 12618 11676 12624 11688
rect 12575 11648 12624 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 13078 11636 13084 11688
rect 13136 11676 13142 11688
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 13136 11648 13829 11676
rect 13136 11636 13142 11648
rect 13817 11645 13829 11648
rect 13863 11645 13875 11679
rect 13924 11676 13952 11716
rect 15580 11676 15608 11772
rect 16574 11744 16580 11756
rect 16535 11716 16580 11744
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 17770 11744 17776 11756
rect 17731 11716 17776 11744
rect 17770 11704 17776 11716
rect 17828 11744 17834 11756
rect 18601 11747 18659 11753
rect 17828 11716 18460 11744
rect 17828 11704 17834 11716
rect 18432 11688 18460 11716
rect 18601 11713 18613 11747
rect 18647 11713 18659 11747
rect 21082 11744 21088 11756
rect 21043 11716 21088 11744
rect 18601 11707 18659 11713
rect 16393 11679 16451 11685
rect 16393 11676 16405 11679
rect 13924 11648 14228 11676
rect 15580 11648 16405 11676
rect 13817 11639 13875 11645
rect 11146 11568 11152 11620
rect 11204 11608 11210 11620
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 11204 11580 11345 11608
rect 11204 11568 11210 11580
rect 11333 11577 11345 11580
rect 11379 11608 11391 11611
rect 12253 11611 12311 11617
rect 12253 11608 12265 11611
rect 11379 11580 12265 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 12253 11577 12265 11580
rect 12299 11577 12311 11611
rect 14062 11611 14120 11617
rect 14062 11608 14074 11611
rect 12253 11571 12311 11577
rect 13740 11580 14074 11608
rect 13740 11552 13768 11580
rect 14062 11577 14074 11580
rect 14108 11577 14120 11611
rect 14200 11608 14228 11648
rect 16393 11645 16405 11648
rect 16439 11676 16451 11679
rect 16482 11676 16488 11688
rect 16439 11648 16488 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 18414 11676 18420 11688
rect 18327 11648 18420 11676
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 14200 11580 17172 11608
rect 14062 11571 14120 11577
rect 17144 11552 17172 11580
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 18616 11608 18644 11707
rect 21082 11704 21088 11716
rect 21140 11704 21146 11756
rect 22462 11704 22468 11756
rect 22520 11744 22526 11756
rect 22664 11753 22692 11784
rect 22649 11747 22707 11753
rect 22649 11744 22661 11747
rect 22520 11716 22661 11744
rect 22520 11704 22526 11716
rect 22649 11713 22661 11716
rect 22695 11713 22707 11747
rect 22649 11707 22707 11713
rect 24118 11704 24124 11756
rect 24176 11744 24182 11756
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 24176 11716 24225 11744
rect 24176 11704 24182 11716
rect 24213 11713 24225 11716
rect 24259 11744 24271 11747
rect 24762 11744 24768 11756
rect 24259 11716 24768 11744
rect 24259 11713 24271 11716
rect 24213 11707 24271 11713
rect 24762 11704 24768 11716
rect 24820 11704 24826 11756
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11713 24915 11747
rect 24857 11707 24915 11713
rect 20346 11636 20352 11688
rect 20404 11676 20410 11688
rect 20809 11679 20867 11685
rect 20809 11676 20821 11679
rect 20404 11648 20821 11676
rect 20404 11636 20410 11648
rect 20809 11645 20821 11648
rect 20855 11645 20867 11679
rect 20809 11639 20867 11645
rect 21913 11679 21971 11685
rect 21913 11645 21925 11679
rect 21959 11676 21971 11679
rect 22922 11676 22928 11688
rect 21959 11648 22928 11676
rect 21959 11645 21971 11648
rect 21913 11639 21971 11645
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 23477 11679 23535 11685
rect 23477 11645 23489 11679
rect 23523 11676 23535 11679
rect 23842 11676 23848 11688
rect 23523 11648 23848 11676
rect 23523 11645 23535 11648
rect 23477 11639 23535 11645
rect 23842 11636 23848 11648
rect 23900 11676 23906 11688
rect 24872 11676 24900 11707
rect 23900 11648 24900 11676
rect 23900 11636 23906 11648
rect 19061 11611 19119 11617
rect 19061 11608 19073 11611
rect 18380 11580 19073 11608
rect 18380 11568 18386 11580
rect 19061 11577 19073 11580
rect 19107 11577 19119 11611
rect 20898 11608 20904 11620
rect 20859 11580 20904 11608
rect 19061 11571 19119 11577
rect 20898 11568 20904 11580
rect 20956 11608 20962 11620
rect 23017 11611 23075 11617
rect 23017 11608 23029 11611
rect 20956 11580 23029 11608
rect 20956 11568 20962 11580
rect 23017 11577 23029 11580
rect 23063 11577 23075 11611
rect 23017 11571 23075 11577
rect 23382 11568 23388 11620
rect 23440 11608 23446 11620
rect 25317 11611 25375 11617
rect 25317 11608 25329 11611
rect 23440 11580 25329 11608
rect 23440 11568 23446 11580
rect 25317 11577 25329 11580
rect 25363 11608 25375 11611
rect 25685 11611 25743 11617
rect 25685 11608 25697 11611
rect 25363 11580 25697 11608
rect 25363 11577 25375 11580
rect 25317 11571 25375 11577
rect 25685 11577 25697 11580
rect 25731 11577 25743 11611
rect 25685 11571 25743 11577
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 13354 11540 13360 11552
rect 11664 11512 13360 11540
rect 11664 11500 11670 11512
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13722 11540 13728 11552
rect 13683 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 15933 11543 15991 11549
rect 15933 11509 15945 11543
rect 15979 11540 15991 11543
rect 16298 11540 16304 11552
rect 15979 11512 16304 11540
rect 15979 11509 15991 11512
rect 15933 11503 15991 11509
rect 16298 11500 16304 11512
rect 16356 11540 16362 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 16356 11512 16497 11540
rect 16356 11500 16362 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16485 11503 16543 11509
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 17037 11543 17095 11549
rect 17037 11540 17049 11543
rect 16816 11512 17049 11540
rect 16816 11500 16822 11512
rect 17037 11509 17049 11512
rect 17083 11509 17095 11543
rect 17037 11503 17095 11509
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 17184 11512 17417 11540
rect 17184 11500 17190 11512
rect 17405 11509 17417 11512
rect 17451 11509 17463 11543
rect 17405 11503 17463 11509
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17920 11512 18061 11540
rect 17920 11500 17926 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11540 18567 11543
rect 18782 11540 18788 11552
rect 18555 11512 18788 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19889 11543 19947 11549
rect 19889 11509 19901 11543
rect 19935 11540 19947 11543
rect 19978 11540 19984 11552
rect 19935 11512 19984 11540
rect 19935 11509 19947 11512
rect 19889 11503 19947 11509
rect 19978 11500 19984 11512
rect 20036 11540 20042 11552
rect 20806 11540 20812 11552
rect 20036 11512 20812 11540
rect 20036 11500 20042 11512
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 22373 11543 22431 11549
rect 22373 11540 22385 11543
rect 22336 11512 22385 11540
rect 22336 11500 22342 11512
rect 22373 11509 22385 11512
rect 22419 11509 22431 11543
rect 22373 11503 22431 11509
rect 22465 11543 22523 11549
rect 22465 11509 22477 11543
rect 22511 11540 22523 11543
rect 22922 11540 22928 11552
rect 22511 11512 22928 11540
rect 22511 11509 22523 11512
rect 22465 11503 22523 11509
rect 22922 11500 22928 11512
rect 22980 11500 22986 11552
rect 24210 11500 24216 11552
rect 24268 11540 24274 11552
rect 24305 11543 24363 11549
rect 24305 11540 24317 11543
rect 24268 11512 24317 11540
rect 24268 11500 24274 11512
rect 24305 11509 24317 11512
rect 24351 11509 24363 11543
rect 24305 11503 24363 11509
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 24673 11543 24731 11549
rect 24673 11540 24685 11543
rect 24636 11512 24685 11540
rect 24636 11500 24642 11512
rect 24673 11509 24685 11512
rect 24719 11509 24731 11543
rect 24673 11503 24731 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12710 11336 12716 11348
rect 12207 11308 12716 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 14090 11336 14096 11348
rect 13495 11308 14096 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14737 11339 14795 11345
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 14826 11336 14832 11348
rect 14783 11308 14832 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15378 11336 15384 11348
rect 15335 11308 15384 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 19150 11336 19156 11348
rect 19111 11308 19156 11336
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19613 11339 19671 11345
rect 19300 11308 19345 11336
rect 19300 11296 19306 11308
rect 19613 11305 19625 11339
rect 19659 11336 19671 11339
rect 20070 11336 20076 11348
rect 19659 11308 20076 11336
rect 19659 11305 19671 11308
rect 19613 11299 19671 11305
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20714 11336 20720 11348
rect 20675 11308 20720 11336
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20864 11308 21005 11336
rect 20864 11296 20870 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 21358 11336 21364 11348
rect 21319 11308 21364 11336
rect 20993 11299 21051 11305
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 22097 11339 22155 11345
rect 22097 11305 22109 11339
rect 22143 11336 22155 11339
rect 22278 11336 22284 11348
rect 22143 11308 22284 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22462 11336 22468 11348
rect 22423 11308 22468 11336
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 23750 11296 23756 11348
rect 23808 11336 23814 11348
rect 24121 11339 24179 11345
rect 24121 11336 24133 11339
rect 23808 11308 24133 11336
rect 23808 11296 23814 11308
rect 24121 11305 24133 11308
rect 24167 11305 24179 11339
rect 24854 11336 24860 11348
rect 24815 11308 24860 11336
rect 24121 11299 24179 11305
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25133 11339 25191 11345
rect 25133 11305 25145 11339
rect 25179 11336 25191 11339
rect 25866 11336 25872 11348
rect 25179 11308 25872 11336
rect 25179 11305 25191 11308
rect 25133 11299 25191 11305
rect 25866 11296 25872 11308
rect 25924 11296 25930 11348
rect 13998 11228 14004 11280
rect 14056 11268 14062 11280
rect 14844 11268 14872 11296
rect 16301 11271 16359 11277
rect 16301 11268 16313 11271
rect 14056 11240 14780 11268
rect 14844 11240 16313 11268
rect 14056 11228 14062 11240
rect 13814 11160 13820 11212
rect 13872 11160 13878 11212
rect 13909 11203 13967 11209
rect 13909 11169 13921 11203
rect 13955 11200 13967 11203
rect 14642 11200 14648 11212
rect 13955 11172 14648 11200
rect 13955 11169 13967 11172
rect 13909 11163 13967 11169
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 14752 11200 14780 11240
rect 16301 11237 16313 11240
rect 16347 11268 16359 11271
rect 16574 11268 16580 11280
rect 16347 11240 16580 11268
rect 16347 11237 16359 11240
rect 16301 11231 16359 11237
rect 16574 11228 16580 11240
rect 16632 11268 16638 11280
rect 16669 11271 16727 11277
rect 16669 11268 16681 11271
rect 16632 11240 16681 11268
rect 16632 11228 16638 11240
rect 16669 11237 16681 11240
rect 16715 11237 16727 11271
rect 20732 11268 20760 11296
rect 20732 11240 21496 11268
rect 16669 11231 16727 11237
rect 14826 11200 14832 11212
rect 14752 11172 14832 11200
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 15470 11160 15476 11212
rect 15528 11200 15534 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15528 11172 15669 11200
rect 15528 11160 15534 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11200 17555 11203
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 17543 11172 17969 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 17957 11169 17969 11172
rect 18003 11200 18015 11203
rect 19242 11200 19248 11212
rect 18003 11172 19248 11200
rect 18003 11169 18015 11172
rect 17957 11163 18015 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 19705 11203 19763 11209
rect 19705 11169 19717 11203
rect 19751 11200 19763 11203
rect 19978 11200 19984 11212
rect 19751 11172 19984 11200
rect 19751 11169 19763 11172
rect 19705 11163 19763 11169
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 21468 11200 21496 11240
rect 22738 11228 22744 11280
rect 22796 11268 22802 11280
rect 22986 11271 23044 11277
rect 22986 11268 22998 11271
rect 22796 11240 22998 11268
rect 22796 11228 22802 11240
rect 22986 11237 22998 11240
rect 23032 11237 23044 11271
rect 22986 11231 23044 11237
rect 23106 11228 23112 11280
rect 23164 11268 23170 11280
rect 23382 11268 23388 11280
rect 23164 11240 23388 11268
rect 23164 11228 23170 11240
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 23124 11200 23152 11228
rect 21468 11172 21588 11200
rect 13832 11132 13860 11160
rect 13998 11132 14004 11144
rect 13832 11104 14004 11132
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 14185 11135 14243 11141
rect 14185 11101 14197 11135
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 12618 11064 12624 11076
rect 12579 11036 12624 11064
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 13814 11064 13820 11076
rect 13587 11036 13820 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 13081 10999 13139 11005
rect 13081 10965 13093 10999
rect 13127 10996 13139 10999
rect 13262 10996 13268 11008
rect 13127 10968 13268 10996
rect 13127 10965 13139 10968
rect 13081 10959 13139 10965
rect 13262 10956 13268 10968
rect 13320 10996 13326 11008
rect 14200 10996 14228 11095
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15344 11104 15761 11132
rect 15344 11092 15350 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15930 11132 15936 11144
rect 15891 11104 15936 11132
rect 15749 11095 15807 11101
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 19886 11132 19892 11144
rect 18279 11104 19380 11132
rect 19847 11104 19892 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 15010 11064 15016 11076
rect 14971 11036 15016 11064
rect 15010 11024 15016 11036
rect 15068 11024 15074 11076
rect 17589 11067 17647 11073
rect 17589 11033 17601 11067
rect 17635 11064 17647 11067
rect 17862 11064 17868 11076
rect 17635 11036 17868 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 14458 10996 14464 11008
rect 13320 10968 14464 10996
rect 13320 10956 13326 10968
rect 14458 10956 14464 10968
rect 14516 10996 14522 11008
rect 15930 10996 15936 11008
rect 14516 10968 15936 10996
rect 14516 10956 14522 10968
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17129 10999 17187 11005
rect 17129 10996 17141 10999
rect 17000 10968 17141 10996
rect 17000 10956 17006 10968
rect 17129 10965 17141 10968
rect 17175 10996 17187 10999
rect 18046 10996 18052 11008
rect 17175 10968 18052 10996
rect 17175 10965 17187 10968
rect 17129 10959 17187 10965
rect 18046 10956 18052 10968
rect 18104 10996 18110 11008
rect 18248 10996 18276 11095
rect 18104 10968 18276 10996
rect 18104 10956 18110 10968
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 18601 10999 18659 11005
rect 18601 10996 18613 10999
rect 18380 10968 18613 10996
rect 18380 10956 18386 10968
rect 18601 10965 18613 10968
rect 18647 10965 18659 10999
rect 19352 10996 19380 11104
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21560 11141 21588 11172
rect 22756 11172 23152 11200
rect 22756 11141 22784 11172
rect 23290 11160 23296 11212
rect 23348 11200 23354 11212
rect 24949 11203 25007 11209
rect 24949 11200 24961 11203
rect 23348 11172 24961 11200
rect 23348 11160 23354 11172
rect 24949 11169 24961 11172
rect 24995 11200 25007 11203
rect 25774 11200 25780 11212
rect 24995 11172 25780 11200
rect 24995 11169 25007 11172
rect 24949 11163 25007 11169
rect 25774 11160 25780 11172
rect 25832 11160 25838 11212
rect 21453 11135 21511 11141
rect 21453 11132 21465 11135
rect 20772 11104 21465 11132
rect 20772 11092 20778 11104
rect 21453 11101 21465 11104
rect 21499 11101 21511 11135
rect 21453 11095 21511 11101
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11101 21603 11135
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 21545 11095 21603 11101
rect 22020 11104 22753 11132
rect 20530 11024 20536 11076
rect 20588 11064 20594 11076
rect 22020 11064 22048 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 20588 11036 22048 11064
rect 24489 11067 24547 11073
rect 20588 11024 20594 11036
rect 24489 11033 24501 11067
rect 24535 11064 24547 11067
rect 24578 11064 24584 11076
rect 24535 11036 24584 11064
rect 24535 11033 24547 11036
rect 24489 11027 24547 11033
rect 24578 11024 24584 11036
rect 24636 11064 24642 11076
rect 24636 11036 24900 11064
rect 24636 11024 24642 11036
rect 19426 10996 19432 11008
rect 19352 10968 19432 10996
rect 18601 10959 18659 10965
rect 19426 10956 19432 10968
rect 19484 10956 19490 11008
rect 24872 10996 24900 11036
rect 25314 10996 25320 11008
rect 24872 10968 25320 10996
rect 25314 10956 25320 10968
rect 25372 10956 25378 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 14642 10792 14648 10804
rect 14603 10764 14648 10792
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 15749 10795 15807 10801
rect 15749 10761 15761 10795
rect 15795 10792 15807 10795
rect 15930 10792 15936 10804
rect 15795 10764 15936 10792
rect 15795 10761 15807 10764
rect 15749 10755 15807 10761
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 17586 10792 17592 10804
rect 17547 10764 17592 10792
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18414 10792 18420 10804
rect 18288 10764 18420 10792
rect 18288 10752 18294 10764
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 19426 10792 19432 10804
rect 19387 10764 19432 10792
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 19797 10795 19855 10801
rect 19797 10761 19809 10795
rect 19843 10792 19855 10795
rect 20070 10792 20076 10804
rect 19843 10764 20076 10792
rect 19843 10761 19855 10764
rect 19797 10755 19855 10761
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 20165 10795 20223 10801
rect 20165 10761 20177 10795
rect 20211 10792 20223 10795
rect 20714 10792 20720 10804
rect 20211 10764 20720 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 21358 10792 21364 10804
rect 21131 10764 21364 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 21726 10752 21732 10804
rect 21784 10792 21790 10804
rect 23385 10795 23443 10801
rect 23385 10792 23397 10795
rect 21784 10764 23397 10792
rect 21784 10752 21790 10764
rect 23385 10761 23397 10764
rect 23431 10761 23443 10795
rect 25774 10792 25780 10804
rect 25735 10764 25780 10792
rect 23385 10755 23443 10761
rect 14660 10656 14688 10752
rect 22738 10724 22744 10736
rect 22699 10696 22744 10724
rect 22738 10684 22744 10696
rect 22796 10684 22802 10736
rect 15197 10659 15255 10665
rect 15197 10656 15209 10659
rect 14660 10628 15209 10656
rect 15197 10625 15209 10628
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 16942 10656 16948 10668
rect 16347 10628 16948 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 19518 10616 19524 10668
rect 19576 10656 19582 10668
rect 20257 10659 20315 10665
rect 20257 10656 20269 10659
rect 19576 10628 20269 10656
rect 19576 10616 19582 10628
rect 20257 10625 20269 10628
rect 20303 10625 20315 10659
rect 23400 10656 23428 10755
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 24302 10656 24308 10668
rect 23400 10628 24308 10656
rect 20257 10619 20315 10625
rect 24302 10616 24308 10628
rect 24360 10616 24366 10668
rect 25314 10656 25320 10668
rect 25275 10628 25320 10656
rect 25314 10616 25320 10628
rect 25372 10616 25378 10668
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 13078 10588 13084 10600
rect 13035 10560 13084 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12710 10520 12716 10532
rect 12299 10492 12716 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12710 10480 12716 10492
rect 12768 10520 12774 10532
rect 13004 10520 13032 10551
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 13262 10597 13268 10600
rect 13256 10588 13268 10597
rect 13223 10560 13268 10588
rect 13256 10551 13268 10560
rect 13262 10548 13268 10551
rect 13320 10548 13326 10600
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14366 10588 14372 10600
rect 14240 10560 14372 10588
rect 14240 10548 14246 10560
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 16761 10591 16819 10597
rect 16761 10557 16773 10591
rect 16807 10588 16819 10591
rect 17034 10588 17040 10600
rect 16807 10560 17040 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 17034 10548 17040 10560
rect 17092 10588 17098 10600
rect 17770 10588 17776 10600
rect 17092 10560 17776 10588
rect 17092 10548 17098 10560
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 18012 10560 18061 10588
rect 18012 10548 18018 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 20530 10548 20536 10600
rect 20588 10588 20594 10600
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 20588 10560 21373 10588
rect 20588 10548 20594 10560
rect 21361 10557 21373 10560
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 21628 10591 21686 10597
rect 21628 10557 21640 10591
rect 21674 10588 21686 10591
rect 22186 10588 22192 10600
rect 21674 10560 22192 10588
rect 21674 10557 21686 10560
rect 21628 10551 21686 10557
rect 22186 10548 22192 10560
rect 22244 10588 22250 10600
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22244 10560 23029 10588
rect 22244 10548 22250 10560
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 24121 10591 24179 10597
rect 24121 10557 24133 10591
rect 24167 10588 24179 10591
rect 24210 10588 24216 10600
rect 24167 10560 24216 10588
rect 24167 10557 24179 10560
rect 24121 10551 24179 10557
rect 24210 10548 24216 10560
rect 24268 10588 24274 10600
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24268 10560 25145 10588
rect 24268 10548 24274 10560
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 12768 10492 13032 10520
rect 12768 10480 12774 10492
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 18322 10529 18328 10532
rect 18316 10520 18328 10529
rect 13780 10492 14412 10520
rect 18283 10492 18328 10520
rect 13780 10480 13786 10492
rect 14384 10464 14412 10492
rect 18316 10483 18328 10492
rect 18322 10480 18328 10483
rect 18380 10480 18386 10532
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12584 10424 12817 10452
rect 12584 10412 12590 10424
rect 12805 10421 12817 10424
rect 12851 10452 12863 10455
rect 13998 10452 14004 10464
rect 12851 10424 14004 10452
rect 12851 10421 12863 10424
rect 12805 10415 12863 10421
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14366 10452 14372 10464
rect 14327 10424 14372 10452
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 15010 10452 15016 10464
rect 14971 10424 15016 10452
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 16390 10452 16396 10464
rect 16351 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16850 10412 16856 10464
rect 16908 10452 16914 10464
rect 23753 10455 23811 10461
rect 16908 10424 16953 10452
rect 16908 10412 16914 10424
rect 23753 10421 23765 10455
rect 23799 10452 23811 10455
rect 24026 10452 24032 10464
rect 23799 10424 24032 10452
rect 23799 10421 23811 10424
rect 23753 10415 23811 10421
rect 24026 10412 24032 10424
rect 24084 10412 24090 10464
rect 24210 10412 24216 10464
rect 24268 10452 24274 10464
rect 24765 10455 24823 10461
rect 24765 10452 24777 10455
rect 24268 10424 24777 10452
rect 24268 10412 24274 10424
rect 24765 10421 24777 10424
rect 24811 10421 24823 10455
rect 26142 10452 26148 10464
rect 26103 10424 26148 10452
rect 24765 10415 24823 10421
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 12621 10251 12679 10257
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 13722 10248 13728 10260
rect 12667 10220 13728 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14093 10251 14151 10257
rect 14093 10217 14105 10251
rect 14139 10248 14151 10251
rect 14458 10248 14464 10260
rect 14139 10220 14464 10248
rect 14139 10217 14151 10220
rect 14093 10211 14151 10217
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 15611 10220 16681 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 16669 10217 16681 10220
rect 16715 10248 16727 10251
rect 16850 10248 16856 10260
rect 16715 10220 16856 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 17034 10248 17040 10260
rect 16995 10220 17040 10248
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18012 10220 18797 10248
rect 18012 10208 18018 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 19334 10248 19340 10260
rect 19295 10220 19340 10248
rect 18785 10211 18843 10217
rect 12894 10180 12900 10192
rect 11992 10152 12900 10180
rect 11238 10072 11244 10124
rect 11296 10112 11302 10124
rect 11514 10112 11520 10124
rect 11296 10084 11520 10112
rect 11296 10072 11302 10084
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 11609 10115 11667 10121
rect 11609 10081 11621 10115
rect 11655 10112 11667 10115
rect 11882 10112 11888 10124
rect 11655 10084 11888 10112
rect 11655 10081 11667 10084
rect 11609 10075 11667 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11756 10016 11805 10044
rect 11756 10004 11762 10016
rect 11793 10013 11805 10016
rect 11839 10044 11851 10047
rect 11992 10044 12020 10152
rect 12894 10140 12900 10152
rect 12952 10189 12958 10192
rect 12952 10183 13016 10189
rect 12952 10149 12970 10183
rect 13004 10149 13016 10183
rect 12952 10143 13016 10149
rect 12952 10140 12958 10143
rect 13354 10140 13360 10192
rect 13412 10180 13418 10192
rect 13412 10152 16896 10180
rect 13412 10140 13418 10152
rect 16868 10124 16896 10152
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 17374 10183 17432 10189
rect 17374 10180 17386 10183
rect 17000 10152 17386 10180
rect 17000 10140 17006 10152
rect 17374 10149 17386 10152
rect 17420 10149 17432 10183
rect 17374 10143 17432 10149
rect 12710 10112 12716 10124
rect 12623 10084 12716 10112
rect 12710 10072 12716 10084
rect 12768 10112 12774 10124
rect 12768 10084 15332 10112
rect 12768 10072 12774 10084
rect 11839 10016 12020 10044
rect 11839 10013 11851 10016
rect 11793 10007 11851 10013
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14734 10044 14740 10056
rect 14516 10016 14740 10044
rect 14516 10004 14522 10016
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15304 9988 15332 10084
rect 15746 10072 15752 10124
rect 15804 10112 15810 10124
rect 15933 10115 15991 10121
rect 15933 10112 15945 10115
rect 15804 10084 15945 10112
rect 15804 10072 15810 10084
rect 15933 10081 15945 10084
rect 15979 10081 15991 10115
rect 15933 10075 15991 10081
rect 16850 10072 16856 10124
rect 16908 10072 16914 10124
rect 18800 10112 18828 10211
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 21361 10251 21419 10257
rect 21361 10248 21373 10251
rect 20364 10220 21373 10248
rect 20364 10192 20392 10220
rect 21361 10217 21373 10220
rect 21407 10248 21419 10251
rect 21818 10248 21824 10260
rect 21407 10220 21824 10248
rect 21407 10217 21419 10220
rect 21361 10211 21419 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 22741 10251 22799 10257
rect 22741 10248 22753 10251
rect 22152 10220 22753 10248
rect 22152 10208 22158 10220
rect 22741 10217 22753 10220
rect 22787 10217 22799 10251
rect 22741 10211 22799 10217
rect 23106 10208 23112 10260
rect 23164 10248 23170 10260
rect 23569 10251 23627 10257
rect 23569 10248 23581 10251
rect 23164 10220 23581 10248
rect 23164 10208 23170 10220
rect 23569 10217 23581 10220
rect 23615 10217 23627 10251
rect 23569 10211 23627 10217
rect 19242 10180 19248 10192
rect 19203 10152 19248 10180
rect 19242 10140 19248 10152
rect 19300 10140 19306 10192
rect 20346 10180 20352 10192
rect 20307 10152 20352 10180
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 22281 10183 22339 10189
rect 22281 10180 22293 10183
rect 21008 10152 22293 10180
rect 21008 10124 21036 10152
rect 22281 10149 22293 10152
rect 22327 10149 22339 10183
rect 22281 10143 22339 10149
rect 19610 10112 19616 10124
rect 18800 10084 19616 10112
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10112 20775 10115
rect 20990 10112 20996 10124
rect 20763 10084 20996 10112
rect 20763 10081 20775 10084
rect 20717 10075 20775 10081
rect 20990 10072 20996 10084
rect 21048 10072 21054 10124
rect 21266 10112 21272 10124
rect 21227 10084 21272 10112
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 22738 10072 22744 10124
rect 22796 10112 22802 10124
rect 23201 10115 23259 10121
rect 23201 10112 23213 10115
rect 22796 10084 23213 10112
rect 22796 10072 22802 10084
rect 23201 10081 23213 10084
rect 23247 10081 23259 10115
rect 23584 10112 23612 10211
rect 24302 10208 24308 10260
rect 24360 10248 24366 10260
rect 25133 10251 25191 10257
rect 25133 10248 25145 10251
rect 24360 10220 25145 10248
rect 24360 10208 24366 10220
rect 25133 10217 25145 10220
rect 25179 10217 25191 10251
rect 25133 10211 25191 10217
rect 23842 10140 23848 10192
rect 23900 10180 23906 10192
rect 23998 10183 24056 10189
rect 23998 10180 24010 10183
rect 23900 10152 24010 10180
rect 23900 10140 23906 10152
rect 23998 10149 24010 10152
rect 24044 10149 24056 10183
rect 23998 10143 24056 10149
rect 23753 10115 23811 10121
rect 23753 10112 23765 10115
rect 23584 10084 23765 10112
rect 23201 10075 23259 10081
rect 23753 10081 23765 10084
rect 23799 10112 23811 10115
rect 25409 10115 25467 10121
rect 25409 10112 25421 10115
rect 23799 10084 25421 10112
rect 23799 10081 23811 10084
rect 23753 10075 23811 10081
rect 25409 10081 25421 10084
rect 25455 10112 25467 10115
rect 26142 10112 26148 10124
rect 25455 10084 26148 10112
rect 25455 10081 25467 10084
rect 25409 10075 25467 10081
rect 26142 10072 26148 10084
rect 26200 10072 26206 10124
rect 16022 10044 16028 10056
rect 15983 10016 16028 10044
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 16206 10044 16212 10056
rect 16167 10016 16212 10044
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16724 10016 17141 10044
rect 16724 10004 16730 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21591 10016 21956 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 15286 9936 15292 9988
rect 15344 9976 15350 9988
rect 16684 9976 16712 10004
rect 15344 9948 16712 9976
rect 15344 9936 15350 9948
rect 21928 9920 21956 10016
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 10962 9908 10968 9920
rect 10919 9880 10968 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11149 9911 11207 9917
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 11195 9880 15025 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 15013 9877 15025 9880
rect 15059 9908 15071 9911
rect 15470 9908 15476 9920
rect 15059 9880 15476 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 18506 9908 18512 9920
rect 18467 9880 18512 9908
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 19886 9908 19892 9920
rect 19847 9880 19892 9908
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20530 9908 20536 9920
rect 20491 9880 20536 9908
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 20898 9908 20904 9920
rect 20859 9880 20904 9908
rect 20898 9868 20904 9880
rect 20956 9868 20962 9920
rect 21910 9908 21916 9920
rect 21871 9880 21916 9908
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 11698 9704 11704 9716
rect 11440 9676 11704 9704
rect 10778 9636 10784 9648
rect 10739 9608 10784 9636
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 11440 9577 11468 9676
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 11882 9704 11888 9716
rect 11843 9676 11888 9704
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 12250 9704 12256 9716
rect 12163 9676 12256 9704
rect 12250 9664 12256 9676
rect 12308 9704 12314 9716
rect 12710 9704 12716 9716
rect 12308 9676 12716 9704
rect 12308 9664 12314 9676
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 14277 9707 14335 9713
rect 14277 9673 14289 9707
rect 14323 9704 14335 9707
rect 14366 9704 14372 9716
rect 14323 9676 14372 9704
rect 14323 9673 14335 9676
rect 14277 9667 14335 9673
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 15013 9707 15071 9713
rect 15013 9673 15025 9707
rect 15059 9704 15071 9707
rect 15286 9704 15292 9716
rect 15059 9676 15292 9704
rect 15059 9673 15071 9676
rect 15013 9667 15071 9673
rect 12618 9596 12624 9648
rect 12676 9636 12682 9648
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 12676 9608 13461 9636
rect 12676 9596 12682 9608
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 13449 9599 13507 9605
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 15028 9636 15056 9667
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 18230 9704 18236 9716
rect 16264 9676 16620 9704
rect 16264 9664 16270 9676
rect 16482 9636 16488 9648
rect 14700 9608 15056 9636
rect 15948 9608 16488 9636
rect 14700 9596 14706 9608
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 9999 9540 10333 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10321 9537 10333 9540
rect 10367 9568 10379 9571
rect 11425 9571 11483 9577
rect 11425 9568 11437 9571
rect 10367 9540 11437 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 11425 9537 11437 9540
rect 11471 9537 11483 9571
rect 12894 9568 12900 9580
rect 12855 9540 12900 9568
rect 11425 9531 11483 9537
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9568 13415 9571
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13403 9540 14013 9568
rect 13403 9537 13415 9540
rect 13357 9531 13415 9537
rect 14001 9537 14013 9540
rect 14047 9568 14059 9571
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14047 9540 14289 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 15948 9577 15976 9608
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 16592 9636 16620 9676
rect 17880 9676 18236 9704
rect 17313 9639 17371 9645
rect 17313 9636 17325 9639
rect 16592 9608 17325 9636
rect 17313 9605 17325 9608
rect 17359 9636 17371 9639
rect 17880 9636 17908 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 19610 9664 19616 9716
rect 19668 9704 19674 9716
rect 20530 9704 20536 9716
rect 19668 9676 20536 9704
rect 19668 9664 19674 9676
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 21637 9707 21695 9713
rect 21637 9704 21649 9707
rect 21416 9676 21649 9704
rect 21416 9664 21422 9676
rect 21637 9673 21649 9676
rect 21683 9673 21695 9707
rect 21637 9667 21695 9673
rect 23845 9707 23903 9713
rect 23845 9673 23857 9707
rect 23891 9704 23903 9707
rect 24210 9704 24216 9716
rect 23891 9676 24216 9704
rect 23891 9673 23903 9676
rect 23845 9667 23903 9673
rect 17359 9608 17908 9636
rect 17359 9605 17371 9608
rect 17313 9599 17371 9605
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 21269 9639 21327 9645
rect 21269 9636 21281 9639
rect 20772 9608 21281 9636
rect 20772 9596 20778 9608
rect 21269 9605 21281 9608
rect 21315 9605 21327 9639
rect 21269 9599 21327 9605
rect 15933 9571 15991 9577
rect 14884 9540 15332 9568
rect 14884 9528 14890 9540
rect 13814 9500 13820 9512
rect 13775 9472 13820 9500
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 15102 9500 15108 9512
rect 13964 9472 15108 9500
rect 13964 9460 13970 9472
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9469 15255 9503
rect 15304 9500 15332 9540
rect 15933 9537 15945 9571
rect 15979 9537 15991 9571
rect 16114 9568 16120 9580
rect 16075 9540 16120 9568
rect 15933 9531 15991 9537
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 17862 9568 17868 9580
rect 17775 9540 17868 9568
rect 17862 9528 17868 9540
rect 17920 9568 17926 9580
rect 18506 9568 18512 9580
rect 17920 9540 18512 9568
rect 17920 9528 17926 9540
rect 18506 9528 18512 9540
rect 18564 9568 18570 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 18564 9540 18613 9568
rect 18564 9528 18570 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 19610 9568 19616 9580
rect 19571 9540 19616 9568
rect 18601 9531 18659 9537
rect 19610 9528 19616 9540
rect 19668 9528 19674 9580
rect 15304 9472 15976 9500
rect 15197 9463 15255 9469
rect 10689 9435 10747 9441
rect 10689 9401 10701 9435
rect 10735 9432 10747 9435
rect 15212 9432 15240 9463
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 10735 9404 11284 9432
rect 10735 9401 10747 9404
rect 10689 9395 10747 9401
rect 11146 9364 11152 9376
rect 11107 9336 11152 9364
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11256 9373 11284 9404
rect 14476 9404 15240 9432
rect 15396 9404 15853 9432
rect 11241 9367 11299 9373
rect 11241 9333 11253 9367
rect 11287 9364 11299 9367
rect 11698 9364 11704 9376
rect 11287 9336 11704 9364
rect 11287 9333 11299 9336
rect 11241 9327 11299 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 13722 9364 13728 9376
rect 12483 9336 13728 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 14476 9373 14504 9404
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14332 9336 14473 9364
rect 14332 9324 14338 9336
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 14461 9327 14519 9333
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14792 9336 14841 9364
rect 14792 9324 14798 9336
rect 14829 9333 14841 9336
rect 14875 9364 14887 9367
rect 15396 9364 15424 9404
rect 15841 9401 15853 9404
rect 15887 9401 15899 9435
rect 15948 9432 15976 9472
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16080 9472 16865 9500
rect 16080 9460 16086 9472
rect 16853 9469 16865 9472
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18417 9503 18475 9509
rect 18417 9500 18429 9503
rect 18012 9472 18429 9500
rect 18012 9460 18018 9472
rect 18417 9469 18429 9472
rect 18463 9500 18475 9503
rect 19061 9503 19119 9509
rect 19061 9500 19073 9503
rect 18463 9472 19073 9500
rect 18463 9469 18475 9472
rect 18417 9463 18475 9469
rect 19061 9469 19073 9472
rect 19107 9469 19119 9503
rect 19061 9463 19119 9469
rect 16206 9432 16212 9444
rect 15948 9404 16212 9432
rect 15841 9395 15899 9401
rect 16206 9392 16212 9404
rect 16264 9392 16270 9444
rect 18322 9392 18328 9444
rect 18380 9432 18386 9444
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 18380 9404 18521 9432
rect 18380 9392 18386 9404
rect 18509 9401 18521 9404
rect 18555 9401 18567 9435
rect 19518 9432 19524 9444
rect 19479 9404 19524 9432
rect 18509 9395 18567 9401
rect 19518 9392 19524 9404
rect 19576 9432 19582 9444
rect 19858 9435 19916 9441
rect 19858 9432 19870 9435
rect 19576 9404 19870 9432
rect 19576 9392 19582 9404
rect 19858 9401 19870 9404
rect 19904 9401 19916 9435
rect 21284 9432 21312 9599
rect 21652 9500 21680 9667
rect 24210 9664 24216 9676
rect 24268 9664 24274 9716
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 21968 9540 22385 9568
rect 21968 9528 21974 9540
rect 22373 9537 22385 9540
rect 22419 9537 22431 9571
rect 22373 9531 22431 9537
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 23900 9540 24501 9568
rect 23900 9528 23906 9540
rect 24489 9537 24501 9540
rect 24535 9568 24547 9571
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24535 9540 24869 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 24857 9537 24869 9540
rect 24903 9568 24915 9571
rect 25130 9568 25136 9580
rect 24903 9540 25136 9568
rect 24903 9537 24915 9540
rect 24857 9531 24915 9537
rect 25130 9528 25136 9540
rect 25188 9568 25194 9580
rect 25225 9571 25283 9577
rect 25225 9568 25237 9571
rect 25188 9540 25237 9568
rect 25188 9528 25194 9540
rect 25225 9537 25237 9540
rect 25271 9537 25283 9571
rect 25225 9531 25283 9537
rect 22189 9503 22247 9509
rect 22189 9500 22201 9503
rect 21652 9472 22201 9500
rect 22189 9469 22201 9472
rect 22235 9469 22247 9503
rect 22189 9463 22247 9469
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9500 22339 9503
rect 23382 9500 23388 9512
rect 22327 9472 23388 9500
rect 22327 9469 22339 9472
rect 22281 9463 22339 9469
rect 22296 9432 22324 9463
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 24305 9435 24363 9441
rect 24305 9432 24317 9435
rect 21284 9404 22324 9432
rect 23032 9404 24317 9432
rect 19858 9395 19916 9401
rect 23032 9376 23060 9404
rect 24305 9401 24317 9404
rect 24351 9401 24363 9435
rect 24305 9395 24363 9401
rect 14875 9336 15424 9364
rect 15473 9367 15531 9373
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 15473 9333 15485 9367
rect 15519 9364 15531 9367
rect 15562 9364 15568 9376
rect 15519 9336 15568 9364
rect 15519 9333 15531 9336
rect 15473 9327 15531 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18049 9367 18107 9373
rect 18049 9364 18061 9367
rect 18012 9336 18061 9364
rect 18012 9324 18018 9336
rect 18049 9333 18061 9336
rect 18095 9333 18107 9367
rect 18049 9327 18107 9333
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 20993 9367 21051 9373
rect 20993 9364 21005 9367
rect 20864 9336 21005 9364
rect 20864 9324 20870 9336
rect 20993 9333 21005 9336
rect 21039 9333 21051 9367
rect 21818 9364 21824 9376
rect 21779 9336 21824 9364
rect 20993 9327 21051 9333
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 23014 9364 23020 9376
rect 22975 9336 23020 9364
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 23474 9364 23480 9376
rect 23387 9336 23480 9364
rect 23474 9324 23480 9336
rect 23532 9364 23538 9376
rect 24210 9364 24216 9376
rect 23532 9336 24216 9364
rect 23532 9324 23538 9336
rect 24210 9324 24216 9336
rect 24268 9324 24274 9376
rect 25406 9364 25412 9376
rect 25367 9336 25412 9364
rect 25406 9324 25412 9336
rect 25464 9324 25470 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 12952 9132 13185 9160
rect 12952 9120 12958 9132
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13814 9160 13820 9172
rect 13775 9132 13820 9160
rect 13173 9123 13231 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 15105 9163 15163 9169
rect 15105 9129 15117 9163
rect 15151 9160 15163 9163
rect 16114 9160 16120 9172
rect 15151 9132 16120 9160
rect 15151 9129 15163 9132
rect 15105 9123 15163 9129
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 16356 9132 17233 9160
rect 16356 9120 16362 9132
rect 17221 9129 17233 9132
rect 17267 9160 17279 9163
rect 17310 9160 17316 9172
rect 17267 9132 17316 9160
rect 17267 9129 17279 9132
rect 17221 9123 17279 9129
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 17957 9163 18015 9169
rect 17957 9129 17969 9163
rect 18003 9160 18015 9163
rect 18046 9160 18052 9172
rect 18003 9132 18052 9160
rect 18003 9129 18015 9132
rect 17957 9123 18015 9129
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 18322 9160 18328 9172
rect 18283 9132 18328 9160
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 20717 9163 20775 9169
rect 20717 9160 20729 9163
rect 20404 9132 20729 9160
rect 20404 9120 20410 9132
rect 20717 9129 20729 9132
rect 20763 9160 20775 9163
rect 21266 9160 21272 9172
rect 20763 9132 21272 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 21266 9120 21272 9132
rect 21324 9120 21330 9172
rect 23017 9163 23075 9169
rect 23017 9129 23029 9163
rect 23063 9160 23075 9163
rect 23106 9160 23112 9172
rect 23063 9132 23112 9160
rect 23063 9129 23075 9132
rect 23017 9123 23075 9129
rect 23106 9120 23112 9132
rect 23164 9160 23170 9172
rect 23477 9163 23535 9169
rect 23477 9160 23489 9163
rect 23164 9132 23489 9160
rect 23164 9120 23170 9132
rect 23477 9129 23489 9132
rect 23523 9160 23535 9163
rect 23569 9163 23627 9169
rect 23569 9160 23581 9163
rect 23523 9132 23581 9160
rect 23523 9129 23535 9132
rect 23477 9123 23535 9129
rect 23569 9129 23581 9132
rect 23615 9129 23627 9163
rect 25130 9160 25136 9172
rect 25091 9132 25136 9160
rect 23569 9123 23627 9129
rect 25130 9120 25136 9132
rect 25188 9120 25194 9172
rect 10781 9095 10839 9101
rect 10781 9061 10793 9095
rect 10827 9092 10839 9095
rect 10870 9092 10876 9104
rect 10827 9064 10876 9092
rect 10827 9061 10839 9064
rect 10781 9055 10839 9061
rect 10870 9052 10876 9064
rect 10928 9052 10934 9104
rect 11701 9095 11759 9101
rect 11701 9061 11713 9095
rect 11747 9092 11759 9095
rect 12250 9092 12256 9104
rect 11747 9064 12256 9092
rect 11747 9061 11759 9064
rect 11701 9055 11759 9061
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10686 9024 10692 9036
rect 10551 8996 10692 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 11808 9033 11836 9064
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 13541 9095 13599 9101
rect 13541 9061 13553 9095
rect 13587 9092 13599 9095
rect 13906 9092 13912 9104
rect 13587 9064 13912 9092
rect 13587 9061 13599 9064
rect 13541 9055 13599 9061
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 14737 9095 14795 9101
rect 14737 9061 14749 9095
rect 14783 9092 14795 9095
rect 18785 9095 18843 9101
rect 14783 9064 15792 9092
rect 14783 9061 14795 9064
rect 14737 9055 14795 9061
rect 12066 9033 12072 9036
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 10796 8996 11805 9024
rect 10796 8968 10824 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 12060 8987 12072 9033
rect 12124 9024 12130 9036
rect 12124 8996 12160 9024
rect 12066 8984 12072 8987
rect 12124 8984 12130 8996
rect 13630 8984 13636 9036
rect 13688 9024 13694 9036
rect 13814 9024 13820 9036
rect 13688 8996 13820 9024
rect 13688 8984 13694 8996
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 15654 9024 15660 9036
rect 15615 8996 15660 9024
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 15764 9033 15792 9064
rect 18785 9061 18797 9095
rect 18831 9092 18843 9095
rect 19613 9095 19671 9101
rect 19613 9092 19625 9095
rect 18831 9064 19625 9092
rect 18831 9061 18843 9064
rect 18785 9055 18843 9061
rect 19613 9061 19625 9064
rect 19659 9092 19671 9095
rect 19978 9092 19984 9104
rect 19659 9064 19984 9092
rect 19659 9061 19671 9064
rect 19613 9055 19671 9061
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 9024 15807 9027
rect 16482 9024 16488 9036
rect 15795 8996 16488 9024
rect 15795 8993 15807 8996
rect 15749 8987 15807 8993
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 20530 9024 20536 9036
rect 19751 8996 20536 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 10778 8916 10784 8968
rect 10836 8916 10842 8968
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8956 14243 8959
rect 14826 8956 14832 8968
rect 14231 8928 14832 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 15930 8956 15936 8968
rect 15891 8928 15936 8956
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16758 8916 16764 8968
rect 16816 8956 16822 8968
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 16816 8928 17325 8956
rect 16816 8916 16822 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 17494 8956 17500 8968
rect 17455 8928 17500 8956
rect 17313 8919 17371 8925
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 19153 8959 19211 8965
rect 19153 8925 19165 8959
rect 19199 8956 19211 8959
rect 19720 8956 19748 8987
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 20864 8996 20913 9024
rect 20864 8984 20870 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 21168 9027 21226 9033
rect 21168 8993 21180 9027
rect 21214 9024 21226 9027
rect 21726 9024 21732 9036
rect 21214 8996 21732 9024
rect 21214 8993 21226 8996
rect 21168 8987 21226 8993
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 23382 8984 23388 9036
rect 23440 9024 23446 9036
rect 24009 9027 24067 9033
rect 24009 9024 24021 9027
rect 23440 8996 24021 9024
rect 23440 8984 23446 8996
rect 24009 8993 24021 8996
rect 24055 8993 24067 9027
rect 24009 8987 24067 8993
rect 19199 8928 19748 8956
rect 19889 8959 19947 8965
rect 19199 8925 19211 8928
rect 19153 8919 19211 8925
rect 19889 8925 19901 8959
rect 19935 8925 19947 8959
rect 19889 8919 19947 8925
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8956 23535 8959
rect 23753 8959 23811 8965
rect 23753 8956 23765 8959
rect 23523 8928 23765 8956
rect 23523 8925 23535 8928
rect 23477 8919 23535 8925
rect 23753 8925 23765 8928
rect 23799 8925 23811 8959
rect 23753 8919 23811 8925
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 13630 8888 13636 8900
rect 12860 8860 13636 8888
rect 12860 8848 12866 8860
rect 13630 8848 13636 8860
rect 13688 8888 13694 8900
rect 15470 8888 15476 8900
rect 13688 8860 15476 8888
rect 13688 8848 13694 8860
rect 15470 8848 15476 8860
rect 15528 8848 15534 8900
rect 15654 8848 15660 8900
rect 15712 8888 15718 8900
rect 16853 8891 16911 8897
rect 16853 8888 16865 8891
rect 15712 8860 16865 8888
rect 15712 8848 15718 8860
rect 16853 8857 16865 8860
rect 16899 8857 16911 8891
rect 16853 8851 16911 8857
rect 19518 8848 19524 8900
rect 19576 8888 19582 8900
rect 19794 8888 19800 8900
rect 19576 8860 19800 8888
rect 19576 8848 19582 8860
rect 19794 8848 19800 8860
rect 19852 8888 19858 8900
rect 19904 8888 19932 8919
rect 19852 8860 20760 8888
rect 19852 8848 19858 8860
rect 11238 8820 11244 8832
rect 11199 8792 11244 8820
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 15286 8820 15292 8832
rect 15247 8792 15292 8820
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15746 8780 15752 8832
rect 15804 8820 15810 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 15804 8792 16405 8820
rect 15804 8780 15810 8792
rect 16393 8789 16405 8792
rect 16439 8820 16451 8823
rect 16482 8820 16488 8832
rect 16439 8792 16488 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 16666 8820 16672 8832
rect 16627 8792 16672 8820
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 18598 8780 18604 8832
rect 18656 8820 18662 8832
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 18656 8792 19257 8820
rect 18656 8780 18662 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 20254 8820 20260 8832
rect 20215 8792 20260 8820
rect 19245 8783 19303 8789
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 20732 8820 20760 8860
rect 22281 8823 22339 8829
rect 22281 8820 22293 8823
rect 20732 8792 22293 8820
rect 22281 8789 22293 8792
rect 22327 8789 22339 8823
rect 22646 8820 22652 8832
rect 22607 8792 22652 8820
rect 22281 8783 22339 8789
rect 22646 8780 22652 8792
rect 22704 8780 22710 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11563 8588 11897 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 11885 8585 11897 8588
rect 11931 8616 11943 8619
rect 12066 8616 12072 8628
rect 11931 8588 12072 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12066 8576 12072 8588
rect 12124 8616 12130 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12124 8588 12173 8616
rect 12124 8576 12130 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 15654 8616 15660 8628
rect 13863 8588 15660 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 12176 8480 12204 8579
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 17368 8588 17417 8616
rect 17368 8576 17374 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17405 8579 17463 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 19794 8616 19800 8628
rect 19755 8588 19800 8616
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 20349 8619 20407 8625
rect 20349 8585 20361 8619
rect 20395 8616 20407 8619
rect 20990 8616 20996 8628
rect 20395 8588 20996 8616
rect 20395 8585 20407 8588
rect 20349 8579 20407 8585
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 23934 8576 23940 8628
rect 23992 8616 23998 8628
rect 24213 8619 24271 8625
rect 24213 8616 24225 8619
rect 23992 8588 24225 8616
rect 23992 8576 23998 8588
rect 24213 8585 24225 8588
rect 24259 8616 24271 8619
rect 24259 8588 24808 8616
rect 24259 8585 24271 8588
rect 24213 8579 24271 8585
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 14274 8548 14280 8560
rect 12492 8520 12537 8548
rect 14235 8520 14280 8548
rect 12492 8508 12498 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12176 8452 13001 8480
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 17880 8480 17908 8576
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 22097 8551 22155 8557
rect 22097 8548 22109 8551
rect 21784 8520 22109 8548
rect 21784 8508 21790 8520
rect 22097 8517 22109 8520
rect 22143 8548 22155 8551
rect 22373 8551 22431 8557
rect 22373 8548 22385 8551
rect 22143 8520 22385 8548
rect 22143 8517 22155 8520
rect 22097 8511 22155 8517
rect 22373 8517 22385 8520
rect 22419 8517 22431 8551
rect 22373 8511 22431 8517
rect 24118 8508 24124 8560
rect 24176 8548 24182 8560
rect 24305 8551 24363 8557
rect 24305 8548 24317 8551
rect 24176 8520 24317 8548
rect 24176 8508 24182 8520
rect 24305 8517 24317 8520
rect 24351 8517 24363 8551
rect 24305 8511 24363 8517
rect 24780 8489 24808 8588
rect 24765 8483 24823 8489
rect 17880 8452 18184 8480
rect 12989 8443 13047 8449
rect 10134 8412 10140 8424
rect 10095 8384 10140 8412
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 13998 8372 14004 8424
rect 14056 8412 14062 8424
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 14056 8384 14473 8412
rect 14056 8372 14062 8384
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 14642 8412 14648 8424
rect 14599 8384 14648 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 14820 8415 14878 8421
rect 14820 8412 14832 8415
rect 14752 8384 14832 8412
rect 10045 8347 10103 8353
rect 10045 8313 10057 8347
rect 10091 8344 10103 8347
rect 10382 8347 10440 8353
rect 10382 8344 10394 8347
rect 10091 8316 10394 8344
rect 10091 8313 10103 8316
rect 10045 8307 10103 8313
rect 10382 8313 10394 8316
rect 10428 8344 10440 8347
rect 10962 8344 10968 8356
rect 10428 8316 10968 8344
rect 10428 8313 10440 8316
rect 10382 8307 10440 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 14185 8347 14243 8353
rect 14185 8313 14197 8347
rect 14231 8344 14243 8347
rect 14752 8344 14780 8384
rect 14820 8381 14832 8384
rect 14866 8412 14878 8415
rect 16114 8412 16120 8424
rect 14866 8384 16120 8412
rect 14866 8381 14878 8384
rect 14820 8375 14878 8381
rect 16114 8372 16120 8384
rect 16172 8412 16178 8424
rect 16485 8415 16543 8421
rect 16485 8412 16497 8415
rect 16172 8384 16497 8412
rect 16172 8372 16178 8384
rect 16485 8381 16497 8384
rect 16531 8412 16543 8415
rect 17494 8412 17500 8424
rect 16531 8384 17500 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18156 8412 18184 8452
rect 24765 8449 24777 8483
rect 24811 8449 24823 8483
rect 24765 8443 24823 8449
rect 24949 8483 25007 8489
rect 24949 8449 24961 8483
rect 24995 8480 25007 8483
rect 25038 8480 25044 8492
rect 24995 8452 25044 8480
rect 24995 8449 25007 8452
rect 24949 8443 25007 8449
rect 25038 8440 25044 8452
rect 25096 8480 25102 8492
rect 25317 8483 25375 8489
rect 25317 8480 25329 8483
rect 25096 8452 25329 8480
rect 25096 8440 25102 8452
rect 25317 8449 25329 8452
rect 25363 8449 25375 8483
rect 25317 8443 25375 8449
rect 18305 8415 18363 8421
rect 18305 8412 18317 8415
rect 18156 8384 18317 8412
rect 18305 8381 18317 8384
rect 18351 8381 18363 8415
rect 18305 8375 18363 8381
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8412 20591 8415
rect 20622 8412 20628 8424
rect 20579 8384 20628 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8412 20775 8415
rect 22646 8412 22652 8424
rect 20763 8384 22652 8412
rect 20763 8381 20775 8384
rect 20717 8375 20775 8381
rect 22646 8372 22652 8384
rect 22704 8412 22710 8424
rect 23198 8412 23204 8424
rect 22704 8384 23204 8412
rect 22704 8372 22710 8384
rect 23198 8372 23204 8384
rect 23256 8372 23262 8424
rect 23477 8415 23535 8421
rect 23477 8381 23489 8415
rect 23523 8412 23535 8415
rect 24673 8415 24731 8421
rect 24673 8412 24685 8415
rect 23523 8384 24685 8412
rect 23523 8381 23535 8384
rect 23477 8375 23535 8381
rect 24673 8381 24685 8384
rect 24719 8412 24731 8415
rect 25406 8412 25412 8424
rect 24719 8384 25412 8412
rect 24719 8381 24731 8384
rect 24673 8375 24731 8381
rect 25406 8372 25412 8384
rect 25464 8372 25470 8424
rect 16758 8344 16764 8356
rect 14231 8316 14780 8344
rect 16719 8316 16764 8344
rect 14231 8313 14243 8316
rect 14185 8307 14243 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 16942 8344 16948 8356
rect 16903 8316 16948 8344
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 20962 8347 21020 8353
rect 20962 8344 20974 8347
rect 20272 8316 20974 8344
rect 20272 8288 20300 8316
rect 20962 8313 20974 8316
rect 21008 8344 21020 8347
rect 21910 8344 21916 8356
rect 21008 8316 21916 8344
rect 21008 8313 21020 8316
rect 20962 8307 21020 8313
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 23109 8347 23167 8353
rect 23109 8313 23121 8347
rect 23155 8344 23167 8347
rect 23382 8344 23388 8356
rect 23155 8316 23388 8344
rect 23155 8313 23167 8316
rect 23109 8307 23167 8313
rect 23382 8304 23388 8316
rect 23440 8344 23446 8356
rect 24854 8344 24860 8356
rect 23440 8316 24860 8344
rect 23440 8304 23446 8316
rect 24854 8304 24860 8316
rect 24912 8304 24918 8356
rect 10870 8236 10876 8288
rect 10928 8276 10934 8288
rect 11330 8276 11336 8288
rect 10928 8248 11336 8276
rect 10928 8236 10934 8248
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 12802 8276 12808 8288
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 15930 8276 15936 8288
rect 12952 8248 12997 8276
rect 15891 8248 15936 8276
rect 12952 8236 12958 8248
rect 15930 8236 15936 8248
rect 15988 8236 15994 8288
rect 20254 8276 20260 8288
rect 20215 8248 20260 8276
rect 20254 8236 20260 8248
rect 20312 8236 20318 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 10686 8072 10692 8084
rect 10643 8044 10692 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 11112 8044 12173 8072
rect 11112 8032 11118 8044
rect 12161 8041 12173 8044
rect 12207 8072 12219 8075
rect 12250 8072 12256 8084
rect 12207 8044 12256 8072
rect 12207 8041 12219 8044
rect 12161 8035 12219 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12802 8072 12808 8084
rect 12763 8044 12808 8072
rect 12802 8032 12808 8044
rect 12860 8072 12866 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12860 8044 13001 8072
rect 12860 8032 12866 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 13998 8032 14004 8084
rect 14056 8072 14062 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 14056 8044 14289 8072
rect 14056 8032 14062 8044
rect 14277 8041 14289 8044
rect 14323 8041 14335 8075
rect 14277 8035 14335 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 14884 8044 15669 8072
rect 14884 8032 14890 8044
rect 15657 8041 15669 8044
rect 15703 8041 15715 8075
rect 15657 8035 15715 8041
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 16853 8075 16911 8081
rect 16853 8072 16865 8075
rect 16632 8044 16865 8072
rect 16632 8032 16638 8044
rect 16853 8041 16865 8044
rect 16899 8041 16911 8075
rect 16853 8035 16911 8041
rect 19245 8075 19303 8081
rect 19245 8041 19257 8075
rect 19291 8072 19303 8075
rect 21361 8075 21419 8081
rect 21361 8072 21373 8075
rect 19291 8044 21373 8072
rect 19291 8041 19303 8044
rect 19245 8035 19303 8041
rect 21361 8041 21373 8044
rect 21407 8072 21419 8075
rect 21913 8075 21971 8081
rect 21913 8072 21925 8075
rect 21407 8044 21925 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 21913 8041 21925 8044
rect 21959 8041 21971 8075
rect 22278 8072 22284 8084
rect 22239 8044 22284 8072
rect 21913 8035 21971 8041
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 24854 8032 24860 8084
rect 24912 8072 24918 8084
rect 25041 8075 25099 8081
rect 25041 8072 25053 8075
rect 24912 8044 25053 8072
rect 24912 8032 24918 8044
rect 25041 8041 25053 8044
rect 25087 8041 25099 8075
rect 25041 8035 25099 8041
rect 12529 8007 12587 8013
rect 12529 7973 12541 8007
rect 12575 8004 12587 8007
rect 12894 8004 12900 8016
rect 12575 7976 12900 8004
rect 12575 7973 12587 7976
rect 12529 7967 12587 7973
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 16666 8004 16672 8016
rect 16627 7976 16672 8004
rect 16666 7964 16672 7976
rect 16724 8004 16730 8016
rect 18046 8004 18052 8016
rect 16724 7976 18052 8004
rect 16724 7964 16730 7976
rect 18046 7964 18052 7976
rect 18104 7964 18110 8016
rect 18690 7964 18696 8016
rect 18748 8004 18754 8016
rect 19705 8007 19763 8013
rect 19705 8004 19717 8007
rect 18748 7976 19717 8004
rect 18748 7964 18754 7976
rect 19705 7973 19717 7976
rect 19751 8004 19763 8007
rect 20438 8004 20444 8016
rect 19751 7976 20444 8004
rect 19751 7973 19763 7976
rect 19705 7967 19763 7973
rect 20438 7964 20444 7976
rect 20496 7964 20502 8016
rect 20625 8007 20683 8013
rect 20625 7973 20637 8007
rect 20671 8004 20683 8007
rect 20898 8004 20904 8016
rect 20671 7976 20904 8004
rect 20671 7973 20683 7976
rect 20625 7967 20683 7973
rect 20898 7964 20904 7976
rect 20956 7964 20962 8016
rect 11048 7939 11106 7945
rect 11048 7905 11060 7939
rect 11094 7936 11106 7939
rect 11422 7936 11428 7948
rect 11094 7908 11428 7936
rect 11094 7905 11106 7908
rect 11048 7899 11106 7905
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 13354 7936 13360 7948
rect 13315 7908 13360 7936
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7936 17279 7939
rect 17586 7936 17592 7948
rect 17267 7908 17592 7936
rect 17267 7905 17279 7908
rect 17221 7899 17279 7905
rect 17586 7896 17592 7908
rect 17644 7896 17650 7948
rect 18874 7936 18880 7948
rect 18835 7908 18880 7936
rect 18874 7896 18880 7908
rect 18932 7896 18938 7948
rect 19610 7936 19616 7948
rect 19571 7908 19616 7936
rect 19610 7896 19616 7908
rect 19668 7896 19674 7948
rect 21266 7936 21272 7948
rect 21227 7908 21272 7936
rect 21266 7896 21272 7908
rect 21324 7896 21330 7948
rect 23750 7896 23756 7948
rect 23808 7936 23814 7948
rect 23928 7939 23986 7945
rect 23928 7936 23940 7939
rect 23808 7908 23940 7936
rect 23808 7896 23814 7908
rect 23928 7905 23940 7908
rect 23974 7936 23986 7939
rect 25038 7936 25044 7948
rect 23974 7908 25044 7936
rect 23974 7905 23986 7908
rect 23928 7899 23986 7905
rect 25038 7896 25044 7908
rect 25096 7896 25102 7948
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 10192 7840 10241 7868
rect 10192 7828 10198 7840
rect 10229 7837 10241 7840
rect 10275 7868 10287 7871
rect 10778 7868 10784 7880
rect 10275 7840 10784 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 12216 7840 13461 7868
rect 12216 7828 12222 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 12710 7760 12716 7812
rect 12768 7800 12774 7812
rect 13556 7800 13584 7831
rect 15562 7828 15568 7880
rect 15620 7868 15626 7880
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 15620 7840 15761 7868
rect 15620 7828 15626 7840
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7868 15899 7871
rect 15930 7868 15936 7880
rect 15887 7840 15936 7868
rect 15887 7837 15899 7840
rect 15841 7831 15899 7837
rect 12768 7772 13584 7800
rect 12768 7760 12774 7772
rect 13998 7760 14004 7812
rect 14056 7800 14062 7812
rect 15289 7803 15347 7809
rect 15289 7800 15301 7803
rect 14056 7772 15301 7800
rect 14056 7760 14062 7772
rect 15289 7769 15301 7772
rect 15335 7769 15347 7803
rect 15856 7800 15884 7831
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7837 17371 7871
rect 17494 7868 17500 7880
rect 17455 7840 17500 7868
rect 17313 7831 17371 7837
rect 15289 7763 15347 7769
rect 15764 7772 15884 7800
rect 14642 7732 14648 7744
rect 14603 7704 14648 7732
rect 14642 7692 14648 7704
rect 14700 7732 14706 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14700 7704 15025 7732
rect 14700 7692 14706 7704
rect 15013 7701 15025 7704
rect 15059 7732 15071 7735
rect 15764 7732 15792 7772
rect 17218 7760 17224 7812
rect 17276 7800 17282 7812
rect 17328 7800 17356 7831
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 18782 7828 18788 7880
rect 18840 7868 18846 7880
rect 19794 7868 19800 7880
rect 18840 7840 19800 7868
rect 18840 7828 18846 7840
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7868 19947 7871
rect 20254 7868 20260 7880
rect 19935 7840 20260 7868
rect 19935 7837 19947 7840
rect 19889 7831 19947 7837
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21726 7868 21732 7880
rect 21591 7840 21732 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22557 7871 22615 7877
rect 22557 7837 22569 7871
rect 22603 7868 22615 7871
rect 23290 7868 23296 7880
rect 22603 7840 23296 7868
rect 22603 7837 22615 7840
rect 22557 7831 22615 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 23661 7871 23719 7877
rect 23661 7868 23673 7871
rect 23492 7840 23673 7868
rect 17276 7772 17356 7800
rect 17276 7760 17282 7772
rect 19978 7760 19984 7812
rect 20036 7800 20042 7812
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 20036 7772 20913 7800
rect 20036 7760 20042 7772
rect 20901 7769 20913 7772
rect 20947 7769 20959 7803
rect 20901 7763 20959 7769
rect 16298 7732 16304 7744
rect 15059 7704 15792 7732
rect 16259 7704 16304 7732
rect 15059 7701 15071 7704
rect 15013 7695 15071 7701
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 18506 7732 18512 7744
rect 18467 7704 18512 7732
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 23198 7692 23204 7744
rect 23256 7732 23262 7744
rect 23492 7741 23520 7840
rect 23661 7837 23673 7840
rect 23707 7837 23719 7871
rect 23661 7831 23719 7837
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 23256 7704 23489 7732
rect 23256 7692 23262 7704
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12710 7528 12716 7540
rect 12308 7500 12716 7528
rect 12308 7488 12314 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 13081 7531 13139 7537
rect 13081 7497 13093 7531
rect 13127 7528 13139 7531
rect 13354 7528 13360 7540
rect 13127 7500 13360 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 10781 7463 10839 7469
rect 10781 7429 10793 7463
rect 10827 7460 10839 7463
rect 12158 7460 12164 7472
rect 10827 7432 12164 7460
rect 10827 7429 10839 7432
rect 10781 7423 10839 7429
rect 12158 7420 12164 7432
rect 12216 7420 12222 7472
rect 11422 7392 11428 7404
rect 11335 7364 11428 7392
rect 11422 7352 11428 7364
rect 11480 7392 11486 7404
rect 11882 7392 11888 7404
rect 11480 7364 11888 7392
rect 11480 7352 11486 7364
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 13096 7324 13124 7491
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15528 7500 15577 7528
rect 15528 7488 15534 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 15565 7491 15623 7497
rect 9815 7296 13124 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 13228 7296 13369 7324
rect 13228 7284 13234 7296
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 15580 7324 15608 7491
rect 17494 7488 17500 7540
rect 17552 7528 17558 7540
rect 17589 7531 17647 7537
rect 17589 7528 17601 7531
rect 17552 7500 17601 7528
rect 17552 7488 17558 7500
rect 17589 7497 17601 7500
rect 17635 7497 17647 7531
rect 18690 7528 18696 7540
rect 18651 7500 18696 7528
rect 17589 7491 17647 7497
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 19610 7488 19616 7540
rect 19668 7528 19674 7540
rect 19797 7531 19855 7537
rect 19797 7528 19809 7531
rect 19668 7500 19809 7528
rect 19668 7488 19674 7500
rect 19797 7497 19809 7500
rect 19843 7497 19855 7531
rect 20530 7528 20536 7540
rect 20491 7500 20536 7528
rect 19797 7491 19855 7497
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 21266 7488 21272 7540
rect 21324 7528 21330 7540
rect 21545 7531 21603 7537
rect 21545 7528 21557 7531
rect 21324 7500 21557 7528
rect 21324 7488 21330 7500
rect 21545 7497 21557 7500
rect 21591 7497 21603 7531
rect 21545 7491 21603 7497
rect 21818 7488 21824 7540
rect 21876 7528 21882 7540
rect 21913 7531 21971 7537
rect 21913 7528 21925 7531
rect 21876 7500 21925 7528
rect 21876 7488 21882 7500
rect 21913 7497 21925 7500
rect 21959 7497 21971 7531
rect 25038 7528 25044 7540
rect 24999 7500 25044 7528
rect 21913 7491 21971 7497
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 16298 7392 16304 7404
rect 16259 7364 16304 7392
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17586 7392 17592 7404
rect 16991 7364 17592 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7392 18383 7395
rect 18874 7392 18880 7404
rect 18371 7364 18880 7392
rect 18371 7361 18383 7364
rect 18325 7355 18383 7361
rect 18874 7352 18880 7364
rect 18932 7392 18938 7404
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 18932 7364 19349 7392
rect 18932 7352 18938 7364
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20956 7364 21005 7392
rect 20956 7352 20962 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 21174 7392 21180 7404
rect 21087 7364 21180 7392
rect 20993 7355 21051 7361
rect 21174 7352 21180 7364
rect 21232 7392 21238 7404
rect 21726 7392 21732 7404
rect 21232 7364 21732 7392
rect 21232 7352 21238 7364
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15580 7296 16129 7324
rect 13357 7287 13415 7293
rect 16117 7293 16129 7296
rect 16163 7293 16175 7327
rect 16117 7287 16175 7293
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7324 16267 7327
rect 16390 7324 16396 7336
rect 16255 7296 16396 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 10318 7256 10324 7268
rect 10231 7228 10324 7256
rect 10318 7216 10324 7228
rect 10376 7256 10382 7268
rect 11241 7259 11299 7265
rect 11241 7256 11253 7259
rect 10376 7228 11253 7256
rect 10376 7216 10382 7228
rect 11241 7225 11253 7228
rect 11287 7256 11299 7259
rect 11606 7256 11612 7268
rect 11287 7228 11612 7256
rect 11287 7225 11299 7228
rect 11241 7219 11299 7225
rect 11606 7216 11612 7228
rect 11664 7216 11670 7268
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 13602 7259 13660 7265
rect 13602 7256 13614 7259
rect 13504 7228 13614 7256
rect 13504 7216 13510 7228
rect 13602 7225 13614 7228
rect 13648 7256 13660 7259
rect 14642 7256 14648 7268
rect 13648 7228 14648 7256
rect 13648 7225 13660 7228
rect 13602 7219 13660 7225
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 15289 7259 15347 7265
rect 15289 7225 15301 7259
rect 15335 7256 15347 7259
rect 16224 7256 16252 7287
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 19150 7324 19156 7336
rect 19111 7296 19156 7324
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7324 22431 7327
rect 22419 7296 23060 7324
rect 22419 7293 22431 7296
rect 22373 7287 22431 7293
rect 15335 7228 16252 7256
rect 15335 7225 15347 7228
rect 15289 7219 15347 7225
rect 18690 7216 18696 7268
rect 18748 7256 18754 7268
rect 19245 7259 19303 7265
rect 19245 7256 19257 7259
rect 18748 7228 19257 7256
rect 18748 7216 18754 7228
rect 19245 7225 19257 7228
rect 19291 7225 19303 7259
rect 19245 7219 19303 7225
rect 20901 7259 20959 7265
rect 20901 7225 20913 7259
rect 20947 7256 20959 7259
rect 21818 7256 21824 7268
rect 20947 7228 21824 7256
rect 20947 7225 20959 7228
rect 20901 7219 20959 7225
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 9180 7160 10609 7188
rect 9180 7148 9186 7160
rect 10597 7157 10609 7160
rect 10643 7188 10655 7191
rect 10870 7188 10876 7200
rect 10643 7160 10876 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 10870 7148 10876 7160
rect 10928 7188 10934 7200
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 10928 7160 11161 7188
rect 10928 7148 10934 7160
rect 11149 7157 11161 7160
rect 11195 7157 11207 7191
rect 11882 7188 11888 7200
rect 11843 7160 11888 7188
rect 11149 7151 11207 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15746 7188 15752 7200
rect 15707 7160 15752 7188
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 17218 7188 17224 7200
rect 17179 7160 17224 7188
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 18785 7191 18843 7197
rect 18785 7157 18797 7191
rect 18831 7188 18843 7191
rect 19058 7188 19064 7200
rect 18831 7160 19064 7188
rect 18831 7157 18843 7160
rect 18785 7151 18843 7157
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 22557 7191 22615 7197
rect 22557 7157 22569 7191
rect 22603 7188 22615 7191
rect 22738 7188 22744 7200
rect 22603 7160 22744 7188
rect 22603 7157 22615 7160
rect 22557 7151 22615 7157
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 23032 7197 23060 7296
rect 23198 7284 23204 7336
rect 23256 7324 23262 7336
rect 23661 7327 23719 7333
rect 23661 7324 23673 7327
rect 23256 7296 23673 7324
rect 23256 7284 23262 7296
rect 23661 7293 23673 7296
rect 23707 7324 23719 7327
rect 25317 7327 25375 7333
rect 25317 7324 25329 7327
rect 23707 7296 25329 7324
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 25317 7293 25329 7296
rect 25363 7293 25375 7327
rect 25317 7287 25375 7293
rect 23934 7265 23940 7268
rect 23477 7259 23535 7265
rect 23477 7225 23489 7259
rect 23523 7256 23535 7259
rect 23928 7256 23940 7265
rect 23523 7228 23940 7256
rect 23523 7225 23535 7228
rect 23477 7219 23535 7225
rect 23928 7219 23940 7228
rect 23934 7216 23940 7219
rect 23992 7216 23998 7268
rect 23017 7191 23075 7197
rect 23017 7157 23029 7191
rect 23063 7188 23075 7191
rect 23382 7188 23388 7200
rect 23063 7160 23388 7188
rect 23063 7157 23075 7160
rect 23017 7151 23075 7157
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 11149 6987 11207 6993
rect 11149 6953 11161 6987
rect 11195 6984 11207 6987
rect 11517 6987 11575 6993
rect 11517 6984 11529 6987
rect 11195 6956 11529 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11517 6953 11529 6956
rect 11563 6984 11575 6987
rect 11882 6984 11888 6996
rect 11563 6956 11888 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 12894 6984 12900 6996
rect 12115 6956 12900 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 13446 6984 13452 6996
rect 13407 6956 13452 6984
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 13998 6984 14004 6996
rect 13780 6956 14004 6984
rect 13780 6944 13786 6956
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 14737 6987 14795 6993
rect 14737 6953 14749 6987
rect 14783 6984 14795 6987
rect 15562 6984 15568 6996
rect 14783 6956 15568 6984
rect 14783 6953 14795 6956
rect 14737 6947 14795 6953
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 18141 6987 18199 6993
rect 18141 6953 18153 6987
rect 18187 6984 18199 6987
rect 18322 6984 18328 6996
rect 18187 6956 18328 6984
rect 18187 6953 18199 6956
rect 18141 6947 18199 6953
rect 18322 6944 18328 6956
rect 18380 6984 18386 6996
rect 19150 6984 19156 6996
rect 18380 6956 19156 6984
rect 18380 6944 18386 6956
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19613 6987 19671 6993
rect 19613 6984 19625 6987
rect 19576 6956 19625 6984
rect 19576 6944 19582 6956
rect 19613 6953 19625 6956
rect 19659 6953 19671 6987
rect 19613 6947 19671 6953
rect 20625 6987 20683 6993
rect 20625 6953 20637 6987
rect 20671 6984 20683 6987
rect 21174 6984 21180 6996
rect 20671 6956 21180 6984
rect 20671 6953 20683 6956
rect 20625 6947 20683 6953
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 22649 6987 22707 6993
rect 22649 6953 22661 6987
rect 22695 6953 22707 6987
rect 23750 6984 23756 6996
rect 23711 6956 23756 6984
rect 22649 6947 22707 6953
rect 9784 6888 10364 6916
rect 9784 6857 9812 6888
rect 10336 6860 10364 6888
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 12492 6888 12537 6916
rect 12492 6876 12498 6888
rect 15654 6876 15660 6928
rect 15712 6916 15718 6928
rect 15841 6919 15899 6925
rect 15841 6916 15853 6919
rect 15712 6888 15853 6916
rect 15712 6876 15718 6888
rect 15841 6885 15853 6888
rect 15887 6916 15899 6919
rect 16485 6919 16543 6925
rect 16485 6916 16497 6919
rect 15887 6888 16497 6916
rect 15887 6885 15899 6888
rect 15841 6879 15899 6885
rect 16485 6885 16497 6888
rect 16531 6885 16543 6919
rect 16485 6879 16543 6885
rect 17862 6876 17868 6928
rect 17920 6916 17926 6928
rect 18049 6919 18107 6925
rect 18049 6916 18061 6919
rect 17920 6888 18061 6916
rect 17920 6876 17926 6888
rect 18049 6885 18061 6888
rect 18095 6916 18107 6919
rect 18095 6888 19380 6916
rect 18095 6885 18107 6888
rect 18049 6879 18107 6885
rect 19352 6860 19380 6888
rect 20254 6876 20260 6928
rect 20312 6916 20318 6928
rect 22664 6916 22692 6947
rect 23750 6944 23756 6956
rect 23808 6944 23814 6996
rect 20312 6888 22692 6916
rect 23768 6916 23796 6944
rect 23768 6888 24348 6916
rect 20312 6876 20318 6888
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10025 6851 10083 6857
rect 10025 6848 10037 6851
rect 9916 6820 10037 6848
rect 9916 6808 9922 6820
rect 10025 6817 10037 6820
rect 10071 6817 10083 6851
rect 10025 6811 10083 6817
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 10376 6820 11989 6848
rect 10376 6808 10382 6820
rect 11977 6817 11989 6820
rect 12023 6848 12035 6851
rect 13170 6848 13176 6860
rect 12023 6820 13176 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 14884 6820 15025 6848
rect 14884 6808 14890 6820
rect 15013 6817 15025 6820
rect 15059 6817 15071 6851
rect 15013 6811 15071 6817
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 17184 6820 17233 6848
rect 17184 6808 17190 6820
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 17494 6848 17500 6860
rect 17455 6820 17500 6848
rect 17221 6811 17279 6817
rect 17494 6808 17500 6820
rect 17552 6848 17558 6860
rect 17552 6820 18276 6848
rect 17552 6808 17558 6820
rect 12526 6780 12532 6792
rect 12487 6752 12532 6780
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 12710 6780 12716 6792
rect 12671 6752 12716 6780
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13320 6752 14105 6780
rect 13320 6740 13326 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14274 6780 14280 6792
rect 14187 6752 14280 6780
rect 14093 6743 14151 6749
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 13004 6684 13645 6712
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 13004 6644 13032 6684
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 14108 6712 14136 6743
rect 14274 6740 14280 6752
rect 14332 6780 14338 6792
rect 14734 6780 14740 6792
rect 14332 6752 14740 6780
rect 14332 6740 14338 6752
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15933 6783 15991 6789
rect 15933 6780 15945 6783
rect 15344 6752 15945 6780
rect 15344 6740 15350 6752
rect 15933 6749 15945 6752
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16666 6780 16672 6792
rect 16163 6752 16672 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 18248 6789 18276 6820
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 19392 6820 19717 6848
rect 19392 6808 19398 6820
rect 19705 6817 19717 6820
rect 19751 6848 19763 6851
rect 20070 6848 20076 6860
rect 19751 6820 20076 6848
rect 19751 6817 19763 6820
rect 19705 6811 19763 6817
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 21082 6808 21088 6860
rect 21140 6848 21146 6860
rect 21525 6851 21583 6857
rect 21525 6848 21537 6851
rect 21140 6820 21537 6848
rect 21140 6808 21146 6820
rect 21525 6817 21537 6820
rect 21571 6817 21583 6851
rect 24210 6848 24216 6860
rect 24171 6820 24216 6848
rect 21525 6811 21583 6817
rect 24210 6808 24216 6820
rect 24268 6808 24274 6860
rect 24320 6848 24348 6888
rect 24320 6820 24440 6848
rect 18233 6783 18291 6789
rect 18233 6749 18245 6783
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 19889 6783 19947 6789
rect 19889 6749 19901 6783
rect 19935 6780 19947 6783
rect 20162 6780 20168 6792
rect 19935 6752 20168 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 21266 6780 21272 6792
rect 21227 6752 21272 6780
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 23106 6740 23112 6792
rect 23164 6780 23170 6792
rect 24412 6789 24440 6820
rect 24305 6783 24363 6789
rect 24305 6780 24317 6783
rect 23164 6752 24317 6780
rect 23164 6740 23170 6752
rect 24305 6749 24317 6752
rect 24351 6749 24363 6783
rect 24305 6743 24363 6749
rect 24397 6783 24455 6789
rect 24397 6749 24409 6783
rect 24443 6749 24455 6783
rect 25406 6780 25412 6792
rect 25367 6752 25412 6780
rect 24397 6743 24455 6749
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 15102 6712 15108 6724
rect 14108 6684 15108 6712
rect 13633 6675 13691 6681
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 15746 6672 15752 6724
rect 15804 6712 15810 6724
rect 16390 6712 16396 6724
rect 15804 6684 16396 6712
rect 15804 6672 15810 6684
rect 16390 6672 16396 6684
rect 16448 6712 16454 6724
rect 16853 6715 16911 6721
rect 16853 6712 16865 6715
rect 16448 6684 16865 6712
rect 16448 6672 16454 6684
rect 16853 6681 16865 6684
rect 16899 6681 16911 6715
rect 17678 6712 17684 6724
rect 17639 6684 17684 6712
rect 16853 6675 16911 6681
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 12400 6616 13032 6644
rect 15473 6647 15531 6653
rect 12400 6604 12406 6616
rect 15473 6613 15485 6647
rect 15519 6644 15531 6647
rect 16022 6644 16028 6656
rect 15519 6616 16028 6644
rect 15519 6613 15531 6616
rect 15473 6607 15531 6613
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 17037 6647 17095 6653
rect 17037 6613 17049 6647
rect 17083 6644 17095 6647
rect 17218 6644 17224 6656
rect 17083 6616 17224 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 18785 6647 18843 6653
rect 18785 6644 18797 6647
rect 18748 6616 18797 6644
rect 18748 6604 18754 6616
rect 18785 6613 18797 6616
rect 18831 6613 18843 6647
rect 19242 6644 19248 6656
rect 19203 6616 19248 6644
rect 18785 6607 18843 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 22278 6644 22284 6656
rect 21324 6616 22284 6644
rect 21324 6604 21330 6616
rect 22278 6604 22284 6616
rect 22336 6644 22342 6656
rect 22925 6647 22983 6653
rect 22925 6644 22937 6647
rect 22336 6616 22937 6644
rect 22336 6604 22342 6616
rect 22925 6613 22937 6616
rect 22971 6644 22983 6647
rect 23198 6644 23204 6656
rect 22971 6616 23204 6644
rect 22971 6613 22983 6616
rect 22925 6607 22983 6613
rect 23198 6604 23204 6616
rect 23256 6644 23262 6656
rect 23293 6647 23351 6653
rect 23293 6644 23305 6647
rect 23256 6616 23305 6644
rect 23256 6604 23262 6616
rect 23293 6613 23305 6616
rect 23339 6613 23351 6647
rect 23842 6644 23848 6656
rect 23803 6616 23848 6644
rect 23293 6607 23351 6613
rect 23842 6604 23848 6616
rect 23900 6604 23906 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 9858 6440 9864 6452
rect 9819 6412 9864 6440
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10229 6443 10287 6449
rect 10229 6409 10241 6443
rect 10275 6440 10287 6443
rect 10318 6440 10324 6452
rect 10275 6412 10324 6440
rect 10275 6409 10287 6412
rect 10229 6403 10287 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10778 6440 10784 6452
rect 10739 6412 10784 6440
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6440 12219 6443
rect 12710 6440 12716 6452
rect 12207 6412 12716 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 12897 6443 12955 6449
rect 12897 6409 12909 6443
rect 12943 6440 12955 6443
rect 13722 6440 13728 6452
rect 12943 6412 13728 6440
rect 12943 6409 12955 6412
rect 12897 6403 12955 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 15105 6443 15163 6449
rect 15105 6409 15117 6443
rect 15151 6440 15163 6443
rect 15562 6440 15568 6452
rect 15151 6412 15568 6440
rect 15151 6409 15163 6412
rect 15105 6403 15163 6409
rect 15562 6400 15568 6412
rect 15620 6440 15626 6452
rect 16298 6440 16304 6452
rect 15620 6412 16304 6440
rect 15620 6400 15626 6412
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 17773 6443 17831 6449
rect 17773 6409 17785 6443
rect 17819 6440 17831 6443
rect 17862 6440 17868 6452
rect 17819 6412 17868 6440
rect 17819 6409 17831 6412
rect 17773 6403 17831 6409
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 18322 6440 18328 6452
rect 18283 6412 18328 6440
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 19668 6412 20361 6440
rect 19668 6400 19674 6412
rect 20349 6409 20361 6412
rect 20395 6409 20407 6443
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 20349 6403 20407 6409
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 23750 6440 23756 6452
rect 23523 6412 23756 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 23750 6400 23756 6412
rect 23808 6400 23814 6452
rect 24210 6400 24216 6452
rect 24268 6440 24274 6452
rect 24489 6443 24547 6449
rect 24489 6440 24501 6443
rect 24268 6412 24501 6440
rect 24268 6400 24274 6412
rect 24489 6409 24501 6412
rect 24535 6440 24547 6443
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 24535 6412 25513 6440
rect 24535 6409 24547 6412
rect 24489 6403 24547 6409
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 11425 6375 11483 6381
rect 11425 6341 11437 6375
rect 11471 6372 11483 6375
rect 12434 6372 12440 6384
rect 11471 6344 12440 6372
rect 11471 6341 11483 6344
rect 11425 6335 11483 6341
rect 12434 6332 12440 6344
rect 12492 6332 12498 6384
rect 13262 6372 13268 6384
rect 13223 6344 13268 6372
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 20993 6375 21051 6381
rect 20993 6372 21005 6375
rect 20732 6344 21005 6372
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6304 11851 6307
rect 12526 6304 12532 6316
rect 11839 6276 12532 6304
rect 11839 6273 11851 6276
rect 11793 6267 11851 6273
rect 12526 6264 12532 6276
rect 12584 6304 12590 6316
rect 13446 6304 13452 6316
rect 12584 6276 13452 6304
rect 12584 6264 12590 6276
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6304 13691 6307
rect 16390 6304 16396 6316
rect 13679 6276 13860 6304
rect 16351 6276 16396 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 13832 6248 13860 6276
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 16577 6307 16635 6313
rect 16577 6273 16589 6307
rect 16623 6304 16635 6307
rect 16666 6304 16672 6316
rect 16623 6276 16672 6304
rect 16623 6273 16635 6276
rect 16577 6267 16635 6273
rect 13170 6196 13176 6248
rect 13228 6236 13234 6248
rect 13722 6236 13728 6248
rect 13228 6208 13728 6236
rect 13228 6196 13234 6208
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 13992 6239 14050 6245
rect 13992 6236 14004 6239
rect 13872 6208 14004 6236
rect 13872 6196 13878 6208
rect 13992 6205 14004 6208
rect 14038 6236 14050 6239
rect 14274 6236 14280 6248
rect 14038 6208 14280 6236
rect 14038 6205 14050 6208
rect 13992 6199 14050 6205
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6236 15531 6239
rect 16592 6236 16620 6267
rect 16666 6264 16672 6276
rect 16724 6304 16730 6316
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16724 6276 16957 6304
rect 16724 6264 16730 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18564 6276 18705 6304
rect 18564 6264 18570 6276
rect 18693 6273 18705 6276
rect 18739 6273 18751 6307
rect 18693 6267 18751 6273
rect 15519 6208 16620 6236
rect 18708 6236 18736 6267
rect 19978 6236 19984 6248
rect 18708 6208 19984 6236
rect 15519 6205 15531 6208
rect 15473 6199 15531 6205
rect 19978 6196 19984 6208
rect 20036 6236 20042 6248
rect 20732 6236 20760 6344
rect 20993 6341 21005 6344
rect 21039 6372 21051 6375
rect 21266 6372 21272 6384
rect 21039 6344 21272 6372
rect 21039 6341 21051 6344
rect 20993 6335 21051 6341
rect 21266 6332 21272 6344
rect 21324 6372 21330 6384
rect 22741 6375 22799 6381
rect 21324 6344 21404 6372
rect 21324 6332 21330 6344
rect 21376 6313 21404 6344
rect 22741 6341 22753 6375
rect 22787 6341 22799 6375
rect 22741 6335 22799 6341
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6273 21419 6307
rect 22756 6304 22784 6335
rect 23934 6304 23940 6316
rect 22756 6276 23940 6304
rect 21361 6267 21419 6273
rect 23934 6264 23940 6276
rect 23992 6304 23998 6316
rect 25130 6304 25136 6316
rect 23992 6276 25136 6304
rect 23992 6264 23998 6276
rect 25130 6264 25136 6276
rect 25188 6264 25194 6316
rect 20036 6208 20760 6236
rect 20036 6196 20042 6208
rect 20990 6196 20996 6248
rect 21048 6236 21054 6248
rect 21177 6239 21235 6245
rect 21177 6236 21189 6239
rect 21048 6208 21189 6236
rect 21048 6196 21054 6208
rect 21177 6205 21189 6208
rect 21223 6236 21235 6239
rect 21450 6236 21456 6248
rect 21223 6208 21456 6236
rect 21223 6205 21235 6208
rect 21177 6199 21235 6205
rect 21450 6196 21456 6208
rect 21508 6196 21514 6248
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 15764 6140 16313 6168
rect 15764 6112 15792 6140
rect 16301 6137 16313 6140
rect 16347 6137 16359 6171
rect 16301 6131 16359 6137
rect 17405 6171 17463 6177
rect 17405 6137 17417 6171
rect 17451 6168 17463 6171
rect 18874 6168 18880 6180
rect 17451 6140 18880 6168
rect 17451 6137 17463 6140
rect 17405 6131 17463 6137
rect 18874 6128 18880 6140
rect 18932 6177 18938 6180
rect 18932 6171 18996 6177
rect 18932 6137 18950 6171
rect 18984 6137 18996 6171
rect 18932 6131 18996 6137
rect 20901 6171 20959 6177
rect 20901 6137 20913 6171
rect 20947 6168 20959 6171
rect 21082 6168 21088 6180
rect 20947 6140 21088 6168
rect 20947 6137 20959 6140
rect 20901 6131 20959 6137
rect 18932 6128 18938 6131
rect 21082 6128 21088 6140
rect 21140 6128 21146 6180
rect 21634 6177 21640 6180
rect 21628 6168 21640 6177
rect 21595 6140 21640 6168
rect 21628 6131 21640 6140
rect 21634 6128 21640 6131
rect 21692 6128 21698 6180
rect 23750 6128 23756 6180
rect 23808 6168 23814 6180
rect 23937 6171 23995 6177
rect 23937 6168 23949 6171
rect 23808 6140 23949 6168
rect 23808 6128 23814 6140
rect 23937 6137 23949 6140
rect 23983 6168 23995 6171
rect 24857 6171 24915 6177
rect 24857 6168 24869 6171
rect 23983 6140 24869 6168
rect 23983 6137 23995 6140
rect 23937 6131 23995 6137
rect 24857 6137 24869 6140
rect 24903 6137 24915 6171
rect 24857 6131 24915 6137
rect 14182 6060 14188 6112
rect 14240 6100 14246 6112
rect 14642 6100 14648 6112
rect 14240 6072 14648 6100
rect 14240 6060 14246 6072
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15746 6100 15752 6112
rect 15707 6072 15752 6100
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 20073 6103 20131 6109
rect 20073 6069 20085 6103
rect 20119 6100 20131 6103
rect 20162 6100 20168 6112
rect 20119 6072 20168 6100
rect 20119 6069 20131 6072
rect 20073 6063 20131 6069
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 22922 6060 22928 6112
rect 22980 6100 22986 6112
rect 24397 6103 24455 6109
rect 24397 6100 24409 6103
rect 22980 6072 24409 6100
rect 22980 6060 22986 6072
rect 24397 6069 24409 6072
rect 24443 6100 24455 6103
rect 24949 6103 25007 6109
rect 24949 6100 24961 6103
rect 24443 6072 24961 6100
rect 24443 6069 24455 6072
rect 24397 6063 24455 6069
rect 24949 6069 24961 6072
rect 24995 6100 25007 6103
rect 25314 6100 25320 6112
rect 24995 6072 25320 6100
rect 24995 6069 25007 6072
rect 24949 6063 25007 6069
rect 25314 6060 25320 6072
rect 25372 6060 25378 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 12066 5896 12072 5908
rect 12027 5868 12072 5896
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 13814 5896 13820 5908
rect 13775 5868 13820 5896
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 14274 5856 14280 5908
rect 14332 5896 14338 5908
rect 15105 5899 15163 5905
rect 15105 5896 15117 5899
rect 14332 5868 15117 5896
rect 14332 5856 14338 5868
rect 15105 5865 15117 5868
rect 15151 5896 15163 5899
rect 15286 5896 15292 5908
rect 15151 5868 15292 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 17126 5896 17132 5908
rect 17087 5868 17132 5896
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 18874 5896 18880 5908
rect 18835 5868 18880 5896
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 19334 5896 19340 5908
rect 19295 5868 19340 5896
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 20714 5896 20720 5908
rect 20675 5868 20720 5896
rect 20714 5856 20720 5868
rect 20772 5896 20778 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 20772 5868 21281 5896
rect 20772 5856 20778 5868
rect 21269 5865 21281 5868
rect 21315 5865 21327 5899
rect 21269 5859 21327 5865
rect 21450 5856 21456 5908
rect 21508 5896 21514 5908
rect 22281 5899 22339 5905
rect 22281 5896 22293 5899
rect 21508 5868 22293 5896
rect 21508 5856 21514 5868
rect 22281 5865 22293 5868
rect 22327 5865 22339 5899
rect 22281 5859 22339 5865
rect 23106 5856 23112 5908
rect 23164 5896 23170 5908
rect 23569 5899 23627 5905
rect 23569 5896 23581 5899
rect 23164 5868 23581 5896
rect 23164 5856 23170 5868
rect 23569 5865 23581 5868
rect 23615 5865 23627 5899
rect 23569 5859 23627 5865
rect 15562 5837 15568 5840
rect 15556 5828 15568 5837
rect 15523 5800 15568 5828
rect 15556 5791 15568 5800
rect 15562 5788 15568 5791
rect 15620 5788 15626 5840
rect 24029 5831 24087 5837
rect 24029 5797 24041 5831
rect 24075 5828 24087 5831
rect 24118 5828 24124 5840
rect 24075 5800 24124 5828
rect 24075 5797 24087 5800
rect 24029 5791 24087 5797
rect 24118 5788 24124 5800
rect 24176 5788 24182 5840
rect 12989 5763 13047 5769
rect 12989 5729 13001 5763
rect 13035 5760 13047 5763
rect 13722 5760 13728 5772
rect 13035 5732 13728 5760
rect 13035 5729 13047 5732
rect 12989 5723 13047 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5760 14151 5763
rect 14182 5760 14188 5772
rect 14139 5732 14188 5760
rect 14139 5729 14151 5732
rect 14093 5723 14151 5729
rect 14182 5720 14188 5732
rect 14240 5760 14246 5772
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 14240 5732 14657 5760
rect 14240 5720 14246 5732
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 17753 5763 17811 5769
rect 17753 5760 17765 5763
rect 17644 5732 17765 5760
rect 17644 5720 17650 5732
rect 17753 5729 17765 5732
rect 17799 5729 17811 5763
rect 19702 5760 19708 5772
rect 19615 5732 19708 5760
rect 17753 5723 17811 5729
rect 19702 5720 19708 5732
rect 19760 5760 19766 5772
rect 20346 5760 20352 5772
rect 19760 5732 20352 5760
rect 19760 5720 19766 5732
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 23106 5720 23112 5772
rect 23164 5760 23170 5772
rect 23937 5763 23995 5769
rect 23937 5760 23949 5763
rect 23164 5732 23949 5760
rect 23164 5720 23170 5732
rect 23937 5729 23949 5732
rect 23983 5729 23995 5763
rect 23937 5723 23995 5729
rect 24854 5720 24860 5772
rect 24912 5760 24918 5772
rect 25133 5763 25191 5769
rect 25133 5760 25145 5763
rect 24912 5732 25145 5760
rect 24912 5720 24918 5732
rect 25133 5729 25145 5732
rect 25179 5729 25191 5763
rect 25133 5723 25191 5729
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13170 5692 13176 5704
rect 13127 5664 13176 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 15286 5692 15292 5704
rect 15247 5664 15292 5692
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 17126 5652 17132 5704
rect 17184 5692 17190 5704
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17184 5664 17509 5692
rect 17184 5652 17190 5664
rect 17497 5661 17509 5664
rect 17543 5661 17555 5695
rect 21358 5692 21364 5704
rect 21319 5664 21364 5692
rect 17497 5655 17555 5661
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21634 5692 21640 5704
rect 21591 5664 21640 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21634 5652 21640 5664
rect 21692 5692 21698 5704
rect 21913 5695 21971 5701
rect 21913 5692 21925 5695
rect 21692 5664 21925 5692
rect 21692 5652 21698 5664
rect 21913 5661 21925 5664
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5661 24271 5695
rect 24213 5655 24271 5661
rect 22649 5627 22707 5633
rect 22649 5593 22661 5627
rect 22695 5624 22707 5627
rect 23934 5624 23940 5636
rect 22695 5596 23940 5624
rect 22695 5593 22707 5596
rect 22649 5587 22707 5593
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 24228 5624 24256 5655
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 24228 5596 24685 5624
rect 24673 5593 24685 5596
rect 24719 5624 24731 5627
rect 25130 5624 25136 5636
rect 24719 5596 25136 5624
rect 24719 5593 24731 5596
rect 24673 5587 24731 5593
rect 25130 5584 25136 5596
rect 25188 5584 25194 5636
rect 14277 5559 14335 5565
rect 14277 5525 14289 5559
rect 14323 5556 14335 5559
rect 14826 5556 14832 5568
rect 14323 5528 14832 5556
rect 14323 5525 14335 5528
rect 14277 5519 14335 5525
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 16666 5556 16672 5568
rect 16627 5528 16672 5556
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5556 19947 5559
rect 20070 5556 20076 5568
rect 19935 5528 20076 5556
rect 19935 5525 19947 5528
rect 19889 5519 19947 5525
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 20162 5516 20168 5568
rect 20220 5556 20226 5568
rect 20257 5559 20315 5565
rect 20257 5556 20269 5559
rect 20220 5528 20269 5556
rect 20220 5516 20226 5528
rect 20257 5525 20269 5528
rect 20303 5525 20315 5559
rect 20898 5556 20904 5568
rect 20859 5528 20904 5556
rect 20257 5519 20315 5525
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 22278 5556 22284 5568
rect 22152 5528 22284 5556
rect 22152 5516 22158 5528
rect 22278 5516 22284 5528
rect 22336 5556 22342 5568
rect 23017 5559 23075 5565
rect 23017 5556 23029 5559
rect 22336 5528 23029 5556
rect 22336 5516 22342 5528
rect 23017 5525 23029 5528
rect 23063 5556 23075 5559
rect 23198 5556 23204 5568
rect 23063 5528 23204 5556
rect 23063 5525 23075 5528
rect 23017 5519 23075 5525
rect 23198 5516 23204 5528
rect 23256 5556 23262 5568
rect 23385 5559 23443 5565
rect 23385 5556 23397 5559
rect 23256 5528 23397 5556
rect 23256 5516 23262 5528
rect 23385 5525 23397 5528
rect 23431 5556 23443 5559
rect 24949 5559 25007 5565
rect 24949 5556 24961 5559
rect 23431 5528 24961 5556
rect 23431 5525 23443 5528
rect 23385 5519 23443 5525
rect 24949 5525 24961 5528
rect 24995 5525 25007 5559
rect 24949 5519 25007 5525
rect 25317 5559 25375 5565
rect 25317 5525 25329 5559
rect 25363 5556 25375 5559
rect 25498 5556 25504 5568
rect 25363 5528 25504 5556
rect 25363 5525 25375 5528
rect 25317 5519 25375 5525
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 13725 5355 13783 5361
rect 13725 5352 13737 5355
rect 12492 5324 13737 5352
rect 12492 5312 12498 5324
rect 13725 5321 13737 5324
rect 13771 5352 13783 5355
rect 13906 5352 13912 5364
rect 13771 5324 13912 5352
rect 13771 5321 13783 5324
rect 13725 5315 13783 5321
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14185 5355 14243 5361
rect 14185 5321 14197 5355
rect 14231 5352 14243 5355
rect 14274 5352 14280 5364
rect 14231 5324 14280 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15562 5352 15568 5364
rect 15427 5324 15568 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 13924 5216 13952 5312
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 13924 5188 14657 5216
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14792 5188 14841 5216
rect 14792 5176 14798 5188
rect 14829 5185 14841 5188
rect 14875 5216 14887 5219
rect 15396 5216 15424 5315
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 21361 5355 21419 5361
rect 21361 5321 21373 5355
rect 21407 5352 21419 5355
rect 21634 5352 21640 5364
rect 21407 5324 21640 5352
rect 21407 5321 21419 5324
rect 21361 5315 21419 5321
rect 21634 5312 21640 5324
rect 21692 5312 21698 5364
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22281 5355 22339 5361
rect 22281 5352 22293 5355
rect 22244 5324 22293 5352
rect 22244 5312 22250 5324
rect 22281 5321 22293 5324
rect 22327 5321 22339 5355
rect 22281 5315 22339 5321
rect 14875 5188 15424 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 18874 5176 18880 5228
rect 18932 5216 18938 5228
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 18932 5188 18981 5216
rect 18932 5176 18938 5188
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 19978 5216 19984 5228
rect 19939 5188 19984 5216
rect 18969 5179 19027 5185
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12912 5120 13093 5148
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 12912 5021 12940 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 14093 5151 14151 5157
rect 14093 5117 14105 5151
rect 14139 5148 14151 5151
rect 14550 5148 14556 5160
rect 14139 5120 14556 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 15286 5108 15292 5160
rect 15344 5148 15350 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15344 5120 15761 5148
rect 15344 5108 15350 5120
rect 15749 5117 15761 5120
rect 15795 5148 15807 5151
rect 17126 5148 17132 5160
rect 15795 5120 17132 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 17126 5108 17132 5120
rect 17184 5108 17190 5160
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5148 18383 5151
rect 18782 5148 18788 5160
rect 18371 5120 18788 5148
rect 18371 5117 18383 5120
rect 18325 5111 18383 5117
rect 18782 5108 18788 5120
rect 18840 5108 18846 5160
rect 22296 5148 22324 5315
rect 22462 5312 22468 5364
rect 22520 5352 22526 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22520 5324 23029 5352
rect 22520 5312 22526 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 23017 5315 23075 5321
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 23164 5324 23397 5352
rect 23164 5312 23170 5324
rect 23385 5321 23397 5324
rect 23431 5352 23443 5355
rect 23431 5324 24716 5352
rect 23431 5321 23443 5324
rect 23385 5315 23443 5321
rect 23198 5176 23204 5228
rect 23256 5216 23262 5228
rect 23661 5219 23719 5225
rect 23661 5216 23673 5219
rect 23256 5188 23673 5216
rect 23256 5176 23262 5188
rect 23661 5185 23673 5188
rect 23707 5185 23719 5219
rect 24688 5216 24716 5324
rect 25130 5312 25136 5364
rect 25188 5352 25194 5364
rect 25317 5355 25375 5361
rect 25317 5352 25329 5355
rect 25188 5324 25329 5352
rect 25188 5312 25194 5324
rect 25317 5321 25329 5324
rect 25363 5321 25375 5355
rect 25317 5315 25375 5321
rect 24762 5244 24768 5296
rect 24820 5284 24826 5296
rect 25038 5284 25044 5296
rect 24820 5256 25044 5284
rect 24820 5244 24826 5256
rect 25038 5244 25044 5256
rect 25096 5244 25102 5296
rect 25130 5216 25136 5228
rect 24688 5188 25136 5216
rect 23661 5179 23719 5185
rect 25130 5176 25136 5188
rect 25188 5176 25194 5228
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22296 5120 22477 5148
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 16016 5083 16074 5089
rect 16016 5049 16028 5083
rect 16062 5080 16074 5083
rect 16666 5080 16672 5092
rect 16062 5052 16672 5080
rect 16062 5049 16074 5052
rect 16016 5043 16074 5049
rect 16666 5040 16672 5052
rect 16724 5040 16730 5092
rect 20162 5040 20168 5092
rect 20220 5089 20226 5092
rect 20220 5083 20284 5089
rect 20220 5049 20238 5083
rect 20272 5049 20284 5083
rect 20220 5043 20284 5049
rect 20220 5040 20226 5043
rect 23750 5040 23756 5092
rect 23808 5080 23814 5092
rect 23906 5083 23964 5089
rect 23906 5080 23918 5083
rect 23808 5052 23918 5080
rect 23808 5040 23814 5052
rect 23906 5049 23918 5052
rect 23952 5049 23964 5083
rect 23906 5043 23964 5049
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12676 4984 12909 5012
rect 12676 4972 12682 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 13262 5012 13268 5024
rect 13223 4984 13268 5012
rect 12897 4975 12955 4981
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 17129 5015 17187 5021
rect 17129 5012 17141 5015
rect 16172 4984 17141 5012
rect 16172 4972 16178 4984
rect 17129 4981 17141 4984
rect 17175 5012 17187 5015
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17175 4984 17509 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17497 4981 17509 4984
rect 17543 5012 17555 5015
rect 17586 5012 17592 5024
rect 17543 4984 17592 5012
rect 17543 4981 17555 4984
rect 17497 4975 17555 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 18840 4984 18889 5012
rect 18840 4972 18846 4984
rect 18877 4981 18889 4984
rect 18923 4981 18935 5015
rect 22646 5012 22652 5024
rect 22607 4984 22652 5012
rect 18877 4975 18935 4981
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 24854 4972 24860 5024
rect 24912 5012 24918 5024
rect 25685 5015 25743 5021
rect 25685 5012 25697 5015
rect 24912 4984 25697 5012
rect 24912 4972 24918 4984
rect 25685 4981 25697 4984
rect 25731 4981 25743 5015
rect 25685 4975 25743 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 13722 4808 13728 4820
rect 13035 4780 13728 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14734 4808 14740 4820
rect 14695 4780 14740 4808
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4808 15163 4811
rect 15930 4808 15936 4820
rect 15151 4780 15936 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16666 4808 16672 4820
rect 16080 4780 16125 4808
rect 16627 4780 16672 4808
rect 16080 4768 16086 4780
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 16758 4768 16764 4820
rect 16816 4808 16822 4820
rect 17313 4811 17371 4817
rect 17313 4808 17325 4811
rect 16816 4780 17325 4808
rect 16816 4768 16822 4780
rect 17313 4777 17325 4780
rect 17359 4777 17371 4811
rect 17678 4808 17684 4820
rect 17639 4780 17684 4808
rect 17313 4771 17371 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18877 4811 18935 4817
rect 18877 4777 18889 4811
rect 18923 4808 18935 4811
rect 21358 4808 21364 4820
rect 18923 4780 21364 4808
rect 18923 4777 18935 4780
rect 18877 4771 18935 4777
rect 21358 4768 21364 4780
rect 21416 4808 21422 4820
rect 21637 4811 21695 4817
rect 21637 4808 21649 4811
rect 21416 4780 21649 4808
rect 21416 4768 21422 4780
rect 21637 4777 21649 4780
rect 21683 4777 21695 4811
rect 21637 4771 21695 4777
rect 22097 4811 22155 4817
rect 22097 4777 22109 4811
rect 22143 4808 22155 4811
rect 22554 4808 22560 4820
rect 22143 4780 22560 4808
rect 22143 4777 22155 4780
rect 22097 4771 22155 4777
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 24670 4808 24676 4820
rect 24631 4780 24676 4808
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 25041 4811 25099 4817
rect 25041 4777 25053 4811
rect 25087 4808 25099 4811
rect 25406 4808 25412 4820
rect 25087 4780 25412 4808
rect 25087 4777 25099 4780
rect 25041 4771 25099 4777
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 14182 4740 14188 4752
rect 14143 4712 14188 4740
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 17034 4700 17040 4752
rect 17092 4740 17098 4752
rect 17770 4740 17776 4752
rect 17092 4712 17776 4740
rect 17092 4700 17098 4712
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 19058 4700 19064 4752
rect 19116 4740 19122 4752
rect 19245 4743 19303 4749
rect 19245 4740 19257 4743
rect 19116 4712 19257 4740
rect 19116 4700 19122 4712
rect 19245 4709 19257 4712
rect 19291 4740 19303 4743
rect 20349 4743 20407 4749
rect 20349 4740 20361 4743
rect 19291 4712 20361 4740
rect 19291 4709 19303 4712
rect 19245 4703 19303 4709
rect 20349 4709 20361 4712
rect 20395 4709 20407 4743
rect 20349 4703 20407 4709
rect 12802 4672 12808 4684
rect 12763 4644 12808 4672
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 14550 4672 14556 4684
rect 13955 4644 14556 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 17494 4632 17500 4684
rect 17552 4672 17558 4684
rect 20898 4672 20904 4684
rect 17552 4644 17908 4672
rect 20859 4644 20904 4672
rect 17552 4632 17558 4644
rect 11790 4604 11796 4616
rect 11751 4576 11796 4604
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 13449 4607 13507 4613
rect 13449 4573 13461 4607
rect 13495 4604 13507 4607
rect 13814 4604 13820 4616
rect 13495 4576 13820 4604
rect 13495 4573 13507 4576
rect 13449 4567 13507 4573
rect 13814 4564 13820 4576
rect 13872 4604 13878 4616
rect 15286 4604 15292 4616
rect 13872 4576 15292 4604
rect 13872 4564 13878 4576
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 16114 4604 16120 4616
rect 16075 4576 16120 4604
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 17880 4613 17908 4644
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 22732 4675 22790 4681
rect 22732 4641 22744 4675
rect 22778 4672 22790 4675
rect 23014 4672 23020 4684
rect 22778 4644 23020 4672
rect 22778 4641 22790 4644
rect 22732 4635 22790 4641
rect 23014 4632 23020 4644
rect 23072 4632 23078 4684
rect 25133 4675 25191 4681
rect 25133 4641 25145 4675
rect 25179 4672 25191 4675
rect 25314 4672 25320 4684
rect 25179 4644 25320 4672
rect 25179 4641 25191 4644
rect 25133 4635 25191 4641
rect 25314 4632 25320 4644
rect 25372 4632 25378 4684
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 18414 4564 18420 4616
rect 18472 4604 18478 4616
rect 19337 4607 19395 4613
rect 19337 4604 19349 4607
rect 18472 4576 19349 4604
rect 18472 4564 18478 4576
rect 19337 4573 19349 4576
rect 19383 4573 19395 4607
rect 19337 4567 19395 4573
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 19981 4607 20039 4613
rect 19981 4604 19993 4607
rect 19484 4576 19993 4604
rect 19484 4564 19490 4576
rect 19981 4573 19993 4576
rect 20027 4604 20039 4607
rect 20162 4604 20168 4616
rect 20027 4576 20168 4604
rect 20027 4573 20039 4576
rect 19981 4567 20039 4573
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 21082 4604 21088 4616
rect 21043 4576 21088 4604
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 22094 4564 22100 4616
rect 22152 4604 22158 4616
rect 22465 4607 22523 4613
rect 22465 4604 22477 4607
rect 22152 4576 22477 4604
rect 22152 4564 22158 4576
rect 22465 4573 22477 4576
rect 22511 4573 22523 4607
rect 22465 4567 22523 4573
rect 25038 4564 25044 4616
rect 25096 4604 25102 4616
rect 25225 4607 25283 4613
rect 25225 4604 25237 4607
rect 25096 4576 25237 4604
rect 25096 4564 25102 4576
rect 25225 4573 25237 4576
rect 25271 4573 25283 4607
rect 25225 4567 25283 4573
rect 16206 4496 16212 4548
rect 16264 4536 16270 4548
rect 24489 4539 24547 4545
rect 24489 4536 24501 4539
rect 16264 4508 17632 4536
rect 16264 4496 16270 4508
rect 17604 4480 17632 4508
rect 23860 4508 24501 4536
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15565 4471 15623 4477
rect 15565 4468 15577 4471
rect 14608 4440 15577 4468
rect 14608 4428 14614 4440
rect 15565 4437 15577 4440
rect 15611 4437 15623 4471
rect 17126 4468 17132 4480
rect 17087 4440 17132 4468
rect 15565 4431 15623 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 17586 4428 17592 4480
rect 17644 4468 17650 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 17644 4440 18429 4468
rect 17644 4428 17650 4440
rect 18417 4437 18429 4440
rect 18463 4468 18475 4471
rect 18782 4468 18788 4480
rect 18463 4440 18788 4468
rect 18463 4437 18475 4440
rect 18417 4431 18475 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 23750 4428 23756 4480
rect 23808 4468 23814 4480
rect 23860 4477 23888 4508
rect 24489 4505 24501 4508
rect 24535 4505 24547 4539
rect 24489 4499 24547 4505
rect 23845 4471 23903 4477
rect 23845 4468 23857 4471
rect 23808 4440 23857 4468
rect 23808 4428 23814 4440
rect 23845 4437 23857 4440
rect 23891 4437 23903 4471
rect 24118 4468 24124 4480
rect 24079 4440 24124 4468
rect 23845 4431 23903 4437
rect 24118 4428 24124 4440
rect 24176 4428 24182 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 14369 4267 14427 4273
rect 14369 4233 14381 4267
rect 14415 4264 14427 4267
rect 14550 4264 14556 4276
rect 14415 4236 14556 4264
rect 14415 4233 14427 4236
rect 14369 4227 14427 4233
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 15654 4264 15660 4276
rect 15615 4236 15660 4264
rect 15654 4224 15660 4236
rect 15712 4224 15718 4276
rect 17405 4267 17463 4273
rect 17405 4233 17417 4267
rect 17451 4264 17463 4267
rect 17678 4264 17684 4276
rect 17451 4236 17684 4264
rect 17451 4233 17463 4236
rect 17405 4227 17463 4233
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 17770 4224 17776 4276
rect 17828 4264 17834 4276
rect 18509 4267 18567 4273
rect 17828 4236 17873 4264
rect 17828 4224 17834 4236
rect 18509 4233 18521 4267
rect 18555 4264 18567 4267
rect 18874 4264 18880 4276
rect 18555 4236 18880 4264
rect 18555 4233 18567 4236
rect 18509 4227 18567 4233
rect 18874 4224 18880 4236
rect 18932 4224 18938 4276
rect 19426 4264 19432 4276
rect 19387 4236 19432 4264
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 20898 4264 20904 4276
rect 20859 4236 20904 4264
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 22830 4264 22836 4276
rect 21376 4236 22836 4264
rect 12802 4196 12808 4208
rect 12360 4168 12808 4196
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12360 4128 12388 4168
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 16114 4196 16120 4208
rect 15120 4168 16120 4196
rect 12299 4100 12388 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13596 4100 13737 4128
rect 13596 4088 13602 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 14458 4128 14464 4140
rect 13955 4100 14464 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 12805 4063 12863 4069
rect 11287 4032 11928 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11900 3936 11928 4032
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13924 4060 13952 4091
rect 14458 4088 14464 4100
rect 14516 4088 14522 4140
rect 14829 4131 14887 4137
rect 14829 4097 14841 4131
rect 14875 4128 14887 4131
rect 15120 4128 15148 4168
rect 16114 4156 16120 4168
rect 16172 4156 16178 4208
rect 17037 4199 17095 4205
rect 17037 4165 17049 4199
rect 17083 4196 17095 4199
rect 17494 4196 17500 4208
rect 17083 4168 17500 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 17494 4156 17500 4168
rect 17552 4156 17558 4208
rect 19889 4199 19947 4205
rect 19889 4165 19901 4199
rect 19935 4196 19947 4199
rect 21376 4196 21404 4236
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 23474 4264 23480 4276
rect 23387 4236 23480 4264
rect 23474 4224 23480 4236
rect 23532 4264 23538 4276
rect 25038 4264 25044 4276
rect 23532 4236 24256 4264
rect 24999 4236 25044 4264
rect 23532 4224 23538 4236
rect 23750 4196 23756 4208
rect 19935 4168 21404 4196
rect 22112 4168 23756 4196
rect 19935 4165 19947 4168
rect 19889 4159 19947 4165
rect 14875 4100 15148 4128
rect 15197 4131 15255 4137
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 15378 4128 15384 4140
rect 15243 4100 15384 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16206 4128 16212 4140
rect 15528 4100 16212 4128
rect 15528 4088 15534 4100
rect 16206 4088 16212 4100
rect 16264 4088 16270 4140
rect 19702 4128 19708 4140
rect 19663 4100 19708 4128
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 20254 4088 20260 4140
rect 20312 4128 20318 4140
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 20312 4100 20453 4128
rect 20312 4088 20318 4100
rect 20441 4097 20453 4100
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 21545 4131 21603 4137
rect 21545 4097 21557 4131
rect 21591 4128 21603 4131
rect 22112 4128 22140 4168
rect 22572 4137 22600 4168
rect 23750 4156 23756 4168
rect 23808 4156 23814 4208
rect 21591 4100 22140 4128
rect 22557 4131 22615 4137
rect 21591 4097 21603 4100
rect 21545 4091 21603 4097
rect 22557 4097 22569 4131
rect 22603 4097 22615 4131
rect 22557 4091 22615 4097
rect 23842 4088 23848 4140
rect 23900 4128 23906 4140
rect 24228 4137 24256 4236
rect 25038 4224 25044 4236
rect 25096 4224 25102 4276
rect 25406 4196 25412 4208
rect 24872 4168 25412 4196
rect 24121 4131 24179 4137
rect 24121 4128 24133 4131
rect 23900 4100 24133 4128
rect 23900 4088 23906 4100
rect 24121 4097 24133 4100
rect 24167 4097 24179 4131
rect 24121 4091 24179 4097
rect 24213 4131 24271 4137
rect 24213 4097 24225 4131
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 24765 4131 24823 4137
rect 24765 4097 24777 4131
rect 24811 4128 24823 4131
rect 24872 4128 24900 4168
rect 25406 4156 25412 4168
rect 25464 4156 25470 4208
rect 24811 4100 24900 4128
rect 24811 4097 24823 4100
rect 24765 4091 24823 4097
rect 12851 4032 13952 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13633 3995 13691 4001
rect 13633 3992 13645 3995
rect 13096 3964 13645 3992
rect 13096 3936 13124 3964
rect 13633 3961 13645 3964
rect 13679 3961 13691 3995
rect 15396 3992 15424 4088
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 15611 4032 16129 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 16117 4029 16129 4032
rect 16163 4060 16175 4063
rect 16298 4060 16304 4072
rect 16163 4032 16304 4060
rect 16163 4029 16175 4032
rect 16117 4023 16175 4029
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 18598 4060 18604 4072
rect 18559 4032 18604 4060
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 16025 3995 16083 4001
rect 16025 3992 16037 3995
rect 15396 3964 16037 3992
rect 13633 3955 13691 3961
rect 16025 3961 16037 3964
rect 16071 3961 16083 3995
rect 18874 3992 18880 4004
rect 18835 3964 18880 3992
rect 16025 3955 16083 3961
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 19720 3992 19748 4088
rect 23566 4020 23572 4072
rect 23624 4060 23630 4072
rect 23750 4060 23756 4072
rect 23624 4032 23756 4060
rect 23624 4020 23630 4032
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 25222 4060 25228 4072
rect 25183 4032 25228 4060
rect 25222 4020 25228 4032
rect 25280 4060 25286 4072
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 25280 4032 25789 4060
rect 25280 4020 25286 4032
rect 25777 4029 25789 4032
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 20257 3995 20315 4001
rect 20257 3992 20269 3995
rect 19720 3964 20269 3992
rect 20257 3961 20269 3964
rect 20303 3961 20315 3995
rect 21818 3992 21824 4004
rect 21779 3964 21824 3992
rect 20257 3955 20315 3961
rect 21818 3952 21824 3964
rect 21876 3992 21882 4004
rect 22373 3995 22431 4001
rect 22373 3992 22385 3995
rect 21876 3964 22385 3992
rect 21876 3952 21882 3964
rect 22373 3961 22385 3964
rect 22419 3961 22431 3995
rect 22373 3955 22431 3961
rect 22465 3995 22523 4001
rect 22465 3961 22477 3995
rect 22511 3992 22523 3995
rect 22554 3992 22560 4004
rect 22511 3964 22560 3992
rect 22511 3961 22523 3964
rect 22465 3955 22523 3961
rect 22554 3952 22560 3964
rect 22612 3952 22618 4004
rect 24029 3995 24087 4001
rect 24029 3961 24041 3995
rect 24075 3992 24087 3995
rect 24210 3992 24216 4004
rect 24075 3964 24216 3992
rect 24075 3961 24087 3964
rect 24029 3955 24087 3961
rect 24210 3952 24216 3964
rect 24268 3952 24274 4004
rect 26142 3992 26148 4004
rect 25424 3964 26148 3992
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 13078 3924 13084 3936
rect 13039 3896 13084 3924
rect 13078 3884 13084 3896
rect 13136 3884 13142 3936
rect 13262 3924 13268 3936
rect 13223 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 22002 3924 22008 3936
rect 20404 3896 20449 3924
rect 21963 3896 22008 3924
rect 20404 3884 20410 3896
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 23014 3924 23020 3936
rect 22975 3896 23020 3924
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23474 3884 23480 3936
rect 23532 3924 23538 3936
rect 25424 3933 25452 3964
rect 26142 3952 26148 3964
rect 26200 3952 26206 4004
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 23532 3896 23673 3924
rect 23532 3884 23538 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 23661 3887 23719 3893
rect 25409 3927 25467 3933
rect 25409 3893 25421 3927
rect 25455 3893 25467 3927
rect 25409 3887 25467 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 13320 3692 14105 3720
rect 13320 3680 13326 3692
rect 14093 3689 14105 3692
rect 14139 3720 14151 3723
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14139 3692 14657 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 16393 3723 16451 3729
rect 16393 3720 16405 3723
rect 16080 3692 16405 3720
rect 16080 3680 16086 3692
rect 16393 3689 16405 3692
rect 16439 3689 16451 3723
rect 16393 3683 16451 3689
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 18414 3720 18420 3732
rect 18371 3692 18420 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 18598 3720 18604 3732
rect 18559 3692 18604 3720
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 19245 3723 19303 3729
rect 19245 3689 19257 3723
rect 19291 3720 19303 3723
rect 20346 3720 20352 3732
rect 19291 3692 20352 3720
rect 19291 3689 19303 3692
rect 19245 3683 19303 3689
rect 20346 3680 20352 3692
rect 20404 3720 20410 3732
rect 21085 3723 21143 3729
rect 21085 3720 21097 3723
rect 20404 3692 21097 3720
rect 20404 3680 20410 3692
rect 21085 3689 21097 3692
rect 21131 3689 21143 3723
rect 21085 3683 21143 3689
rect 23753 3723 23811 3729
rect 23753 3689 23765 3723
rect 23799 3720 23811 3723
rect 23842 3720 23848 3732
rect 23799 3692 23848 3720
rect 23799 3689 23811 3692
rect 23753 3683 23811 3689
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 24949 3723 25007 3729
rect 24949 3720 24961 3723
rect 24268 3692 24961 3720
rect 24268 3680 24274 3692
rect 24949 3689 24961 3692
rect 24995 3689 25007 3723
rect 25314 3720 25320 3732
rect 25275 3692 25320 3720
rect 24949 3683 25007 3689
rect 25314 3680 25320 3692
rect 25372 3680 25378 3732
rect 12250 3652 12256 3664
rect 11256 3624 12256 3652
rect 11256 3593 11284 3624
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 12618 3652 12624 3664
rect 12579 3624 12624 3652
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 13170 3612 13176 3664
rect 13228 3652 13234 3664
rect 14001 3655 14059 3661
rect 14001 3652 14013 3655
rect 13228 3624 14013 3652
rect 13228 3612 13234 3624
rect 14001 3621 14013 3624
rect 14047 3621 14059 3655
rect 15562 3652 15568 3664
rect 15523 3624 15568 3652
rect 14001 3615 14059 3621
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 16117 3655 16175 3661
rect 16117 3621 16129 3655
rect 16163 3652 16175 3655
rect 16206 3652 16212 3664
rect 16163 3624 16212 3652
rect 16163 3621 16175 3624
rect 16117 3615 16175 3621
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 17126 3652 17132 3664
rect 16592 3624 17132 3652
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3553 11299 3587
rect 12342 3584 12348 3596
rect 12303 3556 12348 3584
rect 11241 3547 11299 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3584 13415 3587
rect 13538 3584 13544 3596
rect 13403 3556 13544 3584
rect 13403 3553 13415 3556
rect 13357 3547 13415 3553
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15151 3556 15301 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15289 3553 15301 3556
rect 15335 3584 15347 3587
rect 15470 3584 15476 3596
rect 15335 3556 15476 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 16592 3593 16620 3624
rect 17126 3612 17132 3624
rect 17184 3652 17190 3664
rect 18138 3652 18144 3664
rect 17184 3624 18144 3652
rect 17184 3612 17190 3624
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 23290 3612 23296 3664
rect 23348 3652 23354 3664
rect 24305 3655 24363 3661
rect 24305 3652 24317 3655
rect 23348 3624 24317 3652
rect 23348 3612 23354 3624
rect 23860 3596 23888 3624
rect 24305 3621 24317 3624
rect 24351 3621 24363 3655
rect 24305 3615 24363 3621
rect 16850 3593 16856 3596
rect 16577 3587 16635 3593
rect 16577 3553 16589 3587
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 16844 3547 16856 3593
rect 16908 3584 16914 3596
rect 19610 3584 19616 3596
rect 16908 3556 16944 3584
rect 19571 3556 19616 3584
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8202 3516 8208 3528
rect 7800 3488 8208 3516
rect 7800 3476 7806 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10870 3516 10876 3528
rect 10275 3488 10876 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 14182 3516 14188 3528
rect 14143 3488 14188 3516
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 11422 3448 11428 3460
rect 11383 3420 11428 3448
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 12986 3408 12992 3460
rect 13044 3448 13050 3460
rect 13633 3451 13691 3457
rect 13633 3448 13645 3451
rect 13044 3420 13645 3448
rect 13044 3408 13050 3420
rect 13633 3417 13645 3420
rect 13679 3417 13691 3451
rect 13633 3411 13691 3417
rect 15470 3408 15476 3460
rect 15528 3448 15534 3460
rect 16592 3448 16620 3547
rect 16850 3544 16856 3547
rect 16908 3544 16914 3556
rect 19610 3544 19616 3556
rect 19668 3544 19674 3596
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3584 19763 3587
rect 20346 3584 20352 3596
rect 19751 3556 20352 3584
rect 19751 3553 19763 3556
rect 19705 3547 19763 3553
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 22002 3593 22008 3596
rect 21996 3584 22008 3593
rect 21963 3556 22008 3584
rect 21996 3547 22008 3556
rect 22002 3544 22008 3547
rect 22060 3544 22066 3596
rect 23842 3544 23848 3596
rect 23900 3544 23906 3596
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3485 19855 3519
rect 21726 3516 21732 3528
rect 21687 3488 21732 3516
rect 19797 3479 19855 3485
rect 19812 3448 19840 3479
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 23164 3488 24409 3516
rect 23164 3476 23170 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 24670 3516 24676 3528
rect 24627 3488 24676 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 15528 3420 16620 3448
rect 19168 3420 19840 3448
rect 15528 3408 15534 3420
rect 19168 3392 19196 3420
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 24596 3448 24624 3479
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 23072 3420 24624 3448
rect 23072 3408 23078 3420
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12618 3380 12624 3392
rect 12299 3352 12624 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12618 3340 12624 3352
rect 12676 3380 12682 3392
rect 13262 3380 13268 3392
rect 12676 3352 13268 3380
rect 12676 3340 12682 3352
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 17957 3383 18015 3389
rect 17957 3380 17969 3383
rect 17920 3352 17969 3380
rect 17920 3340 17926 3352
rect 17957 3349 17969 3352
rect 18003 3349 18015 3383
rect 19150 3380 19156 3392
rect 19111 3352 19156 3380
rect 17957 3343 18015 3349
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 20254 3380 20260 3392
rect 20215 3352 20260 3380
rect 20254 3340 20260 3352
rect 20312 3380 20318 3392
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 20312 3352 20637 3380
rect 20312 3340 20318 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 21542 3380 21548 3392
rect 21455 3352 21548 3380
rect 20625 3343 20683 3349
rect 21542 3340 21548 3352
rect 21600 3380 21606 3392
rect 22370 3380 22376 3392
rect 21600 3352 22376 3380
rect 21600 3340 21606 3352
rect 22370 3340 22376 3352
rect 22428 3340 22434 3392
rect 23124 3389 23152 3420
rect 23109 3383 23167 3389
rect 23109 3349 23121 3383
rect 23155 3349 23167 3383
rect 23109 3343 23167 3349
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3380 23995 3383
rect 24946 3380 24952 3392
rect 23983 3352 24952 3380
rect 23983 3349 23995 3352
rect 23937 3343 23995 3349
rect 24946 3340 24952 3352
rect 25004 3340 25010 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 10008 3148 10701 3176
rect 10008 3136 10014 3148
rect 10152 2981 10180 3148
rect 10689 3145 10701 3148
rect 10735 3145 10747 3179
rect 10689 3139 10747 3145
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12342 3176 12348 3188
rect 12299 3148 12348 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12805 3179 12863 3185
rect 12805 3145 12817 3179
rect 12851 3176 12863 3179
rect 14182 3176 14188 3188
rect 12851 3148 14188 3176
rect 12851 3145 12863 3148
rect 12805 3139 12863 3145
rect 14182 3136 14188 3148
rect 14240 3176 14246 3188
rect 14645 3179 14703 3185
rect 14645 3176 14657 3179
rect 14240 3148 14657 3176
rect 14240 3136 14246 3148
rect 14645 3145 14657 3148
rect 14691 3176 14703 3179
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 14691 3148 15301 3176
rect 14691 3145 14703 3148
rect 14645 3139 14703 3145
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 15289 3139 15347 3145
rect 10321 3111 10379 3117
rect 10321 3077 10333 3111
rect 10367 3108 10379 3111
rect 10962 3108 10968 3120
rect 10367 3080 10968 3108
rect 10367 3077 10379 3080
rect 10321 3071 10379 3077
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 13170 3108 13176 3120
rect 13131 3080 13176 3108
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 14458 3068 14464 3120
rect 14516 3108 14522 3120
rect 14921 3111 14979 3117
rect 14921 3108 14933 3111
rect 14516 3080 14933 3108
rect 14516 3068 14522 3080
rect 14921 3077 14933 3080
rect 14967 3077 14979 3111
rect 14921 3071 14979 3077
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12250 3040 12256 3052
rect 11931 3012 12256 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2941 10195 2975
rect 10137 2935 10195 2941
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11195 2944 11253 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11241 2941 11253 2944
rect 11287 2972 11299 2975
rect 12342 2972 12348 2984
rect 11287 2944 12348 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 13262 2972 13268 2984
rect 13175 2944 13268 2972
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13532 2975 13590 2981
rect 13532 2941 13544 2975
rect 13578 2972 13590 2975
rect 14476 2972 14504 3068
rect 15304 3040 15332 3139
rect 16850 3136 16856 3148
rect 16908 3176 16914 3188
rect 17129 3179 17187 3185
rect 17129 3176 17141 3179
rect 16908 3148 17141 3176
rect 16908 3136 16914 3148
rect 17129 3145 17141 3148
rect 17175 3145 17187 3179
rect 17862 3176 17868 3188
rect 17823 3148 17868 3176
rect 17129 3139 17187 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 19150 3136 19156 3188
rect 19208 3176 19214 3188
rect 19521 3179 19579 3185
rect 19521 3176 19533 3179
rect 19208 3148 19533 3176
rect 19208 3136 19214 3148
rect 19521 3145 19533 3148
rect 19567 3145 19579 3179
rect 19521 3139 19579 3145
rect 19610 3136 19616 3188
rect 19668 3176 19674 3188
rect 19797 3179 19855 3185
rect 19797 3176 19809 3179
rect 19668 3148 19809 3176
rect 19668 3136 19674 3148
rect 19797 3145 19809 3148
rect 19843 3145 19855 3179
rect 19797 3139 19855 3145
rect 21913 3179 21971 3185
rect 21913 3145 21925 3179
rect 21959 3176 21971 3179
rect 22002 3176 22008 3188
rect 21959 3148 22008 3176
rect 21959 3145 21971 3148
rect 21913 3139 21971 3145
rect 22002 3136 22008 3148
rect 22060 3176 22066 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 22060 3148 22201 3176
rect 22060 3136 22066 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 22189 3139 22247 3145
rect 22370 3136 22376 3188
rect 22428 3176 22434 3188
rect 22557 3179 22615 3185
rect 22557 3176 22569 3179
rect 22428 3148 22569 3176
rect 22428 3136 22434 3148
rect 22557 3145 22569 3148
rect 22603 3145 22615 3179
rect 23106 3176 23112 3188
rect 23067 3148 23112 3176
rect 22557 3139 22615 3145
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 23474 3176 23480 3188
rect 23435 3148 23480 3176
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 23842 3136 23848 3188
rect 23900 3176 23906 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 23900 3148 24409 3176
rect 23900 3136 23906 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 24397 3139 24455 3145
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 24765 3179 24823 3185
rect 24765 3176 24777 3179
rect 24728 3148 24777 3176
rect 24728 3136 24734 3148
rect 24765 3145 24777 3148
rect 24811 3145 24823 3179
rect 24765 3139 24823 3145
rect 21818 3068 21824 3120
rect 21876 3108 21882 3120
rect 23124 3108 23152 3136
rect 21876 3080 23152 3108
rect 21876 3068 21882 3080
rect 18138 3040 18144 3052
rect 15304 3012 15608 3040
rect 18099 3012 18144 3040
rect 15470 2972 15476 2984
rect 13578 2944 14504 2972
rect 15431 2944 15476 2972
rect 13578 2941 13590 2944
rect 13532 2935 13590 2941
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 15580 2972 15608 3012
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 20257 3043 20315 3049
rect 20257 3009 20269 3043
rect 20303 3040 20315 3043
rect 20346 3040 20352 3052
rect 20303 3012 20352 3040
rect 20303 3009 20315 3012
rect 20257 3003 20315 3009
rect 20346 3000 20352 3012
rect 20404 3000 20410 3052
rect 15729 2975 15787 2981
rect 15729 2972 15741 2975
rect 15580 2944 15741 2972
rect 15729 2941 15741 2944
rect 15775 2941 15787 2975
rect 15729 2935 15787 2941
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 19392 2944 20545 2972
rect 19392 2932 19398 2944
rect 20533 2941 20545 2944
rect 20579 2972 20591 2975
rect 21726 2972 21732 2984
rect 20579 2944 21732 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 21726 2932 21732 2944
rect 21784 2932 21790 2984
rect 23492 2972 23520 3136
rect 25133 3111 25191 3117
rect 25133 3077 25145 3111
rect 25179 3108 25191 3111
rect 26878 3108 26884 3120
rect 25179 3080 26884 3108
rect 25179 3077 25191 3080
rect 25133 3071 25191 3077
rect 26878 3068 26884 3080
rect 26936 3068 26942 3120
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23492 2944 23673 2972
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 24949 2975 25007 2981
rect 24949 2972 24961 2975
rect 24912 2944 24961 2972
rect 24912 2932 24918 2944
rect 24949 2941 24961 2944
rect 24995 2972 25007 2975
rect 25501 2975 25559 2981
rect 25501 2972 25513 2975
rect 24995 2944 25513 2972
rect 24995 2941 25007 2944
rect 24949 2935 25007 2941
rect 25501 2941 25513 2944
rect 25547 2941 25559 2975
rect 25501 2935 25559 2941
rect 13280 2904 13308 2932
rect 15488 2904 15516 2932
rect 13280 2876 15516 2904
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 18386 2907 18444 2913
rect 18386 2904 18398 2907
rect 17828 2876 18398 2904
rect 17828 2864 17834 2876
rect 18386 2873 18398 2876
rect 18432 2873 18444 2907
rect 18386 2867 18444 2873
rect 20254 2864 20260 2916
rect 20312 2904 20318 2916
rect 20778 2907 20836 2913
rect 20778 2904 20790 2907
rect 20312 2876 20790 2904
rect 20312 2864 20318 2876
rect 20778 2873 20790 2876
rect 20824 2873 20836 2907
rect 20778 2867 20836 2873
rect 23382 2864 23388 2916
rect 23440 2904 23446 2916
rect 23937 2907 23995 2913
rect 23937 2904 23949 2907
rect 23440 2876 23949 2904
rect 23440 2864 23446 2876
rect 23937 2873 23949 2876
rect 23983 2873 23995 2907
rect 23937 2867 23995 2873
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 17402 2836 17408 2848
rect 14976 2808 17408 2836
rect 14976 2796 14982 2808
rect 17402 2796 17408 2808
rect 17460 2796 17466 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 10962 2632 10968 2644
rect 10923 2604 10968 2632
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12618 2632 12624 2644
rect 12483 2604 12624 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13081 2635 13139 2641
rect 13081 2601 13093 2635
rect 13127 2632 13139 2635
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 13127 2604 13369 2632
rect 13127 2601 13139 2604
rect 13081 2595 13139 2601
rect 13357 2601 13369 2604
rect 13403 2632 13415 2635
rect 13630 2632 13636 2644
rect 13403 2604 13636 2632
rect 13403 2601 13415 2604
rect 13357 2595 13415 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14918 2632 14924 2644
rect 14323 2604 14924 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 16577 2635 16635 2641
rect 16577 2601 16589 2635
rect 16623 2632 16635 2635
rect 16666 2632 16672 2644
rect 16623 2604 16672 2632
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 16666 2592 16672 2604
rect 16724 2632 16730 2644
rect 17037 2635 17095 2641
rect 17037 2632 17049 2635
rect 16724 2604 17049 2632
rect 16724 2592 16730 2604
rect 17037 2601 17049 2604
rect 17083 2601 17095 2635
rect 17770 2632 17776 2644
rect 17731 2604 17776 2632
rect 17037 2595 17095 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 20254 2632 20260 2644
rect 20215 2604 20260 2632
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 20533 2635 20591 2641
rect 20533 2632 20545 2635
rect 20496 2604 20545 2632
rect 20496 2592 20502 2604
rect 20533 2601 20545 2604
rect 20579 2601 20591 2635
rect 20533 2595 20591 2601
rect 21453 2635 21511 2641
rect 21453 2601 21465 2635
rect 21499 2632 21511 2635
rect 21818 2632 21824 2644
rect 21499 2604 21824 2632
rect 21499 2601 21511 2604
rect 21453 2595 21511 2601
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 9214 2496 9220 2508
rect 8619 2468 9220 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10980 2496 11008 2592
rect 17586 2564 17592 2576
rect 11992 2536 17592 2564
rect 11992 2505 12020 2536
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 19242 2564 19248 2576
rect 18892 2536 19248 2564
rect 10367 2468 11008 2496
rect 11425 2499 11483 2505
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11471 2468 11989 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12713 2499 12771 2505
rect 12713 2465 12725 2499
rect 12759 2496 12771 2499
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 12759 2468 13093 2496
rect 12759 2465 12771 2468
rect 12713 2459 12771 2465
rect 13081 2465 13093 2468
rect 13127 2465 13139 2499
rect 13081 2459 13139 2465
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13688 2468 14197 2496
rect 13688 2456 13694 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 15562 2496 15568 2508
rect 15523 2468 15568 2496
rect 14185 2459 14243 2465
rect 15562 2456 15568 2468
rect 15620 2496 15626 2508
rect 18892 2505 18920 2536
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 20548 2564 20576 2595
rect 21818 2592 21824 2604
rect 21876 2592 21882 2644
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 22833 2635 22891 2641
rect 22833 2632 22845 2635
rect 22152 2604 22845 2632
rect 22152 2592 22158 2604
rect 22833 2601 22845 2604
rect 22879 2632 22891 2635
rect 23201 2635 23259 2641
rect 23201 2632 23213 2635
rect 22879 2604 23213 2632
rect 22879 2601 22891 2604
rect 22833 2595 22891 2601
rect 23201 2601 23213 2604
rect 23247 2632 23259 2635
rect 23569 2635 23627 2641
rect 23569 2632 23581 2635
rect 23247 2604 23581 2632
rect 23247 2601 23259 2604
rect 23201 2595 23259 2601
rect 23569 2601 23581 2604
rect 23615 2601 23627 2635
rect 23569 2595 23627 2601
rect 21910 2564 21916 2576
rect 20548 2536 21916 2564
rect 21910 2524 21916 2536
rect 21968 2524 21974 2576
rect 24305 2567 24363 2573
rect 24305 2533 24317 2567
rect 24351 2564 24363 2567
rect 24670 2564 24676 2576
rect 24351 2536 24676 2564
rect 24351 2533 24363 2536
rect 24305 2527 24363 2533
rect 24670 2524 24676 2536
rect 24728 2524 24734 2576
rect 19150 2505 19156 2508
rect 16117 2499 16175 2505
rect 16117 2496 16129 2499
rect 15620 2468 16129 2496
rect 15620 2456 15626 2468
rect 16117 2465 16129 2468
rect 16163 2465 16175 2499
rect 16117 2459 16175 2465
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2465 18935 2499
rect 19144 2496 19156 2505
rect 18877 2459 18935 2465
rect 18984 2468 19156 2496
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 15289 2431 15347 2437
rect 15289 2428 15301 2431
rect 14507 2400 15301 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 15289 2397 15301 2400
rect 15335 2428 15347 2431
rect 16758 2428 16764 2440
rect 15335 2400 16764 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2397 17187 2431
rect 17129 2391 17187 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2428 17371 2431
rect 17770 2428 17776 2440
rect 17359 2400 17776 2428
rect 17359 2397 17371 2400
rect 17313 2391 17371 2397
rect 12894 2360 12900 2372
rect 12855 2332 12900 2360
rect 12894 2320 12900 2332
rect 12952 2320 12958 2372
rect 13817 2363 13875 2369
rect 13817 2329 13829 2363
rect 13863 2360 13875 2363
rect 17144 2360 17172 2391
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 18785 2431 18843 2437
rect 18785 2397 18797 2431
rect 18831 2428 18843 2431
rect 18984 2428 19012 2468
rect 19144 2459 19156 2468
rect 19150 2456 19156 2459
rect 19208 2456 19214 2508
rect 20898 2496 20904 2508
rect 20859 2468 20904 2496
rect 20898 2456 20904 2468
rect 20956 2496 20962 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 20956 2468 21833 2496
rect 20956 2456 20962 2468
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 24029 2499 24087 2505
rect 24029 2465 24041 2499
rect 24075 2496 24087 2499
rect 24118 2496 24124 2508
rect 24075 2468 24124 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 24118 2456 24124 2468
rect 24176 2496 24182 2508
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24176 2468 24777 2496
rect 24176 2456 24182 2468
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 24765 2459 24823 2465
rect 25130 2456 25136 2508
rect 25188 2496 25194 2508
rect 25317 2499 25375 2505
rect 25317 2496 25329 2499
rect 25188 2468 25329 2496
rect 25188 2456 25194 2468
rect 25317 2465 25329 2468
rect 25363 2496 25375 2499
rect 25869 2499 25927 2505
rect 25869 2496 25881 2499
rect 25363 2468 25881 2496
rect 25363 2465 25375 2468
rect 25317 2459 25375 2465
rect 25869 2465 25881 2468
rect 25915 2465 25927 2499
rect 25869 2459 25927 2465
rect 22002 2428 22008 2440
rect 18831 2400 19012 2428
rect 21915 2400 22008 2428
rect 18831 2397 18843 2400
rect 18785 2391 18843 2397
rect 22002 2388 22008 2400
rect 22060 2428 22066 2440
rect 22465 2431 22523 2437
rect 22465 2428 22477 2431
rect 22060 2400 22477 2428
rect 22060 2388 22066 2400
rect 22465 2397 22477 2400
rect 22511 2397 22523 2431
rect 22465 2391 22523 2397
rect 18049 2363 18107 2369
rect 18049 2360 18061 2363
rect 13863 2332 18061 2360
rect 13863 2329 13875 2332
rect 13817 2323 13875 2329
rect 18049 2329 18061 2332
rect 18095 2329 18107 2363
rect 18049 2323 18107 2329
rect 25501 2363 25559 2369
rect 25501 2329 25513 2363
rect 25547 2360 25559 2363
rect 27522 2360 27528 2372
rect 25547 2332 27528 2360
rect 25547 2329 25559 2332
rect 25501 2323 25559 2329
rect 27522 2320 27528 2332
rect 27580 2320 27586 2372
rect 8754 2292 8760 2304
rect 8715 2264 8760 2292
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 10502 2292 10508 2304
rect 10463 2264 10508 2292
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 13630 2292 13636 2304
rect 13591 2264 13636 2292
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 16666 2292 16672 2304
rect 16627 2264 16672 2292
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 13906 552 13912 604
rect 13964 592 13970 604
rect 14642 592 14648 604
rect 13964 564 14648 592
rect 13964 552 13970 564
rect 14642 552 14648 564
rect 14700 552 14706 604
<< via1 >>
rect 16948 26800 17000 26852
rect 23756 26800 23808 26852
rect 21548 26596 21600 26648
rect 24768 26596 24820 26648
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 17316 25440 17368 25492
rect 22744 25440 22796 25492
rect 24676 25372 24728 25424
rect 14004 25304 14056 25356
rect 16488 25347 16540 25356
rect 16488 25313 16497 25347
rect 16497 25313 16531 25347
rect 16531 25313 16540 25347
rect 16488 25304 16540 25313
rect 19248 25304 19300 25356
rect 19984 25347 20036 25356
rect 19984 25313 19993 25347
rect 19993 25313 20027 25347
rect 20027 25313 20036 25347
rect 19984 25304 20036 25313
rect 22560 25304 22612 25356
rect 24216 25304 24268 25356
rect 18144 25236 18196 25288
rect 26148 25236 26200 25288
rect 23480 25168 23532 25220
rect 24768 25143 24820 25152
rect 24768 25109 24777 25143
rect 24777 25109 24811 25143
rect 24811 25109 24820 25143
rect 24768 25100 24820 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 21364 24896 21416 24948
rect 16028 24828 16080 24880
rect 16488 24828 16540 24880
rect 14556 24692 14608 24744
rect 14924 24667 14976 24676
rect 14924 24633 14933 24667
rect 14933 24633 14967 24667
rect 14967 24633 14976 24667
rect 14924 24624 14976 24633
rect 13452 24599 13504 24608
rect 13452 24565 13461 24599
rect 13461 24565 13495 24599
rect 13495 24565 13504 24599
rect 13452 24556 13504 24565
rect 13728 24599 13780 24608
rect 13728 24565 13737 24599
rect 13737 24565 13771 24599
rect 13771 24565 13780 24599
rect 13728 24556 13780 24565
rect 14004 24556 14056 24608
rect 16396 24556 16448 24608
rect 17316 24556 17368 24608
rect 17408 24556 17460 24608
rect 19432 24692 19484 24744
rect 20168 24692 20220 24744
rect 22192 24735 22244 24744
rect 22192 24701 22201 24735
rect 22201 24701 22235 24735
rect 22235 24701 22244 24735
rect 22192 24692 22244 24701
rect 24584 24735 24636 24744
rect 24584 24701 24593 24735
rect 24593 24701 24627 24735
rect 24627 24701 24636 24735
rect 24584 24692 24636 24701
rect 17960 24556 18012 24608
rect 19248 24556 19300 24608
rect 20076 24624 20128 24676
rect 19984 24599 20036 24608
rect 19984 24565 19993 24599
rect 19993 24565 20027 24599
rect 20027 24565 20036 24599
rect 19984 24556 20036 24565
rect 22008 24556 22060 24608
rect 22560 24599 22612 24608
rect 22560 24565 22569 24599
rect 22569 24565 22603 24599
rect 22603 24565 22612 24599
rect 22560 24556 22612 24565
rect 23112 24556 23164 24608
rect 24216 24556 24268 24608
rect 24768 24599 24820 24608
rect 24768 24565 24777 24599
rect 24777 24565 24811 24599
rect 24811 24565 24820 24599
rect 24768 24556 24820 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 12808 24395 12860 24404
rect 12808 24361 12817 24395
rect 12817 24361 12851 24395
rect 12851 24361 12860 24395
rect 12808 24352 12860 24361
rect 15108 24352 15160 24404
rect 15936 24352 15988 24404
rect 16212 24395 16264 24404
rect 16212 24361 16221 24395
rect 16221 24361 16255 24395
rect 16255 24361 16264 24395
rect 16212 24352 16264 24361
rect 18144 24395 18196 24404
rect 18144 24361 18153 24395
rect 18153 24361 18187 24395
rect 18187 24361 18196 24395
rect 18144 24352 18196 24361
rect 18696 24352 18748 24404
rect 20720 24352 20772 24404
rect 23388 24352 23440 24404
rect 23664 24395 23716 24404
rect 23664 24361 23673 24395
rect 23673 24361 23707 24395
rect 23707 24361 23716 24395
rect 23664 24352 23716 24361
rect 16672 24284 16724 24336
rect 12164 24216 12216 24268
rect 12624 24259 12676 24268
rect 12624 24225 12633 24259
rect 12633 24225 12667 24259
rect 12667 24225 12676 24259
rect 12624 24216 12676 24225
rect 13268 24216 13320 24268
rect 15752 24216 15804 24268
rect 18696 24259 18748 24268
rect 18696 24225 18705 24259
rect 18705 24225 18739 24259
rect 18739 24225 18748 24259
rect 18696 24216 18748 24225
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 22376 24259 22428 24268
rect 22376 24225 22385 24259
rect 22385 24225 22419 24259
rect 22419 24225 22428 24259
rect 22376 24216 22428 24225
rect 23480 24259 23532 24268
rect 23480 24225 23489 24259
rect 23489 24225 23523 24259
rect 23523 24225 23532 24259
rect 23480 24216 23532 24225
rect 24124 24216 24176 24268
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 20628 24148 20680 24200
rect 17868 24123 17920 24132
rect 17868 24089 17877 24123
rect 17877 24089 17911 24123
rect 17911 24089 17920 24123
rect 17868 24080 17920 24089
rect 12992 24012 13044 24064
rect 15752 24012 15804 24064
rect 18604 24055 18656 24064
rect 18604 24021 18613 24055
rect 18613 24021 18647 24055
rect 18647 24021 18656 24055
rect 18604 24012 18656 24021
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 20536 24012 20588 24064
rect 24676 24012 24728 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 12072 23808 12124 23860
rect 12624 23808 12676 23860
rect 15936 23808 15988 23860
rect 19340 23808 19392 23860
rect 21548 23851 21600 23860
rect 21548 23817 21557 23851
rect 21557 23817 21591 23851
rect 21591 23817 21600 23851
rect 21548 23808 21600 23817
rect 23296 23808 23348 23860
rect 23480 23851 23532 23860
rect 23480 23817 23489 23851
rect 23489 23817 23523 23851
rect 23523 23817 23532 23851
rect 23480 23808 23532 23817
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 16672 23672 16724 23724
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 20904 23715 20956 23724
rect 20904 23681 20913 23715
rect 20913 23681 20947 23715
rect 20947 23681 20956 23715
rect 20904 23672 20956 23681
rect 12440 23604 12492 23656
rect 14832 23604 14884 23656
rect 16212 23604 16264 23656
rect 18144 23604 18196 23656
rect 19432 23604 19484 23656
rect 20812 23604 20864 23656
rect 12072 23536 12124 23588
rect 12532 23536 12584 23588
rect 14372 23536 14424 23588
rect 15936 23536 15988 23588
rect 16120 23536 16172 23588
rect 19984 23536 20036 23588
rect 8392 23468 8444 23520
rect 9680 23468 9732 23520
rect 12808 23468 12860 23520
rect 15568 23468 15620 23520
rect 16488 23468 16540 23520
rect 17776 23511 17828 23520
rect 17776 23477 17785 23511
rect 17785 23477 17819 23511
rect 17819 23477 17828 23511
rect 17776 23468 17828 23477
rect 18052 23511 18104 23520
rect 18052 23477 18061 23511
rect 18061 23477 18095 23511
rect 18095 23477 18104 23511
rect 18052 23468 18104 23477
rect 18696 23468 18748 23520
rect 19524 23511 19576 23520
rect 19524 23477 19533 23511
rect 19533 23477 19567 23511
rect 19567 23477 19576 23511
rect 19524 23468 19576 23477
rect 22468 23468 22520 23520
rect 22652 23468 22704 23520
rect 24124 23468 24176 23520
rect 24860 23468 24912 23520
rect 25412 23468 25464 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 12440 23307 12492 23316
rect 12440 23273 12449 23307
rect 12449 23273 12483 23307
rect 12483 23273 12492 23307
rect 12440 23264 12492 23273
rect 11980 23103 12032 23112
rect 11980 23069 11989 23103
rect 11989 23069 12023 23103
rect 12023 23069 12032 23103
rect 11980 23060 12032 23069
rect 12440 23060 12492 23112
rect 14096 23264 14148 23316
rect 14832 23264 14884 23316
rect 12992 23196 13044 23248
rect 16580 23264 16632 23316
rect 20720 23264 20772 23316
rect 23388 23264 23440 23316
rect 17868 23239 17920 23248
rect 17868 23205 17902 23239
rect 17902 23205 17920 23239
rect 17868 23196 17920 23205
rect 25228 23239 25280 23248
rect 25228 23205 25237 23239
rect 25237 23205 25271 23239
rect 25271 23205 25280 23239
rect 25228 23196 25280 23205
rect 15568 23171 15620 23180
rect 15568 23137 15602 23171
rect 15602 23137 15620 23171
rect 15568 23128 15620 23137
rect 19524 23128 19576 23180
rect 21272 23128 21324 23180
rect 22836 23128 22888 23180
rect 23940 23128 23992 23180
rect 25044 23128 25096 23180
rect 20628 23060 20680 23112
rect 21364 23103 21416 23112
rect 21364 23069 21373 23103
rect 21373 23069 21407 23103
rect 21407 23069 21416 23103
rect 21364 23060 21416 23069
rect 16672 23035 16724 23044
rect 16672 23001 16681 23035
rect 16681 23001 16715 23035
rect 16715 23001 16724 23035
rect 16672 22992 16724 23001
rect 22376 23060 22428 23112
rect 14372 22967 14424 22976
rect 14372 22933 14381 22967
rect 14381 22933 14415 22967
rect 14415 22933 14424 22967
rect 14372 22924 14424 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 18880 22924 18932 22976
rect 20444 22924 20496 22976
rect 20904 22967 20956 22976
rect 20904 22933 20913 22967
rect 20913 22933 20947 22967
rect 20947 22933 20956 22967
rect 20904 22924 20956 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 14556 22720 14608 22772
rect 10876 22584 10928 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 15568 22584 15620 22636
rect 16580 22584 16632 22636
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17868 22720 17920 22772
rect 21088 22720 21140 22772
rect 21364 22720 21416 22772
rect 25044 22720 25096 22772
rect 17040 22584 17092 22593
rect 18236 22516 18288 22568
rect 24216 22584 24268 22636
rect 14188 22491 14240 22500
rect 14188 22457 14197 22491
rect 14197 22457 14231 22491
rect 14231 22457 14240 22491
rect 14188 22448 14240 22457
rect 16856 22448 16908 22500
rect 19524 22516 19576 22568
rect 21272 22516 21324 22568
rect 22836 22559 22888 22568
rect 22836 22525 22845 22559
rect 22845 22525 22879 22559
rect 22879 22525 22888 22559
rect 22836 22516 22888 22525
rect 18880 22448 18932 22500
rect 25044 22516 25096 22568
rect 12256 22423 12308 22432
rect 12256 22389 12265 22423
rect 12265 22389 12299 22423
rect 12299 22389 12308 22423
rect 12256 22380 12308 22389
rect 12992 22380 13044 22432
rect 15108 22423 15160 22432
rect 15108 22389 15117 22423
rect 15117 22389 15151 22423
rect 15151 22389 15160 22423
rect 15108 22380 15160 22389
rect 16488 22380 16540 22432
rect 19524 22380 19576 22432
rect 20444 22380 20496 22432
rect 22560 22423 22612 22432
rect 22560 22389 22569 22423
rect 22569 22389 22603 22423
rect 22603 22389 22612 22423
rect 22560 22380 22612 22389
rect 23848 22380 23900 22432
rect 24400 22423 24452 22432
rect 24400 22389 24409 22423
rect 24409 22389 24443 22423
rect 24443 22389 24452 22423
rect 24400 22380 24452 22389
rect 24860 22380 24912 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 10876 22219 10928 22228
rect 10876 22185 10885 22219
rect 10885 22185 10919 22219
rect 10919 22185 10928 22219
rect 10876 22176 10928 22185
rect 12256 22176 12308 22228
rect 12992 22219 13044 22228
rect 12992 22185 13001 22219
rect 13001 22185 13035 22219
rect 13035 22185 13044 22219
rect 12992 22176 13044 22185
rect 14648 22176 14700 22228
rect 15108 22176 15160 22228
rect 17040 22176 17092 22228
rect 18052 22219 18104 22228
rect 18052 22185 18061 22219
rect 18061 22185 18095 22219
rect 18095 22185 18104 22219
rect 18052 22176 18104 22185
rect 20720 22219 20772 22228
rect 20720 22185 20729 22219
rect 20729 22185 20763 22219
rect 20763 22185 20772 22219
rect 20720 22176 20772 22185
rect 24952 22176 25004 22228
rect 25136 22176 25188 22228
rect 1400 22040 1452 22092
rect 2320 22040 2372 22092
rect 11244 22083 11296 22092
rect 11244 22049 11278 22083
rect 11278 22049 11296 22083
rect 11244 22040 11296 22049
rect 12808 22040 12860 22092
rect 13544 22040 13596 22092
rect 14648 22083 14700 22092
rect 14648 22049 14657 22083
rect 14657 22049 14691 22083
rect 14691 22049 14700 22083
rect 14648 22040 14700 22049
rect 15292 22040 15344 22092
rect 14372 21972 14424 22024
rect 14740 21972 14792 22024
rect 15568 21972 15620 22024
rect 16488 21972 16540 22024
rect 16580 21972 16632 22024
rect 17776 21972 17828 22024
rect 19616 22083 19668 22092
rect 19616 22049 19625 22083
rect 19625 22049 19659 22083
rect 19659 22049 19668 22083
rect 19616 22040 19668 22049
rect 20904 22040 20956 22092
rect 21180 22040 21232 22092
rect 22560 22108 22612 22160
rect 23848 22083 23900 22092
rect 23848 22049 23857 22083
rect 23857 22049 23891 22083
rect 23891 22049 23900 22083
rect 23848 22040 23900 22049
rect 24768 22040 24820 22092
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 25412 22083 25464 22092
rect 25412 22049 25421 22083
rect 25421 22049 25455 22083
rect 25455 22049 25464 22083
rect 25412 22040 25464 22049
rect 18236 22015 18288 22024
rect 18236 21981 18245 22015
rect 18245 21981 18279 22015
rect 18279 21981 18288 22015
rect 18236 21972 18288 21981
rect 19708 22015 19760 22024
rect 19708 21981 19717 22015
rect 19717 21981 19751 22015
rect 19751 21981 19760 22015
rect 19708 21972 19760 21981
rect 17684 21947 17736 21956
rect 17684 21913 17693 21947
rect 17693 21913 17727 21947
rect 17727 21913 17736 21947
rect 17684 21904 17736 21913
rect 19340 21904 19392 21956
rect 19524 21904 19576 21956
rect 10692 21836 10744 21888
rect 15660 21879 15712 21888
rect 15660 21845 15669 21879
rect 15669 21845 15703 21879
rect 15703 21845 15712 21879
rect 15660 21836 15712 21845
rect 16304 21836 16356 21888
rect 18604 21836 18656 21888
rect 18880 21836 18932 21888
rect 20352 21836 20404 21888
rect 24584 21904 24636 21956
rect 21272 21836 21324 21888
rect 22560 21836 22612 21888
rect 22744 21879 22796 21888
rect 22744 21845 22753 21879
rect 22753 21845 22787 21879
rect 22787 21845 22796 21879
rect 22744 21836 22796 21845
rect 24676 21836 24728 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 9680 21632 9732 21684
rect 11244 21675 11296 21684
rect 10232 21607 10284 21616
rect 10232 21573 10241 21607
rect 10241 21573 10275 21607
rect 10275 21573 10284 21607
rect 10232 21564 10284 21573
rect 11244 21641 11253 21675
rect 11253 21641 11287 21675
rect 11287 21641 11296 21675
rect 11244 21632 11296 21641
rect 14188 21675 14240 21684
rect 14188 21641 14197 21675
rect 14197 21641 14231 21675
rect 14231 21641 14240 21675
rect 14188 21632 14240 21641
rect 15292 21675 15344 21684
rect 15292 21641 15301 21675
rect 15301 21641 15335 21675
rect 15335 21641 15344 21675
rect 15292 21632 15344 21641
rect 15568 21632 15620 21684
rect 18236 21632 18288 21684
rect 19616 21632 19668 21684
rect 23848 21675 23900 21684
rect 23848 21641 23857 21675
rect 23857 21641 23891 21675
rect 23891 21641 23900 21675
rect 23848 21632 23900 21641
rect 20444 21607 20496 21616
rect 20444 21573 20453 21607
rect 20453 21573 20487 21607
rect 20487 21573 20496 21607
rect 20444 21564 20496 21573
rect 20628 21564 20680 21616
rect 22008 21564 22060 21616
rect 25136 21607 25188 21616
rect 25136 21573 25145 21607
rect 25145 21573 25179 21607
rect 25179 21573 25188 21607
rect 25136 21564 25188 21573
rect 10692 21496 10744 21548
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 14740 21539 14792 21548
rect 14740 21505 14749 21539
rect 14749 21505 14783 21539
rect 14783 21505 14792 21539
rect 14740 21496 14792 21505
rect 15660 21496 15712 21548
rect 18880 21539 18932 21548
rect 14648 21428 14700 21480
rect 10140 21292 10192 21344
rect 10784 21292 10836 21344
rect 11060 21292 11112 21344
rect 12440 21335 12492 21344
rect 12440 21301 12449 21335
rect 12449 21301 12483 21335
rect 12483 21301 12492 21335
rect 12440 21292 12492 21301
rect 12716 21292 12768 21344
rect 13544 21292 13596 21344
rect 13820 21292 13872 21344
rect 14832 21292 14884 21344
rect 15844 21335 15896 21344
rect 15844 21301 15853 21335
rect 15853 21301 15887 21335
rect 15887 21301 15896 21335
rect 15844 21292 15896 21301
rect 16304 21292 16356 21344
rect 18880 21505 18889 21539
rect 18889 21505 18923 21539
rect 18923 21505 18932 21539
rect 18880 21496 18932 21505
rect 19524 21496 19576 21548
rect 19708 21496 19760 21548
rect 21180 21496 21232 21548
rect 22560 21539 22612 21548
rect 22560 21505 22569 21539
rect 22569 21505 22603 21539
rect 22603 21505 22612 21539
rect 22560 21496 22612 21505
rect 20904 21428 20956 21480
rect 23940 21428 23992 21480
rect 25504 21471 25556 21480
rect 25504 21437 25513 21471
rect 25513 21437 25547 21471
rect 25547 21437 25556 21471
rect 25504 21428 25556 21437
rect 18236 21360 18288 21412
rect 20996 21360 21048 21412
rect 24492 21403 24544 21412
rect 24492 21369 24501 21403
rect 24501 21369 24535 21403
rect 24535 21369 24544 21403
rect 24492 21360 24544 21369
rect 17224 21292 17276 21344
rect 18328 21335 18380 21344
rect 18328 21301 18337 21335
rect 18337 21301 18371 21335
rect 18371 21301 18380 21335
rect 18328 21292 18380 21301
rect 18604 21292 18656 21344
rect 20352 21292 20404 21344
rect 22008 21335 22060 21344
rect 22008 21301 22017 21335
rect 22017 21301 22051 21335
rect 22051 21301 22060 21335
rect 22008 21292 22060 21301
rect 22100 21292 22152 21344
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 10876 21088 10928 21140
rect 11244 21088 11296 21140
rect 12716 21131 12768 21140
rect 12716 21097 12725 21131
rect 12725 21097 12759 21131
rect 12759 21097 12768 21131
rect 12716 21088 12768 21097
rect 13176 21131 13228 21140
rect 13176 21097 13185 21131
rect 13185 21097 13219 21131
rect 13219 21097 13228 21131
rect 13176 21088 13228 21097
rect 14740 21131 14792 21140
rect 14740 21097 14749 21131
rect 14749 21097 14783 21131
rect 14783 21097 14792 21131
rect 14740 21088 14792 21097
rect 17776 21131 17828 21140
rect 17776 21097 17785 21131
rect 17785 21097 17819 21131
rect 17819 21097 17828 21131
rect 17776 21088 17828 21097
rect 19340 21131 19392 21140
rect 19340 21097 19349 21131
rect 19349 21097 19383 21131
rect 19383 21097 19392 21131
rect 19340 21088 19392 21097
rect 20076 21088 20128 21140
rect 20352 21088 20404 21140
rect 21180 21131 21232 21140
rect 21180 21097 21189 21131
rect 21189 21097 21223 21131
rect 21223 21097 21232 21131
rect 21180 21088 21232 21097
rect 24032 21131 24084 21140
rect 24032 21097 24041 21131
rect 24041 21097 24075 21131
rect 24075 21097 24084 21131
rect 24032 21088 24084 21097
rect 10692 21020 10744 21072
rect 11060 21020 11112 21072
rect 14004 21020 14056 21072
rect 14648 21020 14700 21072
rect 13084 20995 13136 21004
rect 13084 20961 13093 20995
rect 13093 20961 13127 20995
rect 13127 20961 13136 20995
rect 13084 20952 13136 20961
rect 14464 20995 14516 21004
rect 14464 20961 14473 20995
rect 14473 20961 14507 20995
rect 14507 20961 14516 20995
rect 14464 20952 14516 20961
rect 16488 20952 16540 21004
rect 17960 20952 18012 21004
rect 13268 20927 13320 20936
rect 13268 20893 13277 20927
rect 13277 20893 13311 20927
rect 13311 20893 13320 20927
rect 13268 20884 13320 20893
rect 13636 20816 13688 20868
rect 14188 20816 14240 20868
rect 15568 20816 15620 20868
rect 18144 20884 18196 20936
rect 19432 20952 19484 21004
rect 19708 20995 19760 21004
rect 19708 20961 19717 20995
rect 19717 20961 19751 20995
rect 19751 20961 19760 20995
rect 19708 20952 19760 20961
rect 21272 20952 21324 21004
rect 21732 20995 21784 21004
rect 21732 20961 21766 20995
rect 21766 20961 21784 20995
rect 21732 20952 21784 20961
rect 25228 20995 25280 21004
rect 25228 20961 25237 20995
rect 25237 20961 25271 20995
rect 25271 20961 25280 20995
rect 25228 20952 25280 20961
rect 18880 20884 18932 20936
rect 24032 20884 24084 20936
rect 24216 20927 24268 20936
rect 24216 20893 24225 20927
rect 24225 20893 24259 20927
rect 24259 20893 24268 20927
rect 24216 20884 24268 20893
rect 10692 20748 10744 20800
rect 13912 20748 13964 20800
rect 17224 20791 17276 20800
rect 17224 20757 17233 20791
rect 17233 20757 17267 20791
rect 17267 20757 17276 20791
rect 17224 20748 17276 20757
rect 18052 20791 18104 20800
rect 18052 20757 18061 20791
rect 18061 20757 18095 20791
rect 18095 20757 18104 20791
rect 18052 20748 18104 20757
rect 22376 20748 22428 20800
rect 22744 20748 22796 20800
rect 24952 20816 25004 20868
rect 24216 20748 24268 20800
rect 24768 20748 24820 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 9404 20587 9456 20596
rect 9404 20553 9413 20587
rect 9413 20553 9447 20587
rect 9447 20553 9456 20587
rect 9404 20544 9456 20553
rect 10968 20544 11020 20596
rect 11060 20544 11112 20596
rect 11520 20544 11572 20596
rect 11888 20544 11940 20596
rect 15292 20544 15344 20596
rect 16488 20544 16540 20596
rect 17868 20544 17920 20596
rect 18420 20544 18472 20596
rect 21272 20544 21324 20596
rect 22008 20587 22060 20596
rect 22008 20553 22017 20587
rect 22017 20553 22051 20587
rect 22051 20553 22060 20587
rect 22008 20544 22060 20553
rect 25044 20587 25096 20596
rect 25044 20553 25053 20587
rect 25053 20553 25087 20587
rect 25087 20553 25096 20587
rect 25044 20544 25096 20553
rect 25228 20544 25280 20596
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 11244 20408 11296 20460
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13636 20451 13688 20460
rect 13636 20417 13645 20451
rect 13645 20417 13679 20451
rect 13679 20417 13688 20451
rect 13636 20408 13688 20417
rect 15844 20408 15896 20460
rect 21916 20476 21968 20528
rect 9404 20340 9456 20392
rect 13912 20383 13964 20392
rect 13912 20349 13946 20383
rect 13946 20349 13964 20383
rect 13912 20340 13964 20349
rect 21732 20408 21784 20460
rect 22560 20451 22612 20460
rect 22560 20417 22569 20451
rect 22569 20417 22603 20451
rect 22603 20417 22612 20451
rect 22560 20408 22612 20417
rect 25412 20451 25464 20460
rect 16948 20340 17000 20392
rect 19156 20383 19208 20392
rect 9864 20204 9916 20256
rect 11244 20247 11296 20256
rect 11244 20213 11253 20247
rect 11253 20213 11287 20247
rect 11287 20213 11296 20247
rect 11244 20204 11296 20213
rect 13084 20204 13136 20256
rect 14740 20204 14792 20256
rect 14832 20204 14884 20256
rect 16580 20272 16632 20324
rect 16396 20247 16448 20256
rect 16396 20213 16405 20247
rect 16405 20213 16439 20247
rect 16439 20213 16448 20247
rect 16396 20204 16448 20213
rect 16764 20204 16816 20256
rect 18144 20204 18196 20256
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 20720 20340 20772 20392
rect 23664 20340 23716 20392
rect 25412 20417 25421 20451
rect 25421 20417 25455 20451
rect 25455 20417 25464 20451
rect 25412 20408 25464 20417
rect 24584 20340 24636 20392
rect 24952 20340 25004 20392
rect 19064 20315 19116 20324
rect 19064 20281 19073 20315
rect 19073 20281 19107 20315
rect 19107 20281 19116 20315
rect 19064 20272 19116 20281
rect 21272 20272 21324 20324
rect 22284 20272 22336 20324
rect 18788 20204 18840 20256
rect 18880 20204 18932 20256
rect 21088 20204 21140 20256
rect 22100 20204 22152 20256
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 23664 20247 23716 20256
rect 23664 20213 23673 20247
rect 23673 20213 23707 20247
rect 23707 20213 23716 20247
rect 23664 20204 23716 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 11520 20043 11572 20052
rect 11520 20009 11529 20043
rect 11529 20009 11563 20043
rect 11563 20009 11572 20043
rect 11520 20000 11572 20009
rect 13176 20000 13228 20052
rect 14464 20000 14516 20052
rect 16396 20000 16448 20052
rect 18052 20000 18104 20052
rect 18328 20000 18380 20052
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 20076 20000 20128 20052
rect 20352 20043 20404 20052
rect 20352 20009 20361 20043
rect 20361 20009 20395 20043
rect 20395 20009 20404 20043
rect 20352 20000 20404 20009
rect 20720 20043 20772 20052
rect 20720 20009 20729 20043
rect 20729 20009 20763 20043
rect 20763 20009 20772 20043
rect 20720 20000 20772 20009
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 24032 20000 24084 20052
rect 24124 20000 24176 20052
rect 24952 20000 25004 20052
rect 10876 19932 10928 19984
rect 10232 19864 10284 19916
rect 13636 19932 13688 19984
rect 25320 19932 25372 19984
rect 12808 19864 12860 19916
rect 14832 19864 14884 19916
rect 15568 19907 15620 19916
rect 15568 19873 15577 19907
rect 15577 19873 15611 19907
rect 15611 19873 15620 19907
rect 15568 19864 15620 19873
rect 15660 19864 15712 19916
rect 19708 19907 19760 19916
rect 19708 19873 19717 19907
rect 19717 19873 19751 19907
rect 19751 19873 19760 19907
rect 19708 19864 19760 19873
rect 21272 19864 21324 19916
rect 22376 19864 22428 19916
rect 24216 19864 24268 19916
rect 24952 19907 25004 19916
rect 24952 19873 24961 19907
rect 24961 19873 24995 19907
rect 24995 19873 25004 19907
rect 24952 19864 25004 19873
rect 18144 19796 18196 19848
rect 19156 19796 19208 19848
rect 22284 19839 22336 19848
rect 22284 19805 22293 19839
rect 22293 19805 22327 19839
rect 22327 19805 22336 19839
rect 22284 19796 22336 19805
rect 24584 19796 24636 19848
rect 25964 19796 26016 19848
rect 13912 19728 13964 19780
rect 16948 19771 17000 19780
rect 16948 19737 16957 19771
rect 16957 19737 16991 19771
rect 16991 19737 17000 19771
rect 16948 19728 17000 19737
rect 23480 19728 23532 19780
rect 14188 19660 14240 19712
rect 19340 19660 19392 19712
rect 22100 19703 22152 19712
rect 22100 19669 22109 19703
rect 22109 19669 22143 19703
rect 22143 19669 22152 19703
rect 22100 19660 22152 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 10876 19456 10928 19508
rect 296 19320 348 19372
rect 388 19320 440 19372
rect 12808 19456 12860 19508
rect 15292 19456 15344 19508
rect 17132 19456 17184 19508
rect 17408 19456 17460 19508
rect 18328 19456 18380 19508
rect 22376 19456 22428 19508
rect 24676 19456 24728 19508
rect 24952 19456 25004 19508
rect 25964 19499 26016 19508
rect 25964 19465 25973 19499
rect 25973 19465 26007 19499
rect 26007 19465 26016 19499
rect 25964 19456 26016 19465
rect 14740 19388 14792 19440
rect 14832 19320 14884 19372
rect 10232 19295 10284 19304
rect 10232 19261 10241 19295
rect 10241 19261 10275 19295
rect 10275 19261 10284 19295
rect 10232 19252 10284 19261
rect 14280 19252 14332 19304
rect 12624 19184 12676 19236
rect 13912 19184 13964 19236
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 16488 19320 16540 19372
rect 18880 19388 18932 19440
rect 17776 19320 17828 19372
rect 16856 19252 16908 19304
rect 17408 19252 17460 19304
rect 18144 19320 18196 19372
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 22560 19363 22612 19372
rect 22560 19329 22569 19363
rect 22569 19329 22603 19363
rect 22603 19329 22612 19363
rect 22560 19320 22612 19329
rect 22652 19320 22704 19372
rect 22836 19320 22888 19372
rect 15660 19184 15712 19236
rect 17224 19184 17276 19236
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 16304 19116 16356 19168
rect 16488 19116 16540 19168
rect 17316 19116 17368 19168
rect 18880 19116 18932 19168
rect 19708 19252 19760 19304
rect 22744 19252 22796 19304
rect 19340 19184 19392 19236
rect 22100 19184 22152 19236
rect 24032 19320 24084 19372
rect 23664 19252 23716 19304
rect 25228 19295 25280 19304
rect 25228 19261 25237 19295
rect 25237 19261 25271 19295
rect 25271 19261 25280 19295
rect 25228 19252 25280 19261
rect 25504 19227 25556 19236
rect 25504 19193 25513 19227
rect 25513 19193 25547 19227
rect 25547 19193 25556 19227
rect 25504 19184 25556 19193
rect 19064 19116 19116 19168
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 22744 19116 22796 19168
rect 24124 19116 24176 19168
rect 25320 19116 25372 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 13636 18912 13688 18964
rect 14464 18912 14516 18964
rect 15660 18955 15712 18964
rect 15660 18921 15669 18955
rect 15669 18921 15703 18955
rect 15703 18921 15712 18955
rect 15660 18912 15712 18921
rect 16580 18912 16632 18964
rect 17868 18955 17920 18964
rect 17868 18921 17877 18955
rect 17877 18921 17911 18955
rect 17911 18921 17920 18955
rect 17868 18912 17920 18921
rect 19340 18912 19392 18964
rect 19984 18912 20036 18964
rect 20720 18955 20772 18964
rect 20720 18921 20729 18955
rect 20729 18921 20763 18955
rect 20763 18921 20772 18955
rect 20720 18912 20772 18921
rect 21456 18912 21508 18964
rect 22560 18912 22612 18964
rect 23204 18912 23256 18964
rect 25228 18912 25280 18964
rect 14004 18844 14056 18896
rect 11704 18776 11756 18828
rect 12716 18776 12768 18828
rect 14740 18819 14792 18828
rect 14740 18785 14749 18819
rect 14749 18785 14783 18819
rect 14783 18785 14792 18819
rect 14740 18776 14792 18785
rect 16396 18776 16448 18828
rect 19156 18844 19208 18896
rect 25044 18844 25096 18896
rect 18512 18776 18564 18828
rect 21180 18819 21232 18828
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 22376 18776 22428 18828
rect 24032 18776 24084 18828
rect 11520 18708 11572 18760
rect 12256 18708 12308 18760
rect 11428 18683 11480 18692
rect 11428 18649 11437 18683
rect 11437 18649 11471 18683
rect 11471 18649 11480 18683
rect 11428 18640 11480 18649
rect 12624 18640 12676 18692
rect 14188 18708 14240 18760
rect 16212 18708 16264 18760
rect 22284 18751 22336 18760
rect 16488 18640 16540 18692
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 24952 18751 25004 18760
rect 24952 18717 24961 18751
rect 24961 18717 24995 18751
rect 24995 18717 25004 18751
rect 24952 18708 25004 18717
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 24216 18640 24268 18692
rect 12900 18615 12952 18624
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 13176 18572 13228 18624
rect 15568 18572 15620 18624
rect 15660 18572 15712 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 17960 18572 18012 18624
rect 20076 18615 20128 18624
rect 20076 18581 20085 18615
rect 20085 18581 20119 18615
rect 20119 18581 20128 18615
rect 20076 18572 20128 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 11336 18368 11388 18420
rect 12716 18411 12768 18420
rect 12716 18377 12725 18411
rect 12725 18377 12759 18411
rect 12759 18377 12768 18411
rect 12716 18368 12768 18377
rect 14004 18368 14056 18420
rect 14188 18411 14240 18420
rect 14188 18377 14197 18411
rect 14197 18377 14231 18411
rect 14231 18377 14240 18411
rect 14188 18368 14240 18377
rect 14556 18368 14608 18420
rect 19064 18411 19116 18420
rect 11520 18300 11572 18352
rect 11704 18300 11756 18352
rect 12440 18300 12492 18352
rect 14280 18300 14332 18352
rect 12900 18232 12952 18284
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 13820 18232 13872 18284
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 19984 18368 20036 18420
rect 22376 18411 22428 18420
rect 15568 18275 15620 18284
rect 15568 18241 15577 18275
rect 15577 18241 15611 18275
rect 15611 18241 15620 18275
rect 15568 18232 15620 18241
rect 16396 18232 16448 18284
rect 19432 18300 19484 18352
rect 20076 18300 20128 18352
rect 20260 18275 20312 18284
rect 20260 18241 20269 18275
rect 20269 18241 20303 18275
rect 20303 18241 20312 18275
rect 20260 18232 20312 18241
rect 22376 18377 22385 18411
rect 22385 18377 22419 18411
rect 22419 18377 22428 18411
rect 22376 18368 22428 18377
rect 22652 18411 22704 18420
rect 22652 18377 22661 18411
rect 22661 18377 22695 18411
rect 22695 18377 22704 18411
rect 22652 18368 22704 18377
rect 22744 18368 22796 18420
rect 24124 18368 24176 18420
rect 24952 18368 25004 18420
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 24032 18232 24084 18284
rect 11428 18207 11480 18216
rect 11428 18173 11437 18207
rect 11437 18173 11471 18207
rect 11471 18173 11480 18207
rect 11428 18164 11480 18173
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13176 18164 13228 18173
rect 16580 18207 16632 18216
rect 16580 18173 16589 18207
rect 16589 18173 16623 18207
rect 16623 18173 16632 18207
rect 16580 18164 16632 18173
rect 20076 18164 20128 18216
rect 15200 18096 15252 18148
rect 15844 18096 15896 18148
rect 16856 18139 16908 18148
rect 16856 18105 16865 18139
rect 16865 18105 16899 18139
rect 16899 18105 16908 18139
rect 16856 18096 16908 18105
rect 17960 18096 18012 18148
rect 18512 18096 18564 18148
rect 20720 18164 20772 18216
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 22744 18164 22796 18216
rect 23020 18207 23072 18216
rect 23020 18173 23029 18207
rect 23029 18173 23063 18207
rect 23063 18173 23072 18207
rect 25228 18207 25280 18216
rect 23020 18164 23072 18173
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 15108 18028 15160 18080
rect 16488 18028 16540 18080
rect 18052 18028 18104 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 19340 18028 19392 18080
rect 23020 18028 23072 18080
rect 25044 18071 25096 18080
rect 25044 18037 25053 18071
rect 25053 18037 25087 18071
rect 25087 18037 25096 18071
rect 25044 18028 25096 18037
rect 25412 18071 25464 18080
rect 25412 18037 25421 18071
rect 25421 18037 25455 18071
rect 25455 18037 25464 18071
rect 25412 18028 25464 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 12900 17824 12952 17876
rect 14648 17824 14700 17876
rect 15016 17867 15068 17876
rect 15016 17833 15025 17867
rect 15025 17833 15059 17867
rect 15059 17833 15068 17867
rect 15016 17824 15068 17833
rect 16212 17867 16264 17876
rect 16212 17833 16221 17867
rect 16221 17833 16255 17867
rect 16255 17833 16264 17867
rect 16212 17824 16264 17833
rect 17960 17867 18012 17876
rect 17960 17833 17969 17867
rect 17969 17833 18003 17867
rect 18003 17833 18012 17867
rect 17960 17824 18012 17833
rect 22100 17867 22152 17876
rect 22100 17833 22109 17867
rect 22109 17833 22143 17867
rect 22143 17833 22152 17867
rect 22100 17824 22152 17833
rect 24032 17824 24084 17876
rect 25136 17824 25188 17876
rect 14740 17756 14792 17808
rect 16580 17756 16632 17808
rect 16948 17756 17000 17808
rect 18512 17756 18564 17808
rect 11704 17731 11756 17740
rect 11704 17697 11713 17731
rect 11713 17697 11747 17731
rect 11747 17697 11756 17731
rect 11704 17688 11756 17697
rect 12348 17688 12400 17740
rect 13544 17688 13596 17740
rect 14372 17688 14424 17740
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 13452 17620 13504 17672
rect 14188 17620 14240 17672
rect 15936 17620 15988 17672
rect 17776 17688 17828 17740
rect 17960 17688 18012 17740
rect 18328 17688 18380 17740
rect 19340 17756 19392 17808
rect 20168 17756 20220 17808
rect 23204 17799 23256 17808
rect 23204 17765 23238 17799
rect 23238 17765 23256 17799
rect 23204 17756 23256 17765
rect 21272 17731 21324 17740
rect 12624 17552 12676 17604
rect 18052 17552 18104 17604
rect 19248 17595 19300 17604
rect 19248 17561 19257 17595
rect 19257 17561 19291 17595
rect 19291 17561 19300 17595
rect 19248 17552 19300 17561
rect 19984 17620 20036 17672
rect 21272 17697 21281 17731
rect 21281 17697 21315 17731
rect 21315 17697 21324 17731
rect 21272 17688 21324 17697
rect 25228 17688 25280 17740
rect 20904 17620 20956 17672
rect 21548 17620 21600 17672
rect 22928 17663 22980 17672
rect 22928 17629 22937 17663
rect 22937 17629 22971 17663
rect 22971 17629 22980 17663
rect 22928 17620 22980 17629
rect 11888 17484 11940 17536
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 18972 17527 19024 17536
rect 18972 17493 18981 17527
rect 18981 17493 19015 17527
rect 19015 17493 19024 17527
rect 18972 17484 19024 17493
rect 22468 17527 22520 17536
rect 22468 17493 22477 17527
rect 22477 17493 22511 17527
rect 22511 17493 22520 17527
rect 22468 17484 22520 17493
rect 25320 17527 25372 17536
rect 25320 17493 25329 17527
rect 25329 17493 25363 17527
rect 25363 17493 25372 17527
rect 25320 17484 25372 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 11704 17280 11756 17332
rect 14188 17323 14240 17332
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 19984 17280 20036 17332
rect 21272 17280 21324 17332
rect 23204 17280 23256 17332
rect 14648 17255 14700 17264
rect 11612 17144 11664 17196
rect 11980 17076 12032 17128
rect 14648 17221 14657 17255
rect 14657 17221 14691 17255
rect 14691 17221 14700 17255
rect 14648 17212 14700 17221
rect 14464 17076 14516 17128
rect 14832 17119 14884 17128
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 21916 17212 21968 17264
rect 25320 17255 25372 17264
rect 25320 17221 25329 17255
rect 25329 17221 25363 17255
rect 25363 17221 25372 17255
rect 25320 17212 25372 17221
rect 18236 17144 18288 17196
rect 19984 17187 20036 17196
rect 19984 17153 19993 17187
rect 19993 17153 20027 17187
rect 20027 17153 20036 17187
rect 19984 17144 20036 17153
rect 20720 17144 20772 17196
rect 15660 17076 15712 17128
rect 17316 17076 17368 17128
rect 12348 17008 12400 17060
rect 12808 17008 12860 17060
rect 13176 17008 13228 17060
rect 14372 17008 14424 17060
rect 16580 17008 16632 17060
rect 11244 16940 11296 16992
rect 13452 16940 13504 16992
rect 13544 16940 13596 16992
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 17960 16940 18012 16992
rect 19432 17076 19484 17128
rect 18696 17008 18748 17060
rect 20904 17008 20956 17060
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 22100 17076 22152 17128
rect 22192 17076 22244 17128
rect 22928 17076 22980 17128
rect 21456 17051 21508 17060
rect 21456 17017 21465 17051
rect 21465 17017 21499 17051
rect 21499 17017 21508 17051
rect 21456 17008 21508 17017
rect 24032 17008 24084 17060
rect 24124 17008 24176 17060
rect 18604 16940 18656 16992
rect 19248 16940 19300 16992
rect 20996 16983 21048 16992
rect 20996 16949 21005 16983
rect 21005 16949 21039 16983
rect 21039 16949 21048 16983
rect 20996 16940 21048 16949
rect 22100 16940 22152 16992
rect 23296 16940 23348 16992
rect 25044 16983 25096 16992
rect 25044 16949 25053 16983
rect 25053 16949 25087 16983
rect 25087 16949 25096 16983
rect 25044 16940 25096 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 10876 16779 10928 16788
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 14464 16779 14516 16788
rect 14464 16745 14473 16779
rect 14473 16745 14507 16779
rect 14507 16745 14516 16779
rect 14464 16736 14516 16745
rect 14832 16779 14884 16788
rect 14832 16745 14841 16779
rect 14841 16745 14875 16779
rect 14875 16745 14884 16779
rect 14832 16736 14884 16745
rect 16580 16736 16632 16788
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 17776 16736 17828 16788
rect 18052 16736 18104 16788
rect 18512 16779 18564 16788
rect 18512 16745 18521 16779
rect 18521 16745 18555 16779
rect 18555 16745 18564 16779
rect 19340 16779 19392 16788
rect 18512 16736 18564 16745
rect 12532 16668 12584 16720
rect 15568 16711 15620 16720
rect 15568 16677 15602 16711
rect 15602 16677 15620 16711
rect 15568 16668 15620 16677
rect 15660 16668 15712 16720
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 11612 16600 11664 16652
rect 11704 16532 11756 16584
rect 13544 16600 13596 16652
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 18972 16668 19024 16720
rect 19340 16745 19349 16779
rect 19349 16745 19383 16779
rect 19383 16745 19392 16779
rect 19340 16736 19392 16745
rect 19432 16736 19484 16788
rect 20720 16779 20772 16788
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 23940 16779 23992 16788
rect 23940 16745 23949 16779
rect 23949 16745 23983 16779
rect 23983 16745 23992 16779
rect 23940 16736 23992 16745
rect 24216 16736 24268 16788
rect 24952 16736 25004 16788
rect 21732 16668 21784 16720
rect 24124 16668 24176 16720
rect 11980 16464 12032 16516
rect 18420 16532 18472 16584
rect 19156 16600 19208 16652
rect 19984 16600 20036 16652
rect 21180 16600 21232 16652
rect 22652 16643 22704 16652
rect 22652 16609 22661 16643
rect 22661 16609 22695 16643
rect 22695 16609 22704 16643
rect 22652 16600 22704 16609
rect 18236 16464 18288 16516
rect 21272 16464 21324 16516
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 22928 16575 22980 16584
rect 21456 16532 21508 16541
rect 22928 16541 22937 16575
rect 22937 16541 22971 16575
rect 22971 16541 22980 16575
rect 22928 16532 22980 16541
rect 24216 16532 24268 16584
rect 25044 16600 25096 16652
rect 23572 16464 23624 16516
rect 12808 16396 12860 16448
rect 13820 16439 13872 16448
rect 13820 16405 13829 16439
rect 13829 16405 13863 16439
rect 13863 16405 13872 16439
rect 13820 16396 13872 16405
rect 19892 16439 19944 16448
rect 19892 16405 19901 16439
rect 19901 16405 19935 16439
rect 19935 16405 19944 16439
rect 19892 16396 19944 16405
rect 20904 16439 20956 16448
rect 20904 16405 20913 16439
rect 20913 16405 20947 16439
rect 20947 16405 20956 16439
rect 20904 16396 20956 16405
rect 22008 16439 22060 16448
rect 22008 16405 22017 16439
rect 22017 16405 22051 16439
rect 22051 16405 22060 16439
rect 22008 16396 22060 16405
rect 22192 16396 22244 16448
rect 25044 16439 25096 16448
rect 25044 16405 25053 16439
rect 25053 16405 25087 16439
rect 25087 16405 25096 16439
rect 25044 16396 25096 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 11244 16235 11296 16244
rect 11244 16201 11253 16235
rect 11253 16201 11287 16235
rect 11287 16201 11296 16235
rect 11244 16192 11296 16201
rect 11704 16235 11756 16244
rect 11704 16201 11713 16235
rect 11713 16201 11747 16235
rect 11747 16201 11756 16235
rect 11704 16192 11756 16201
rect 12440 16235 12492 16244
rect 12440 16201 12449 16235
rect 12449 16201 12483 16235
rect 12483 16201 12492 16235
rect 13544 16235 13596 16244
rect 12440 16192 12492 16201
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 15568 16192 15620 16244
rect 16212 16192 16264 16244
rect 18236 16192 18288 16244
rect 22928 16192 22980 16244
rect 23572 16192 23624 16244
rect 24216 16192 24268 16244
rect 12808 16056 12860 16108
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 13820 15988 13872 16040
rect 15292 16056 15344 16108
rect 23388 16124 23440 16176
rect 24952 16124 25004 16176
rect 16304 16056 16356 16108
rect 16488 16056 16540 16108
rect 23204 16056 23256 16108
rect 17776 15988 17828 16040
rect 20076 15988 20128 16040
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 22928 15988 22980 16040
rect 24032 16056 24084 16108
rect 24400 16056 24452 16108
rect 25596 16099 25648 16108
rect 25596 16065 25605 16099
rect 25605 16065 25639 16099
rect 25639 16065 25648 16099
rect 25596 16056 25648 16065
rect 11888 15920 11940 15972
rect 13084 15920 13136 15972
rect 18144 15920 18196 15972
rect 11612 15852 11664 15904
rect 12532 15852 12584 15904
rect 12900 15852 12952 15904
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 17500 15895 17552 15904
rect 17500 15861 17509 15895
rect 17509 15861 17543 15895
rect 17543 15861 17552 15895
rect 17500 15852 17552 15861
rect 19156 15852 19208 15904
rect 19984 15852 20036 15904
rect 20628 15920 20680 15972
rect 21272 15920 21324 15972
rect 23848 15920 23900 15972
rect 24216 15920 24268 15972
rect 21456 15852 21508 15904
rect 21548 15852 21600 15904
rect 21732 15852 21784 15904
rect 24768 15852 24820 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 13084 15648 13136 15700
rect 14188 15648 14240 15700
rect 14648 15691 14700 15700
rect 14648 15657 14657 15691
rect 14657 15657 14691 15691
rect 14691 15657 14700 15691
rect 14648 15648 14700 15657
rect 16120 15648 16172 15700
rect 17868 15648 17920 15700
rect 18144 15691 18196 15700
rect 18144 15657 18153 15691
rect 18153 15657 18187 15691
rect 18187 15657 18196 15691
rect 18144 15648 18196 15657
rect 19248 15691 19300 15700
rect 19248 15657 19257 15691
rect 19257 15657 19291 15691
rect 19291 15657 19300 15691
rect 19248 15648 19300 15657
rect 20444 15648 20496 15700
rect 20628 15648 20680 15700
rect 22008 15648 22060 15700
rect 24400 15691 24452 15700
rect 16028 15580 16080 15632
rect 16304 15580 16356 15632
rect 17132 15623 17184 15632
rect 17132 15589 17141 15623
rect 17141 15589 17175 15623
rect 17175 15589 17184 15623
rect 17132 15580 17184 15589
rect 17316 15580 17368 15632
rect 19984 15580 20036 15632
rect 11980 15512 12032 15564
rect 12164 15555 12216 15564
rect 12164 15521 12198 15555
rect 12198 15521 12216 15555
rect 12164 15512 12216 15521
rect 15292 15512 15344 15564
rect 16488 15512 16540 15564
rect 19524 15512 19576 15564
rect 10968 15308 11020 15360
rect 11152 15308 11204 15360
rect 13820 15444 13872 15496
rect 20260 15512 20312 15564
rect 20904 15512 20956 15564
rect 15568 15376 15620 15428
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 20076 15444 20128 15496
rect 24400 15657 24409 15691
rect 24409 15657 24443 15691
rect 24443 15657 24452 15691
rect 24400 15648 24452 15657
rect 24676 15648 24728 15700
rect 25044 15648 25096 15700
rect 23020 15512 23072 15564
rect 24952 15555 25004 15564
rect 24952 15521 24961 15555
rect 24961 15521 24995 15555
rect 24995 15521 25004 15555
rect 24952 15512 25004 15521
rect 26148 15512 26200 15564
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 25136 15487 25188 15496
rect 25136 15453 25145 15487
rect 25145 15453 25179 15487
rect 25179 15453 25188 15487
rect 25136 15444 25188 15453
rect 18236 15376 18288 15428
rect 23480 15376 23532 15428
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 16764 15308 16816 15360
rect 20812 15308 20864 15360
rect 23296 15308 23348 15360
rect 24768 15308 24820 15360
rect 26056 15308 26108 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 12532 15104 12584 15156
rect 15476 15104 15528 15156
rect 16488 15104 16540 15156
rect 18236 15104 18288 15156
rect 18604 15104 18656 15156
rect 20904 15104 20956 15156
rect 15568 15079 15620 15088
rect 15568 15045 15577 15079
rect 15577 15045 15611 15079
rect 15611 15045 15620 15079
rect 15568 15036 15620 15045
rect 16396 15079 16448 15088
rect 16396 15045 16405 15079
rect 16405 15045 16439 15079
rect 16439 15045 16448 15079
rect 16396 15036 16448 15045
rect 21456 15036 21508 15088
rect 11428 15011 11480 15020
rect 11428 14977 11437 15011
rect 11437 14977 11471 15011
rect 11471 14977 11480 15011
rect 11428 14968 11480 14977
rect 12164 14968 12216 15020
rect 13636 15011 13688 15020
rect 13636 14977 13645 15011
rect 13645 14977 13679 15011
rect 13679 14977 13688 15011
rect 13636 14968 13688 14977
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 16304 14968 16356 15020
rect 18604 15011 18656 15020
rect 18604 14977 18613 15011
rect 18613 14977 18647 15011
rect 18647 14977 18656 15011
rect 18604 14968 18656 14977
rect 11060 14900 11112 14952
rect 12532 14900 12584 14952
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 13728 14900 13780 14952
rect 16764 14943 16816 14952
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 17868 14900 17920 14952
rect 19984 14900 20036 14952
rect 23388 15104 23440 15156
rect 23020 15079 23072 15088
rect 23020 15045 23029 15079
rect 23029 15045 23063 15079
rect 23063 15045 23072 15079
rect 25136 15104 25188 15156
rect 26240 15147 26292 15156
rect 26240 15113 26249 15147
rect 26249 15113 26283 15147
rect 26283 15113 26292 15147
rect 26240 15104 26292 15113
rect 23020 15036 23072 15045
rect 22468 15011 22520 15020
rect 22468 14977 22477 15011
rect 22477 14977 22511 15011
rect 22511 14977 22520 15011
rect 22468 14968 22520 14977
rect 24676 14900 24728 14952
rect 12348 14832 12400 14884
rect 14280 14832 14332 14884
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 13268 14764 13320 14816
rect 17316 14764 17368 14816
rect 17500 14764 17552 14816
rect 19800 14832 19852 14884
rect 21548 14832 21600 14884
rect 24400 14875 24452 14884
rect 24400 14841 24434 14875
rect 24434 14841 24452 14875
rect 24400 14832 24452 14841
rect 25044 14832 25096 14884
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 19524 14764 19576 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 12992 14560 13044 14612
rect 15108 14603 15160 14612
rect 15108 14569 15117 14603
rect 15117 14569 15151 14603
rect 15151 14569 15160 14603
rect 15108 14560 15160 14569
rect 16304 14560 16356 14612
rect 16580 14560 16632 14612
rect 21272 14560 21324 14612
rect 21640 14560 21692 14612
rect 22560 14560 22612 14612
rect 23388 14560 23440 14612
rect 24952 14560 25004 14612
rect 11888 14492 11940 14544
rect 14004 14535 14056 14544
rect 14004 14501 14013 14535
rect 14013 14501 14047 14535
rect 14047 14501 14056 14535
rect 14004 14492 14056 14501
rect 15752 14492 15804 14544
rect 16856 14492 16908 14544
rect 10968 14467 11020 14476
rect 10968 14433 10977 14467
rect 10977 14433 11011 14467
rect 11011 14433 11020 14467
rect 10968 14424 11020 14433
rect 13176 14424 13228 14476
rect 14648 14424 14700 14476
rect 16580 14424 16632 14476
rect 19432 14424 19484 14476
rect 20812 14492 20864 14544
rect 23020 14492 23072 14544
rect 23756 14492 23808 14544
rect 19984 14424 20036 14476
rect 20996 14424 21048 14476
rect 23940 14424 23992 14476
rect 25596 14424 25648 14476
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 14188 14356 14240 14365
rect 21548 14399 21600 14408
rect 19340 14288 19392 14340
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 23296 14356 23348 14408
rect 21824 14288 21876 14340
rect 22744 14288 22796 14340
rect 24400 14288 24452 14340
rect 25228 14356 25280 14408
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 15384 14220 15436 14272
rect 15844 14220 15896 14272
rect 17960 14220 18012 14272
rect 18604 14220 18656 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 20812 14220 20864 14272
rect 22560 14220 22612 14272
rect 23572 14263 23624 14272
rect 23572 14229 23581 14263
rect 23581 14229 23615 14263
rect 23615 14229 23624 14263
rect 23572 14220 23624 14229
rect 25136 14220 25188 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 11888 14059 11940 14068
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 11888 14016 11940 14025
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 13176 14016 13228 14068
rect 14188 14016 14240 14068
rect 14648 14059 14700 14068
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 15568 14016 15620 14068
rect 19340 14016 19392 14068
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 21548 14016 21600 14068
rect 23388 14059 23440 14068
rect 23388 14025 23397 14059
rect 23397 14025 23431 14059
rect 23431 14025 23440 14059
rect 23388 14016 23440 14025
rect 23756 14016 23808 14068
rect 25044 14016 25096 14068
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 16580 13991 16632 14000
rect 16580 13957 16589 13991
rect 16589 13957 16623 13991
rect 16623 13957 16632 13991
rect 16580 13948 16632 13957
rect 20444 13948 20496 14000
rect 21824 13991 21876 14000
rect 9772 13923 9824 13932
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 10876 13880 10928 13932
rect 11888 13880 11940 13932
rect 13452 13880 13504 13932
rect 10784 13812 10836 13864
rect 15108 13880 15160 13932
rect 21824 13957 21833 13991
rect 21833 13957 21867 13991
rect 21867 13957 21876 13991
rect 21824 13948 21876 13957
rect 14372 13812 14424 13864
rect 15476 13855 15528 13864
rect 15476 13821 15510 13855
rect 15510 13821 15528 13855
rect 15476 13812 15528 13821
rect 17960 13812 18012 13864
rect 18880 13812 18932 13864
rect 22560 13923 22612 13932
rect 22560 13889 22569 13923
rect 22569 13889 22603 13923
rect 22603 13889 22612 13923
rect 22560 13880 22612 13889
rect 23296 13880 23348 13932
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 25596 13880 25648 13932
rect 23020 13855 23072 13864
rect 23020 13821 23029 13855
rect 23029 13821 23063 13855
rect 23063 13821 23072 13855
rect 23020 13812 23072 13821
rect 23940 13812 23992 13864
rect 25044 13855 25096 13864
rect 12440 13744 12492 13796
rect 13636 13744 13688 13796
rect 16764 13744 16816 13796
rect 20076 13744 20128 13796
rect 22100 13744 22152 13796
rect 22744 13744 22796 13796
rect 25044 13821 25053 13855
rect 25053 13821 25087 13855
rect 25087 13821 25096 13855
rect 25044 13812 25096 13821
rect 10692 13719 10744 13728
rect 10692 13685 10701 13719
rect 10701 13685 10735 13719
rect 10735 13685 10744 13719
rect 10692 13676 10744 13685
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 14004 13719 14056 13728
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 17592 13676 17644 13728
rect 18972 13676 19024 13728
rect 20812 13676 20864 13728
rect 22560 13676 22612 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 10048 13515 10100 13524
rect 10048 13481 10057 13515
rect 10057 13481 10091 13515
rect 10091 13481 10100 13515
rect 10048 13472 10100 13481
rect 10692 13472 10744 13524
rect 11888 13472 11940 13524
rect 11796 13404 11848 13456
rect 12348 13404 12400 13456
rect 12440 13404 12492 13456
rect 14004 13472 14056 13524
rect 16488 13472 16540 13524
rect 16764 13472 16816 13524
rect 16856 13515 16908 13524
rect 16856 13481 16865 13515
rect 16865 13481 16899 13515
rect 16899 13481 16908 13515
rect 18328 13515 18380 13524
rect 16856 13472 16908 13481
rect 18328 13481 18337 13515
rect 18337 13481 18371 13515
rect 18371 13481 18380 13515
rect 18328 13472 18380 13481
rect 18696 13472 18748 13524
rect 20996 13472 21048 13524
rect 21640 13515 21692 13524
rect 21640 13481 21649 13515
rect 21649 13481 21683 13515
rect 21683 13481 21692 13515
rect 21640 13472 21692 13481
rect 23296 13515 23348 13524
rect 23296 13481 23305 13515
rect 23305 13481 23339 13515
rect 23339 13481 23348 13515
rect 23296 13472 23348 13481
rect 13268 13404 13320 13456
rect 14556 13404 14608 13456
rect 16028 13404 16080 13456
rect 16212 13404 16264 13456
rect 17040 13447 17092 13456
rect 17040 13413 17049 13447
rect 17049 13413 17083 13447
rect 17083 13413 17092 13447
rect 17040 13404 17092 13413
rect 18972 13404 19024 13456
rect 24032 13404 24084 13456
rect 12624 13336 12676 13388
rect 14004 13379 14056 13388
rect 14004 13345 14013 13379
rect 14013 13345 14047 13379
rect 14047 13345 14056 13379
rect 14004 13336 14056 13345
rect 11060 13268 11112 13320
rect 15108 13336 15160 13388
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 16948 13336 17000 13388
rect 18880 13379 18932 13388
rect 18880 13345 18889 13379
rect 18889 13345 18923 13379
rect 18923 13345 18932 13379
rect 18880 13336 18932 13345
rect 20904 13379 20956 13388
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 22560 13336 22612 13388
rect 13636 13243 13688 13252
rect 13636 13209 13645 13243
rect 13645 13209 13679 13243
rect 13679 13209 13688 13243
rect 13636 13200 13688 13209
rect 14740 13243 14792 13252
rect 14740 13209 14749 13243
rect 14749 13209 14783 13243
rect 14783 13209 14792 13243
rect 14740 13200 14792 13209
rect 11152 13132 11204 13184
rect 12072 13132 12124 13184
rect 15384 13200 15436 13252
rect 16580 13268 16632 13320
rect 20720 13268 20772 13320
rect 21916 13268 21968 13320
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 23572 13268 23624 13320
rect 20812 13200 20864 13252
rect 22652 13200 22704 13252
rect 18328 13132 18380 13184
rect 19156 13132 19208 13184
rect 20168 13132 20220 13184
rect 22100 13175 22152 13184
rect 22100 13141 22109 13175
rect 22109 13141 22143 13175
rect 22143 13141 22152 13175
rect 22284 13175 22336 13184
rect 22100 13132 22152 13141
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 23388 13132 23440 13184
rect 25228 13175 25280 13184
rect 25228 13141 25237 13175
rect 25237 13141 25271 13175
rect 25271 13141 25280 13175
rect 25228 13132 25280 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 14004 12928 14056 12980
rect 14280 12928 14332 12980
rect 17868 12928 17920 12980
rect 18972 12928 19024 12980
rect 11888 12860 11940 12912
rect 19340 12860 19392 12912
rect 19708 12903 19760 12912
rect 19708 12869 19717 12903
rect 19717 12869 19751 12903
rect 19751 12869 19760 12903
rect 19708 12860 19760 12869
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 17500 12792 17552 12844
rect 17592 12835 17644 12844
rect 17592 12801 17601 12835
rect 17601 12801 17635 12835
rect 17635 12801 17644 12835
rect 18788 12835 18840 12844
rect 17592 12792 17644 12801
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 13084 12724 13136 12776
rect 14740 12724 14792 12776
rect 16856 12724 16908 12776
rect 18972 12792 19024 12844
rect 20536 12928 20588 12980
rect 22928 12971 22980 12980
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 24032 12928 24084 12980
rect 23664 12860 23716 12912
rect 23112 12792 23164 12844
rect 23480 12792 23532 12844
rect 11980 12656 12032 12708
rect 14832 12656 14884 12708
rect 17684 12656 17736 12708
rect 18880 12656 18932 12708
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 14740 12588 14792 12640
rect 19708 12724 19760 12776
rect 20168 12767 20220 12776
rect 20168 12733 20191 12767
rect 20191 12733 20220 12767
rect 21548 12767 21600 12776
rect 20168 12724 20220 12733
rect 21548 12733 21557 12767
rect 21557 12733 21591 12767
rect 21591 12733 21600 12767
rect 21548 12724 21600 12733
rect 22284 12724 22336 12776
rect 22928 12724 22980 12776
rect 23388 12724 23440 12776
rect 20720 12656 20772 12708
rect 21916 12699 21968 12708
rect 21916 12665 21925 12699
rect 21925 12665 21959 12699
rect 21959 12665 21968 12699
rect 21916 12656 21968 12665
rect 23756 12656 23808 12708
rect 19432 12588 19484 12640
rect 21456 12588 21508 12640
rect 22376 12588 22428 12640
rect 23572 12588 23624 12640
rect 24216 12588 24268 12640
rect 24676 12588 24728 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 10140 12384 10192 12436
rect 11060 12384 11112 12436
rect 12348 12384 12400 12436
rect 12532 12384 12584 12436
rect 13820 12384 13872 12436
rect 15108 12384 15160 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 15752 12384 15804 12436
rect 10968 12316 11020 12368
rect 12256 12248 12308 12300
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 12164 12180 12216 12232
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 15384 12316 15436 12368
rect 17040 12384 17092 12436
rect 19156 12384 19208 12436
rect 21088 12384 21140 12436
rect 22560 12427 22612 12436
rect 22560 12393 22569 12427
rect 22569 12393 22603 12427
rect 22603 12393 22612 12427
rect 22560 12384 22612 12393
rect 22928 12427 22980 12436
rect 22928 12393 22937 12427
rect 22937 12393 22971 12427
rect 22971 12393 22980 12427
rect 22928 12384 22980 12393
rect 25596 12427 25648 12436
rect 25596 12393 25605 12427
rect 25605 12393 25639 12427
rect 25639 12393 25648 12427
rect 25596 12384 25648 12393
rect 14004 12291 14056 12300
rect 14004 12257 14013 12291
rect 14013 12257 14047 12291
rect 14047 12257 14056 12291
rect 14004 12248 14056 12257
rect 14096 12291 14148 12300
rect 14096 12257 14105 12291
rect 14105 12257 14139 12291
rect 14139 12257 14148 12291
rect 14096 12248 14148 12257
rect 14280 12223 14332 12232
rect 12716 12180 12768 12189
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 11060 12112 11112 12164
rect 13452 12112 13504 12164
rect 14924 12248 14976 12300
rect 15292 12180 15344 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 17868 12316 17920 12368
rect 17960 12316 18012 12368
rect 18604 12316 18656 12368
rect 18880 12359 18932 12368
rect 18880 12325 18889 12359
rect 18889 12325 18923 12359
rect 18923 12325 18932 12359
rect 18880 12316 18932 12325
rect 22192 12316 22244 12368
rect 23296 12316 23348 12368
rect 24860 12316 24912 12368
rect 25228 12316 25280 12368
rect 16764 12248 16816 12300
rect 18788 12248 18840 12300
rect 19340 12248 19392 12300
rect 20260 12248 20312 12300
rect 21456 12248 21508 12300
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 17132 12180 17184 12232
rect 19156 12180 19208 12232
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 20536 12180 20588 12232
rect 23388 12180 23440 12232
rect 18144 12155 18196 12164
rect 12440 12044 12492 12096
rect 13084 12044 13136 12096
rect 14280 12044 14332 12096
rect 15752 12044 15804 12096
rect 16028 12044 16080 12096
rect 16580 12044 16632 12096
rect 18144 12121 18153 12155
rect 18153 12121 18187 12155
rect 18187 12121 18196 12155
rect 18144 12112 18196 12121
rect 18788 12112 18840 12164
rect 23480 12112 23532 12164
rect 24124 12112 24176 12164
rect 18236 12044 18288 12096
rect 22192 12044 22244 12096
rect 23756 12087 23808 12096
rect 23756 12053 23765 12087
rect 23765 12053 23799 12087
rect 23799 12053 23808 12087
rect 23756 12044 23808 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 10968 11840 11020 11892
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 12716 11840 12768 11892
rect 13452 11840 13504 11892
rect 14004 11840 14056 11892
rect 19892 11840 19944 11892
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 20628 11840 20680 11892
rect 21456 11883 21508 11892
rect 21456 11849 21465 11883
rect 21465 11849 21499 11883
rect 21499 11849 21508 11883
rect 21456 11840 21508 11849
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 24860 11840 24912 11892
rect 11060 11772 11112 11824
rect 12256 11704 12308 11756
rect 13360 11704 13412 11756
rect 14832 11772 14884 11824
rect 15568 11815 15620 11824
rect 15568 11781 15577 11815
rect 15577 11781 15611 11815
rect 15611 11781 15620 11815
rect 15568 11772 15620 11781
rect 12624 11636 12676 11688
rect 13084 11636 13136 11688
rect 16580 11747 16632 11756
rect 16580 11713 16589 11747
rect 16589 11713 16623 11747
rect 16623 11713 16632 11747
rect 16580 11704 16632 11713
rect 17776 11747 17828 11756
rect 17776 11713 17785 11747
rect 17785 11713 17819 11747
rect 17819 11713 17828 11747
rect 17776 11704 17828 11713
rect 21088 11747 21140 11756
rect 11152 11568 11204 11620
rect 16488 11636 16540 11688
rect 18420 11679 18472 11688
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 18328 11568 18380 11620
rect 21088 11713 21097 11747
rect 21097 11713 21131 11747
rect 21131 11713 21140 11747
rect 21088 11704 21140 11713
rect 22468 11704 22520 11756
rect 24124 11704 24176 11756
rect 24768 11747 24820 11756
rect 24768 11713 24777 11747
rect 24777 11713 24811 11747
rect 24811 11713 24820 11747
rect 24768 11704 24820 11713
rect 20352 11636 20404 11688
rect 22928 11636 22980 11688
rect 23848 11636 23900 11688
rect 20904 11611 20956 11620
rect 20904 11577 20913 11611
rect 20913 11577 20947 11611
rect 20947 11577 20956 11611
rect 20904 11568 20956 11577
rect 23388 11568 23440 11620
rect 11612 11500 11664 11552
rect 13360 11500 13412 11552
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 16304 11500 16356 11552
rect 16764 11500 16816 11552
rect 17132 11500 17184 11552
rect 17868 11500 17920 11552
rect 18788 11500 18840 11552
rect 19984 11500 20036 11552
rect 20812 11500 20864 11552
rect 22284 11500 22336 11552
rect 22928 11500 22980 11552
rect 24216 11500 24268 11552
rect 24584 11500 24636 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 12716 11296 12768 11348
rect 14096 11296 14148 11348
rect 14832 11296 14884 11348
rect 15384 11296 15436 11348
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19156 11339 19208 11348
rect 19156 11305 19165 11339
rect 19165 11305 19199 11339
rect 19199 11305 19208 11339
rect 19156 11296 19208 11305
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 20076 11296 20128 11348
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 20720 11339 20772 11348
rect 20720 11305 20729 11339
rect 20729 11305 20763 11339
rect 20763 11305 20772 11339
rect 20720 11296 20772 11305
rect 20812 11296 20864 11348
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 22284 11296 22336 11348
rect 22468 11339 22520 11348
rect 22468 11305 22477 11339
rect 22477 11305 22511 11339
rect 22511 11305 22520 11339
rect 22468 11296 22520 11305
rect 23756 11296 23808 11348
rect 24860 11339 24912 11348
rect 24860 11305 24869 11339
rect 24869 11305 24903 11339
rect 24903 11305 24912 11339
rect 24860 11296 24912 11305
rect 25872 11296 25924 11348
rect 14004 11228 14056 11280
rect 13820 11160 13872 11212
rect 14648 11160 14700 11212
rect 16580 11228 16632 11280
rect 14832 11160 14884 11212
rect 15476 11160 15528 11212
rect 19248 11160 19300 11212
rect 19984 11160 20036 11212
rect 22744 11228 22796 11280
rect 23112 11228 23164 11280
rect 23388 11228 23440 11280
rect 14004 11135 14056 11144
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 12624 11067 12676 11076
rect 12624 11033 12633 11067
rect 12633 11033 12667 11067
rect 12667 11033 12676 11067
rect 12624 11024 12676 11033
rect 13820 11024 13872 11076
rect 13268 10956 13320 11008
rect 15292 11092 15344 11144
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 19892 11135 19944 11144
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 17868 11024 17920 11076
rect 14464 10956 14516 11008
rect 15936 10956 15988 11008
rect 16948 10956 17000 11008
rect 18052 10956 18104 11008
rect 18328 10956 18380 11008
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 20720 11092 20772 11144
rect 23296 11160 23348 11212
rect 25780 11160 25832 11212
rect 20536 11024 20588 11076
rect 24584 11024 24636 11076
rect 19432 10956 19484 11008
rect 25320 10956 25372 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 15936 10752 15988 10804
rect 17592 10795 17644 10804
rect 17592 10761 17601 10795
rect 17601 10761 17635 10795
rect 17635 10761 17644 10795
rect 17592 10752 17644 10761
rect 18236 10752 18288 10804
rect 18420 10752 18472 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 20076 10752 20128 10804
rect 20720 10752 20772 10804
rect 21364 10752 21416 10804
rect 21732 10752 21784 10804
rect 25780 10795 25832 10804
rect 22744 10727 22796 10736
rect 22744 10693 22753 10727
rect 22753 10693 22787 10727
rect 22787 10693 22796 10727
rect 22744 10684 22796 10693
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 16948 10616 17000 10625
rect 19524 10616 19576 10668
rect 25780 10761 25789 10795
rect 25789 10761 25823 10795
rect 25823 10761 25832 10795
rect 25780 10752 25832 10761
rect 24308 10659 24360 10668
rect 24308 10625 24317 10659
rect 24317 10625 24351 10659
rect 24351 10625 24360 10659
rect 24308 10616 24360 10625
rect 25320 10659 25372 10668
rect 25320 10625 25329 10659
rect 25329 10625 25363 10659
rect 25363 10625 25372 10659
rect 25320 10616 25372 10625
rect 12716 10480 12768 10532
rect 13084 10548 13136 10600
rect 13268 10591 13320 10600
rect 13268 10557 13302 10591
rect 13302 10557 13320 10591
rect 13268 10548 13320 10557
rect 14188 10548 14240 10600
rect 14372 10548 14424 10600
rect 17040 10548 17092 10600
rect 17776 10548 17828 10600
rect 17960 10548 18012 10600
rect 20536 10548 20588 10600
rect 22192 10548 22244 10600
rect 24216 10548 24268 10600
rect 13728 10480 13780 10532
rect 18328 10523 18380 10532
rect 18328 10489 18362 10523
rect 18362 10489 18380 10523
rect 18328 10480 18380 10489
rect 12532 10412 12584 10464
rect 14004 10412 14056 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15016 10455 15068 10464
rect 15016 10421 15025 10455
rect 15025 10421 15059 10455
rect 15059 10421 15068 10455
rect 15016 10412 15068 10421
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 24032 10412 24084 10464
rect 24216 10455 24268 10464
rect 24216 10421 24225 10455
rect 24225 10421 24259 10455
rect 24259 10421 24268 10455
rect 24216 10412 24268 10421
rect 26148 10455 26200 10464
rect 26148 10421 26157 10455
rect 26157 10421 26191 10455
rect 26191 10421 26200 10455
rect 26148 10412 26200 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 13728 10208 13780 10260
rect 14464 10251 14516 10260
rect 14464 10217 14473 10251
rect 14473 10217 14507 10251
rect 14507 10217 14516 10251
rect 14464 10208 14516 10217
rect 16856 10208 16908 10260
rect 17040 10251 17092 10260
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 17960 10208 18012 10260
rect 19340 10251 19392 10260
rect 11244 10072 11296 10124
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 11888 10072 11940 10124
rect 11704 10004 11756 10056
rect 12900 10140 12952 10192
rect 13360 10140 13412 10192
rect 16948 10140 17000 10192
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 14464 10004 14516 10056
rect 14740 10004 14792 10056
rect 15752 10072 15804 10124
rect 16856 10072 16908 10124
rect 19340 10217 19349 10251
rect 19349 10217 19383 10251
rect 19383 10217 19392 10251
rect 19340 10208 19392 10217
rect 21824 10208 21876 10260
rect 22100 10208 22152 10260
rect 23112 10208 23164 10260
rect 19248 10183 19300 10192
rect 19248 10149 19257 10183
rect 19257 10149 19291 10183
rect 19291 10149 19300 10183
rect 19248 10140 19300 10149
rect 20352 10183 20404 10192
rect 20352 10149 20361 10183
rect 20361 10149 20395 10183
rect 20395 10149 20404 10183
rect 20352 10140 20404 10149
rect 19616 10072 19668 10124
rect 20996 10072 21048 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 22744 10072 22796 10124
rect 24308 10208 24360 10260
rect 23848 10140 23900 10192
rect 26148 10072 26200 10124
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 16672 10004 16724 10056
rect 15292 9936 15344 9988
rect 10968 9868 11020 9920
rect 15476 9868 15528 9920
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 20904 9911 20956 9920
rect 20904 9877 20913 9911
rect 20913 9877 20947 9911
rect 20947 9877 20956 9911
rect 20904 9868 20956 9877
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 10784 9639 10836 9648
rect 10784 9605 10793 9639
rect 10793 9605 10827 9639
rect 10827 9605 10836 9639
rect 10784 9596 10836 9605
rect 11704 9664 11756 9716
rect 11888 9707 11940 9716
rect 11888 9673 11897 9707
rect 11897 9673 11931 9707
rect 11931 9673 11940 9707
rect 11888 9664 11940 9673
rect 12256 9707 12308 9716
rect 12256 9673 12265 9707
rect 12265 9673 12299 9707
rect 12299 9673 12308 9707
rect 12256 9664 12308 9673
rect 12716 9664 12768 9716
rect 14372 9664 14424 9716
rect 12624 9596 12676 9648
rect 14648 9596 14700 9648
rect 15292 9664 15344 9716
rect 16212 9664 16264 9716
rect 16488 9639 16540 9648
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 14832 9528 14884 9580
rect 16488 9605 16497 9639
rect 16497 9605 16531 9639
rect 16531 9605 16540 9639
rect 16488 9596 16540 9605
rect 18236 9664 18288 9716
rect 19616 9664 19668 9716
rect 20536 9664 20588 9716
rect 21364 9664 21416 9716
rect 20720 9596 20772 9648
rect 13820 9503 13872 9512
rect 13820 9469 13829 9503
rect 13829 9469 13863 9503
rect 13863 9469 13872 9503
rect 13820 9460 13872 9469
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 15108 9460 15160 9512
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 17868 9571 17920 9580
rect 17868 9537 17877 9571
rect 17877 9537 17911 9571
rect 17911 9537 17920 9571
rect 17868 9528 17920 9537
rect 18512 9528 18564 9580
rect 19616 9571 19668 9580
rect 19616 9537 19625 9571
rect 19625 9537 19659 9571
rect 19659 9537 19668 9571
rect 19616 9528 19668 9537
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 11704 9324 11756 9376
rect 13728 9324 13780 9376
rect 14280 9324 14332 9376
rect 14740 9324 14792 9376
rect 16028 9460 16080 9512
rect 17960 9460 18012 9512
rect 16212 9392 16264 9444
rect 18328 9392 18380 9444
rect 19524 9435 19576 9444
rect 19524 9401 19533 9435
rect 19533 9401 19567 9435
rect 19567 9401 19576 9435
rect 19524 9392 19576 9401
rect 24216 9664 24268 9716
rect 21916 9528 21968 9580
rect 23848 9528 23900 9580
rect 25136 9528 25188 9580
rect 23388 9460 23440 9512
rect 15568 9324 15620 9376
rect 17960 9324 18012 9376
rect 20812 9324 20864 9376
rect 21824 9367 21876 9376
rect 21824 9333 21833 9367
rect 21833 9333 21867 9367
rect 21867 9333 21876 9367
rect 21824 9324 21876 9333
rect 23020 9367 23072 9376
rect 23020 9333 23029 9367
rect 23029 9333 23063 9367
rect 23063 9333 23072 9367
rect 23020 9324 23072 9333
rect 23480 9367 23532 9376
rect 23480 9333 23489 9367
rect 23489 9333 23523 9367
rect 23523 9333 23532 9367
rect 24216 9367 24268 9376
rect 23480 9324 23532 9333
rect 24216 9333 24225 9367
rect 24225 9333 24259 9367
rect 24259 9333 24268 9367
rect 24216 9324 24268 9333
rect 25412 9367 25464 9376
rect 25412 9333 25421 9367
rect 25421 9333 25455 9367
rect 25455 9333 25464 9367
rect 25412 9324 25464 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 12900 9120 12952 9172
rect 13820 9163 13872 9172
rect 13820 9129 13829 9163
rect 13829 9129 13863 9163
rect 13863 9129 13872 9163
rect 13820 9120 13872 9129
rect 16120 9120 16172 9172
rect 16304 9120 16356 9172
rect 17316 9120 17368 9172
rect 18052 9120 18104 9172
rect 18328 9163 18380 9172
rect 18328 9129 18337 9163
rect 18337 9129 18371 9163
rect 18371 9129 18380 9163
rect 18328 9120 18380 9129
rect 20352 9120 20404 9172
rect 21272 9120 21324 9172
rect 23112 9120 23164 9172
rect 25136 9163 25188 9172
rect 25136 9129 25145 9163
rect 25145 9129 25179 9163
rect 25179 9129 25188 9163
rect 25136 9120 25188 9129
rect 10876 9052 10928 9104
rect 10692 8984 10744 9036
rect 12256 9052 12308 9104
rect 13912 9052 13964 9104
rect 12072 9027 12124 9036
rect 12072 8993 12106 9027
rect 12106 8993 12124 9027
rect 12072 8984 12124 8993
rect 13636 8984 13688 9036
rect 13820 8984 13872 9036
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 19984 9052 20036 9104
rect 16488 8984 16540 9036
rect 10784 8916 10836 8968
rect 14832 8916 14884 8968
rect 15936 8959 15988 8968
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 16764 8916 16816 8968
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 20536 8984 20588 9036
rect 20812 8984 20864 9036
rect 21732 8984 21784 9036
rect 23388 8984 23440 9036
rect 12808 8848 12860 8900
rect 13636 8848 13688 8900
rect 15476 8848 15528 8900
rect 15660 8848 15712 8900
rect 19524 8848 19576 8900
rect 19800 8848 19852 8900
rect 11244 8823 11296 8832
rect 11244 8789 11253 8823
rect 11253 8789 11287 8823
rect 11287 8789 11296 8823
rect 11244 8780 11296 8789
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 15752 8780 15804 8832
rect 16488 8780 16540 8832
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 18604 8780 18656 8832
rect 20260 8823 20312 8832
rect 20260 8789 20269 8823
rect 20269 8789 20303 8823
rect 20303 8789 20312 8823
rect 20260 8780 20312 8789
rect 22652 8823 22704 8832
rect 22652 8789 22661 8823
rect 22661 8789 22695 8823
rect 22695 8789 22704 8823
rect 22652 8780 22704 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 12072 8576 12124 8628
rect 15660 8576 15712 8628
rect 17316 8576 17368 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 19800 8619 19852 8628
rect 19800 8585 19809 8619
rect 19809 8585 19843 8619
rect 19843 8585 19852 8619
rect 19800 8576 19852 8585
rect 20996 8576 21048 8628
rect 23940 8576 23992 8628
rect 12440 8551 12492 8560
rect 12440 8517 12449 8551
rect 12449 8517 12483 8551
rect 12483 8517 12492 8551
rect 14280 8551 14332 8560
rect 12440 8508 12492 8517
rect 14280 8517 14289 8551
rect 14289 8517 14323 8551
rect 14323 8517 14332 8551
rect 14280 8508 14332 8517
rect 21732 8508 21784 8560
rect 24124 8508 24176 8560
rect 10140 8415 10192 8424
rect 10140 8381 10149 8415
rect 10149 8381 10183 8415
rect 10183 8381 10192 8415
rect 10140 8372 10192 8381
rect 14004 8372 14056 8424
rect 14648 8372 14700 8424
rect 10968 8304 11020 8356
rect 16120 8372 16172 8424
rect 17500 8372 17552 8424
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 25044 8440 25096 8492
rect 20628 8372 20680 8424
rect 22652 8372 22704 8424
rect 23204 8372 23256 8424
rect 25412 8372 25464 8424
rect 16764 8347 16816 8356
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 16948 8347 17000 8356
rect 16948 8313 16957 8347
rect 16957 8313 16991 8347
rect 16991 8313 17000 8347
rect 16948 8304 17000 8313
rect 21916 8304 21968 8356
rect 23388 8304 23440 8356
rect 24860 8304 24912 8356
rect 10876 8236 10928 8288
rect 11336 8236 11388 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 15936 8279 15988 8288
rect 12900 8236 12952 8245
rect 15936 8245 15945 8279
rect 15945 8245 15979 8279
rect 15979 8245 15988 8279
rect 15936 8236 15988 8245
rect 20260 8279 20312 8288
rect 20260 8245 20269 8279
rect 20269 8245 20303 8279
rect 20303 8245 20312 8279
rect 20260 8236 20312 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 10692 8032 10744 8084
rect 11060 8032 11112 8084
rect 12256 8032 12308 8084
rect 12808 8075 12860 8084
rect 12808 8041 12817 8075
rect 12817 8041 12851 8075
rect 12851 8041 12860 8075
rect 12808 8032 12860 8041
rect 14004 8032 14056 8084
rect 14832 8032 14884 8084
rect 16580 8032 16632 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 24860 8032 24912 8084
rect 12900 7964 12952 8016
rect 16672 8007 16724 8016
rect 16672 7973 16681 8007
rect 16681 7973 16715 8007
rect 16715 7973 16724 8007
rect 18052 8007 18104 8016
rect 16672 7964 16724 7973
rect 18052 7973 18061 8007
rect 18061 7973 18095 8007
rect 18095 7973 18104 8007
rect 18052 7964 18104 7973
rect 18696 7964 18748 8016
rect 20444 7964 20496 8016
rect 20904 7964 20956 8016
rect 11428 7896 11480 7948
rect 13360 7939 13412 7948
rect 13360 7905 13369 7939
rect 13369 7905 13403 7939
rect 13403 7905 13412 7939
rect 13360 7896 13412 7905
rect 17592 7896 17644 7948
rect 18880 7939 18932 7948
rect 18880 7905 18889 7939
rect 18889 7905 18923 7939
rect 18923 7905 18932 7939
rect 18880 7896 18932 7905
rect 19616 7939 19668 7948
rect 19616 7905 19625 7939
rect 19625 7905 19659 7939
rect 19659 7905 19668 7939
rect 19616 7896 19668 7905
rect 21272 7939 21324 7948
rect 21272 7905 21281 7939
rect 21281 7905 21315 7939
rect 21315 7905 21324 7939
rect 21272 7896 21324 7905
rect 23756 7896 23808 7948
rect 25044 7896 25096 7948
rect 10140 7828 10192 7880
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 12164 7828 12216 7880
rect 12716 7760 12768 7812
rect 15568 7828 15620 7880
rect 14004 7760 14056 7812
rect 15936 7828 15988 7880
rect 17500 7871 17552 7880
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 17224 7760 17276 7812
rect 17500 7837 17509 7871
rect 17509 7837 17543 7871
rect 17543 7837 17552 7871
rect 17500 7828 17552 7837
rect 18788 7828 18840 7880
rect 19800 7828 19852 7880
rect 20260 7828 20312 7880
rect 21732 7828 21784 7880
rect 23296 7828 23348 7880
rect 19984 7760 20036 7812
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 23204 7692 23256 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 12256 7488 12308 7540
rect 12716 7531 12768 7540
rect 12716 7497 12725 7531
rect 12725 7497 12759 7531
rect 12759 7497 12768 7531
rect 12716 7488 12768 7497
rect 12164 7463 12216 7472
rect 12164 7429 12173 7463
rect 12173 7429 12207 7463
rect 12207 7429 12216 7463
rect 12164 7420 12216 7429
rect 11428 7395 11480 7404
rect 11428 7361 11437 7395
rect 11437 7361 11471 7395
rect 11471 7361 11480 7395
rect 11428 7352 11480 7361
rect 11888 7352 11940 7404
rect 13360 7488 13412 7540
rect 15476 7488 15528 7540
rect 13176 7284 13228 7336
rect 17500 7488 17552 7540
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 19616 7488 19668 7540
rect 20536 7531 20588 7540
rect 20536 7497 20545 7531
rect 20545 7497 20579 7531
rect 20579 7497 20588 7531
rect 20536 7488 20588 7497
rect 21272 7488 21324 7540
rect 21824 7488 21876 7540
rect 25044 7531 25096 7540
rect 25044 7497 25053 7531
rect 25053 7497 25087 7531
rect 25087 7497 25096 7531
rect 25044 7488 25096 7497
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 17592 7352 17644 7404
rect 18880 7352 18932 7404
rect 20904 7352 20956 7404
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 21732 7352 21784 7404
rect 10324 7259 10376 7268
rect 10324 7225 10333 7259
rect 10333 7225 10367 7259
rect 10367 7225 10376 7259
rect 10324 7216 10376 7225
rect 11612 7216 11664 7268
rect 13452 7216 13504 7268
rect 14648 7216 14700 7268
rect 16396 7284 16448 7336
rect 19156 7327 19208 7336
rect 19156 7293 19165 7327
rect 19165 7293 19199 7327
rect 19199 7293 19208 7327
rect 19156 7284 19208 7293
rect 18696 7216 18748 7268
rect 21824 7216 21876 7268
rect 9128 7148 9180 7200
rect 10876 7148 10928 7200
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 15752 7148 15804 7157
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 19064 7148 19116 7200
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 22744 7148 22796 7200
rect 23204 7284 23256 7336
rect 23940 7259 23992 7268
rect 23940 7225 23974 7259
rect 23974 7225 23992 7259
rect 23940 7216 23992 7225
rect 23388 7148 23440 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 11888 6944 11940 6996
rect 12900 6944 12952 6996
rect 13452 6987 13504 6996
rect 13452 6953 13461 6987
rect 13461 6953 13495 6987
rect 13495 6953 13504 6987
rect 13452 6944 13504 6953
rect 13728 6944 13780 6996
rect 14004 6987 14056 6996
rect 14004 6953 14013 6987
rect 14013 6953 14047 6987
rect 14047 6953 14056 6987
rect 14004 6944 14056 6953
rect 15568 6944 15620 6996
rect 18328 6944 18380 6996
rect 19156 6944 19208 6996
rect 19524 6944 19576 6996
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 23756 6987 23808 6996
rect 12440 6919 12492 6928
rect 12440 6885 12449 6919
rect 12449 6885 12483 6919
rect 12483 6885 12492 6919
rect 12440 6876 12492 6885
rect 15660 6876 15712 6928
rect 17868 6876 17920 6928
rect 20260 6876 20312 6928
rect 23756 6953 23765 6987
rect 23765 6953 23799 6987
rect 23799 6953 23808 6987
rect 23756 6944 23808 6953
rect 9864 6808 9916 6860
rect 10324 6808 10376 6860
rect 13176 6808 13228 6860
rect 14832 6808 14884 6860
rect 17132 6808 17184 6860
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 12532 6783 12584 6792
rect 12532 6749 12541 6783
rect 12541 6749 12575 6783
rect 12575 6749 12584 6783
rect 12532 6740 12584 6749
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 13268 6740 13320 6792
rect 14280 6783 14332 6792
rect 12348 6604 12400 6656
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 14740 6740 14792 6792
rect 15292 6740 15344 6792
rect 16672 6740 16724 6792
rect 19340 6808 19392 6860
rect 20076 6808 20128 6860
rect 21088 6808 21140 6860
rect 24216 6851 24268 6860
rect 24216 6817 24225 6851
rect 24225 6817 24259 6851
rect 24259 6817 24268 6851
rect 24216 6808 24268 6817
rect 20168 6740 20220 6792
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 23112 6740 23164 6792
rect 25412 6783 25464 6792
rect 25412 6749 25421 6783
rect 25421 6749 25455 6783
rect 25455 6749 25464 6783
rect 25412 6740 25464 6749
rect 15108 6672 15160 6724
rect 15752 6672 15804 6724
rect 16396 6672 16448 6724
rect 17684 6715 17736 6724
rect 17684 6681 17693 6715
rect 17693 6681 17727 6715
rect 17727 6681 17736 6715
rect 17684 6672 17736 6681
rect 16028 6604 16080 6656
rect 17224 6604 17276 6656
rect 18696 6604 18748 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 21272 6604 21324 6656
rect 22284 6604 22336 6656
rect 23204 6604 23256 6656
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 10324 6400 10376 6452
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 12716 6400 12768 6452
rect 13728 6400 13780 6452
rect 15568 6400 15620 6452
rect 16304 6400 16356 6452
rect 17868 6400 17920 6452
rect 18328 6443 18380 6452
rect 18328 6409 18337 6443
rect 18337 6409 18371 6443
rect 18371 6409 18380 6443
rect 18328 6400 18380 6409
rect 19616 6400 19668 6452
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23756 6400 23808 6452
rect 24216 6400 24268 6452
rect 12440 6332 12492 6384
rect 13268 6375 13320 6384
rect 13268 6341 13277 6375
rect 13277 6341 13311 6375
rect 13311 6341 13320 6375
rect 13268 6332 13320 6341
rect 12532 6264 12584 6316
rect 13452 6264 13504 6316
rect 16396 6307 16448 6316
rect 16396 6273 16405 6307
rect 16405 6273 16439 6307
rect 16439 6273 16448 6307
rect 16396 6264 16448 6273
rect 13176 6196 13228 6248
rect 13728 6239 13780 6248
rect 13728 6205 13737 6239
rect 13737 6205 13771 6239
rect 13771 6205 13780 6239
rect 13728 6196 13780 6205
rect 13820 6196 13872 6248
rect 14280 6196 14332 6248
rect 16672 6264 16724 6316
rect 18512 6264 18564 6316
rect 19984 6196 20036 6248
rect 21272 6332 21324 6384
rect 23940 6264 23992 6316
rect 25136 6307 25188 6316
rect 25136 6273 25145 6307
rect 25145 6273 25179 6307
rect 25179 6273 25188 6307
rect 25136 6264 25188 6273
rect 20996 6196 21048 6248
rect 21456 6196 21508 6248
rect 18880 6128 18932 6180
rect 21088 6128 21140 6180
rect 21640 6171 21692 6180
rect 21640 6137 21674 6171
rect 21674 6137 21692 6171
rect 21640 6128 21692 6137
rect 23756 6128 23808 6180
rect 14188 6060 14240 6112
rect 14648 6060 14700 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 20168 6060 20220 6112
rect 22928 6060 22980 6112
rect 25320 6060 25372 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 12072 5899 12124 5908
rect 12072 5865 12081 5899
rect 12081 5865 12115 5899
rect 12115 5865 12124 5899
rect 12072 5856 12124 5865
rect 13820 5899 13872 5908
rect 13820 5865 13829 5899
rect 13829 5865 13863 5899
rect 13863 5865 13872 5899
rect 13820 5856 13872 5865
rect 14280 5856 14332 5908
rect 15292 5856 15344 5908
rect 17132 5899 17184 5908
rect 17132 5865 17141 5899
rect 17141 5865 17175 5899
rect 17175 5865 17184 5899
rect 17132 5856 17184 5865
rect 18880 5899 18932 5908
rect 18880 5865 18889 5899
rect 18889 5865 18923 5899
rect 18923 5865 18932 5899
rect 18880 5856 18932 5865
rect 19340 5899 19392 5908
rect 19340 5865 19349 5899
rect 19349 5865 19383 5899
rect 19383 5865 19392 5899
rect 19340 5856 19392 5865
rect 20720 5899 20772 5908
rect 20720 5865 20729 5899
rect 20729 5865 20763 5899
rect 20763 5865 20772 5899
rect 20720 5856 20772 5865
rect 21456 5856 21508 5908
rect 23112 5856 23164 5908
rect 15568 5831 15620 5840
rect 15568 5797 15602 5831
rect 15602 5797 15620 5831
rect 15568 5788 15620 5797
rect 24124 5788 24176 5840
rect 13728 5720 13780 5772
rect 14188 5720 14240 5772
rect 17592 5720 17644 5772
rect 19708 5763 19760 5772
rect 19708 5729 19717 5763
rect 19717 5729 19751 5763
rect 19751 5729 19760 5763
rect 19708 5720 19760 5729
rect 20352 5720 20404 5772
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 23112 5720 23164 5772
rect 24860 5720 24912 5772
rect 13176 5652 13228 5704
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 17132 5652 17184 5704
rect 21364 5695 21416 5704
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 21640 5652 21692 5704
rect 23940 5584 23992 5636
rect 25136 5584 25188 5636
rect 14832 5516 14884 5568
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 20076 5516 20128 5568
rect 20168 5516 20220 5568
rect 20904 5559 20956 5568
rect 20904 5525 20913 5559
rect 20913 5525 20947 5559
rect 20947 5525 20956 5559
rect 20904 5516 20956 5525
rect 22100 5516 22152 5568
rect 22284 5516 22336 5568
rect 23204 5516 23256 5568
rect 25504 5516 25556 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 12440 5312 12492 5364
rect 13912 5312 13964 5364
rect 14280 5312 14332 5364
rect 14740 5176 14792 5228
rect 15568 5312 15620 5364
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 21640 5355 21692 5364
rect 21640 5321 21649 5355
rect 21649 5321 21683 5355
rect 21683 5321 21692 5355
rect 21640 5312 21692 5321
rect 22192 5312 22244 5364
rect 18880 5176 18932 5228
rect 19984 5219 20036 5228
rect 19984 5185 19993 5219
rect 19993 5185 20027 5219
rect 20027 5185 20036 5219
rect 19984 5176 20036 5185
rect 12624 4972 12676 5024
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 15292 5108 15344 5160
rect 17132 5108 17184 5160
rect 18788 5151 18840 5160
rect 18788 5117 18797 5151
rect 18797 5117 18831 5151
rect 18831 5117 18840 5151
rect 18788 5108 18840 5117
rect 22468 5312 22520 5364
rect 23112 5312 23164 5364
rect 23204 5176 23256 5228
rect 25136 5312 25188 5364
rect 24768 5244 24820 5296
rect 25044 5287 25096 5296
rect 25044 5253 25053 5287
rect 25053 5253 25087 5287
rect 25087 5253 25096 5287
rect 25044 5244 25096 5253
rect 25136 5176 25188 5228
rect 16672 5040 16724 5092
rect 20168 5040 20220 5092
rect 23756 5040 23808 5092
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 16120 4972 16172 5024
rect 17592 4972 17644 5024
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 18788 4972 18840 5024
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 24860 4972 24912 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 13728 4768 13780 4820
rect 14740 4811 14792 4820
rect 14740 4777 14749 4811
rect 14749 4777 14783 4811
rect 14783 4777 14792 4811
rect 14740 4768 14792 4777
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16672 4811 16724 4820
rect 16028 4768 16080 4777
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 16764 4768 16816 4820
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 21364 4768 21416 4820
rect 22560 4768 22612 4820
rect 24676 4811 24728 4820
rect 24676 4777 24685 4811
rect 24685 4777 24719 4811
rect 24719 4777 24728 4811
rect 24676 4768 24728 4777
rect 25412 4768 25464 4820
rect 14188 4743 14240 4752
rect 14188 4709 14197 4743
rect 14197 4709 14231 4743
rect 14231 4709 14240 4743
rect 14188 4700 14240 4709
rect 17040 4700 17092 4752
rect 17776 4743 17828 4752
rect 17776 4709 17785 4743
rect 17785 4709 17819 4743
rect 17819 4709 17828 4743
rect 17776 4700 17828 4709
rect 19064 4700 19116 4752
rect 12808 4675 12860 4684
rect 12808 4641 12817 4675
rect 12817 4641 12851 4675
rect 12851 4641 12860 4675
rect 12808 4632 12860 4641
rect 14556 4632 14608 4684
rect 17500 4632 17552 4684
rect 20904 4675 20956 4684
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 15292 4564 15344 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 23020 4632 23072 4684
rect 25320 4632 25372 4684
rect 18420 4564 18472 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20168 4564 20220 4616
rect 21088 4607 21140 4616
rect 21088 4573 21097 4607
rect 21097 4573 21131 4607
rect 21131 4573 21140 4607
rect 21088 4564 21140 4573
rect 22100 4564 22152 4616
rect 25044 4564 25096 4616
rect 16212 4496 16264 4548
rect 14556 4428 14608 4480
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 17592 4428 17644 4480
rect 18788 4428 18840 4480
rect 23756 4428 23808 4480
rect 24124 4471 24176 4480
rect 24124 4437 24133 4471
rect 24133 4437 24167 4471
rect 24167 4437 24176 4471
rect 24124 4428 24176 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 14556 4224 14608 4276
rect 15660 4267 15712 4276
rect 15660 4233 15669 4267
rect 15669 4233 15703 4267
rect 15703 4233 15712 4267
rect 15660 4224 15712 4233
rect 17684 4224 17736 4276
rect 17776 4267 17828 4276
rect 17776 4233 17785 4267
rect 17785 4233 17819 4267
rect 17819 4233 17828 4267
rect 17776 4224 17828 4233
rect 18880 4224 18932 4276
rect 19432 4267 19484 4276
rect 19432 4233 19441 4267
rect 19441 4233 19475 4267
rect 19475 4233 19484 4267
rect 19432 4224 19484 4233
rect 20904 4267 20956 4276
rect 20904 4233 20913 4267
rect 20913 4233 20947 4267
rect 20947 4233 20956 4267
rect 20904 4224 20956 4233
rect 12808 4156 12860 4208
rect 13544 4088 13596 4140
rect 14464 4088 14516 4140
rect 16120 4156 16172 4208
rect 17500 4156 17552 4208
rect 22836 4224 22888 4276
rect 23480 4267 23532 4276
rect 23480 4233 23489 4267
rect 23489 4233 23523 4267
rect 23523 4233 23532 4267
rect 25044 4267 25096 4276
rect 23480 4224 23532 4233
rect 15384 4088 15436 4140
rect 15476 4088 15528 4140
rect 16212 4131 16264 4140
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 19708 4131 19760 4140
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 20260 4088 20312 4140
rect 23756 4156 23808 4208
rect 23848 4088 23900 4140
rect 25044 4233 25053 4267
rect 25053 4233 25087 4267
rect 25087 4233 25096 4267
rect 25044 4224 25096 4233
rect 25412 4156 25464 4208
rect 16304 4020 16356 4072
rect 18604 4063 18656 4072
rect 18604 4029 18613 4063
rect 18613 4029 18647 4063
rect 18647 4029 18656 4063
rect 18604 4020 18656 4029
rect 18880 3995 18932 4004
rect 18880 3961 18889 3995
rect 18889 3961 18923 3995
rect 18923 3961 18932 3995
rect 18880 3952 18932 3961
rect 23572 4020 23624 4072
rect 23756 4020 23808 4072
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 21824 3995 21876 4004
rect 21824 3961 21833 3995
rect 21833 3961 21867 3995
rect 21867 3961 21876 3995
rect 21824 3952 21876 3961
rect 22560 3952 22612 4004
rect 24216 3952 24268 4004
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 13084 3927 13136 3936
rect 13084 3893 13093 3927
rect 13093 3893 13127 3927
rect 13127 3893 13136 3927
rect 13084 3884 13136 3893
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 22008 3927 22060 3936
rect 20352 3884 20404 3893
rect 22008 3893 22017 3927
rect 22017 3893 22051 3927
rect 22051 3893 22060 3927
rect 22008 3884 22060 3893
rect 23020 3927 23072 3936
rect 23020 3893 23029 3927
rect 23029 3893 23063 3927
rect 23063 3893 23072 3927
rect 23020 3884 23072 3893
rect 23480 3884 23532 3936
rect 26148 3952 26200 4004
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 13268 3680 13320 3732
rect 16028 3680 16080 3732
rect 18420 3680 18472 3732
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 20352 3680 20404 3732
rect 23848 3680 23900 3732
rect 24216 3680 24268 3732
rect 25320 3723 25372 3732
rect 25320 3689 25329 3723
rect 25329 3689 25363 3723
rect 25363 3689 25372 3723
rect 25320 3680 25372 3689
rect 12256 3612 12308 3664
rect 12624 3655 12676 3664
rect 12624 3621 12633 3655
rect 12633 3621 12667 3655
rect 12667 3621 12676 3655
rect 12624 3612 12676 3621
rect 13176 3612 13228 3664
rect 15568 3655 15620 3664
rect 15568 3621 15577 3655
rect 15577 3621 15611 3655
rect 15611 3621 15620 3655
rect 15568 3612 15620 3621
rect 16212 3612 16264 3664
rect 12348 3587 12400 3596
rect 12348 3553 12357 3587
rect 12357 3553 12391 3587
rect 12391 3553 12400 3587
rect 12348 3544 12400 3553
rect 13544 3544 13596 3596
rect 15476 3544 15528 3596
rect 17132 3612 17184 3664
rect 18144 3612 18196 3664
rect 23296 3612 23348 3664
rect 16856 3587 16908 3596
rect 16856 3553 16890 3587
rect 16890 3553 16908 3587
rect 19616 3587 19668 3596
rect 7748 3476 7800 3528
rect 8208 3476 8260 3528
rect 10876 3476 10928 3528
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 11428 3451 11480 3460
rect 11428 3417 11437 3451
rect 11437 3417 11471 3451
rect 11471 3417 11480 3451
rect 11428 3408 11480 3417
rect 12992 3408 13044 3460
rect 15476 3408 15528 3460
rect 16856 3544 16908 3553
rect 19616 3553 19625 3587
rect 19625 3553 19659 3587
rect 19659 3553 19668 3587
rect 19616 3544 19668 3553
rect 20352 3544 20404 3596
rect 22008 3587 22060 3596
rect 22008 3553 22042 3587
rect 22042 3553 22060 3587
rect 22008 3544 22060 3553
rect 23848 3544 23900 3596
rect 21732 3519 21784 3528
rect 21732 3485 21741 3519
rect 21741 3485 21775 3519
rect 21775 3485 21784 3519
rect 21732 3476 21784 3485
rect 23112 3476 23164 3528
rect 23020 3408 23072 3460
rect 24676 3476 24728 3528
rect 12624 3340 12676 3392
rect 13268 3340 13320 3392
rect 17868 3340 17920 3392
rect 19156 3383 19208 3392
rect 19156 3349 19165 3383
rect 19165 3349 19199 3383
rect 19199 3349 19208 3383
rect 19156 3340 19208 3349
rect 20260 3383 20312 3392
rect 20260 3349 20269 3383
rect 20269 3349 20303 3383
rect 20303 3349 20312 3383
rect 20260 3340 20312 3349
rect 21548 3383 21600 3392
rect 21548 3349 21557 3383
rect 21557 3349 21591 3383
rect 21591 3349 21600 3383
rect 21548 3340 21600 3349
rect 22376 3340 22428 3392
rect 24952 3340 25004 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 9956 3136 10008 3188
rect 12348 3136 12400 3188
rect 14188 3136 14240 3188
rect 16856 3179 16908 3188
rect 10968 3068 11020 3120
rect 13176 3111 13228 3120
rect 13176 3077 13185 3111
rect 13185 3077 13219 3111
rect 13219 3077 13228 3111
rect 13176 3068 13228 3077
rect 14464 3068 14516 3120
rect 12256 3000 12308 3052
rect 12348 2932 12400 2984
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17868 3179 17920 3188
rect 17868 3145 17877 3179
rect 17877 3145 17911 3179
rect 17911 3145 17920 3179
rect 17868 3136 17920 3145
rect 19156 3136 19208 3188
rect 19616 3136 19668 3188
rect 22008 3136 22060 3188
rect 22376 3136 22428 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 23480 3136 23532 3145
rect 23848 3136 23900 3188
rect 24676 3136 24728 3188
rect 21824 3068 21876 3120
rect 18144 3043 18196 3052
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 20352 3000 20404 3052
rect 19340 2932 19392 2984
rect 21732 2932 21784 2984
rect 26884 3068 26936 3120
rect 24860 2932 24912 2984
rect 17776 2864 17828 2916
rect 20260 2864 20312 2916
rect 23388 2864 23440 2916
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 14924 2796 14976 2848
rect 17408 2796 17460 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 10968 2635 11020 2644
rect 10968 2601 10977 2635
rect 10977 2601 11011 2635
rect 11011 2601 11020 2635
rect 10968 2592 11020 2601
rect 12624 2592 12676 2644
rect 13636 2592 13688 2644
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 16672 2592 16724 2644
rect 17776 2635 17828 2644
rect 17776 2601 17785 2635
rect 17785 2601 17819 2635
rect 17819 2601 17828 2635
rect 17776 2592 17828 2601
rect 20260 2635 20312 2644
rect 20260 2601 20269 2635
rect 20269 2601 20303 2635
rect 20303 2601 20312 2635
rect 20260 2592 20312 2601
rect 20444 2592 20496 2644
rect 9220 2456 9272 2508
rect 17592 2524 17644 2576
rect 13636 2456 13688 2508
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 19248 2524 19300 2576
rect 21824 2592 21876 2644
rect 22100 2592 22152 2644
rect 21916 2567 21968 2576
rect 21916 2533 21925 2567
rect 21925 2533 21959 2567
rect 21959 2533 21968 2567
rect 21916 2524 21968 2533
rect 24676 2524 24728 2576
rect 15568 2456 15620 2465
rect 19156 2499 19208 2508
rect 16764 2388 16816 2440
rect 12900 2363 12952 2372
rect 12900 2329 12909 2363
rect 12909 2329 12943 2363
rect 12943 2329 12952 2363
rect 12900 2320 12952 2329
rect 17776 2388 17828 2440
rect 19156 2465 19190 2499
rect 19190 2465 19208 2499
rect 19156 2456 19208 2465
rect 20904 2499 20956 2508
rect 20904 2465 20913 2499
rect 20913 2465 20947 2499
rect 20947 2465 20956 2499
rect 20904 2456 20956 2465
rect 24124 2456 24176 2508
rect 25136 2456 25188 2508
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 27528 2320 27580 2372
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 10508 2295 10560 2304
rect 10508 2261 10517 2295
rect 10517 2261 10551 2295
rect 10551 2261 10560 2295
rect 10508 2252 10560 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 16672 2295 16724 2304
rect 16672 2261 16681 2295
rect 16681 2261 16715 2295
rect 16715 2261 16724 2295
rect 16672 2252 16724 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 13912 552 13964 604
rect 14648 552 14700 604
<< metal2 >>
rect 294 27520 350 28000
rect 938 27520 994 28000
rect 1582 27520 1638 28000
rect 2318 27520 2374 28000
rect 2962 27520 3018 28000
rect 3698 27520 3754 28000
rect 4342 27520 4398 28000
rect 4986 27520 5042 28000
rect 5722 27520 5778 28000
rect 6366 27520 6422 28000
rect 7102 27520 7158 28000
rect 7746 27520 7802 28000
rect 8390 27520 8446 28000
rect 9126 27520 9182 28000
rect 9770 27520 9826 28000
rect 10506 27520 10562 28000
rect 11150 27520 11206 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13174 27520 13230 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15290 27520 15346 28000
rect 15934 27520 15990 28000
rect 16578 27520 16634 28000
rect 17314 27520 17370 28000
rect 17958 27520 18014 28000
rect 18694 27520 18750 28000
rect 19338 27520 19394 28000
rect 20074 27520 20130 28000
rect 20718 27520 20774 28000
rect 21362 27520 21418 28000
rect 22098 27520 22154 28000
rect 22742 27520 22798 28000
rect 23478 27520 23534 28000
rect 23754 27704 23810 27713
rect 23754 27639 23810 27648
rect 308 19378 336 27520
rect 952 24449 980 27520
rect 938 24440 994 24449
rect 938 24375 994 24384
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 296 19372 348 19378
rect 296 19314 348 19320
rect 388 19372 440 19378
rect 388 19314 440 19320
rect 400 11665 428 19314
rect 386 11656 442 11665
rect 386 11591 442 11600
rect 1412 10169 1440 22034
rect 1596 18193 1624 27520
rect 2332 22098 2360 27520
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2976 22001 3004 27520
rect 3712 23769 3740 27520
rect 3698 23760 3754 23769
rect 3698 23695 3754 23704
rect 2962 21992 3018 22001
rect 2962 21927 3018 21936
rect 4066 21040 4122 21049
rect 4066 20975 4122 20984
rect 1582 18184 1638 18193
rect 1582 18119 1638 18128
rect 4080 15473 4108 20975
rect 4356 18873 4384 27520
rect 5000 22681 5028 27520
rect 5736 25514 5764 27520
rect 5736 25486 6040 25514
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24857 6040 25486
rect 5998 24848 6054 24857
rect 5998 24783 6054 24792
rect 5998 24440 6054 24449
rect 5998 24375 6054 24384
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 4986 22672 5042 22681
rect 4986 22607 5042 22616
rect 6012 22545 6040 24375
rect 6090 23760 6146 23769
rect 6090 23695 6146 23704
rect 5998 22536 6054 22545
rect 5998 22471 6054 22480
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6104 21593 6132 23695
rect 6380 23225 6408 27520
rect 7116 23497 7144 27520
rect 7760 23905 7788 27520
rect 7746 23896 7802 23905
rect 7746 23831 7802 23840
rect 8404 23526 8432 27520
rect 9140 24177 9168 27520
rect 9126 24168 9182 24177
rect 9126 24103 9182 24112
rect 8392 23520 8444 23526
rect 7102 23488 7158 23497
rect 8392 23462 8444 23468
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 7102 23423 7158 23432
rect 6366 23216 6422 23225
rect 6366 23151 6422 23160
rect 9692 21690 9720 23462
rect 9784 21729 9812 27520
rect 10520 27418 10548 27520
rect 10520 27390 10732 27418
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10138 23488 10194 23497
rect 10138 23423 10194 23432
rect 9770 21720 9826 21729
rect 9680 21684 9732 21690
rect 9770 21655 9826 21664
rect 9680 21626 9732 21632
rect 6090 21584 6146 21593
rect 6090 21519 6146 21528
rect 10152 21350 10180 23423
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10704 23089 10732 27390
rect 11164 23497 11192 27520
rect 11610 23624 11666 23633
rect 11610 23559 11666 23568
rect 11150 23488 11206 23497
rect 11150 23423 11206 23432
rect 11150 23352 11206 23361
rect 11150 23287 11206 23296
rect 10690 23080 10746 23089
rect 10690 23015 10746 23024
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10888 22234 10916 22578
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 10244 21457 10272 21558
rect 10704 21554 10732 21830
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10230 21448 10286 21457
rect 10230 21383 10286 21392
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21078 10732 21490
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10692 21072 10744 21078
rect 10692 21014 10744 21020
rect 10796 20890 10824 21286
rect 10888 21146 10916 22170
rect 11060 21344 11112 21350
rect 10980 21304 11060 21332
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10704 20862 10824 20890
rect 10704 20806 10732 20862
rect 10692 20800 10744 20806
rect 9402 20768 9458 20777
rect 5622 20700 5918 20720
rect 10692 20742 10744 20748
rect 9402 20703 9458 20712
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 9416 20602 9444 20703
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9416 20398 9444 20538
rect 9770 20496 9826 20505
rect 9770 20431 9772 20440
rect 9824 20431 9826 20440
rect 9772 20402 9824 20408
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9770 19816 9826 19825
rect 9770 19751 9826 19760
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 4342 18864 4398 18873
rect 4342 18799 4398 18808
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 8206 16280 8262 16289
rect 8206 16215 8262 16224
rect 4066 15464 4122 15473
rect 4066 15399 4122 15408
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 1398 10160 1454 10169
rect 1398 10095 1454 10104
rect 4986 10160 5042 10169
rect 4986 10095 5042 10104
rect 294 8120 350 8129
rect 294 8055 350 8064
rect 308 480 336 8055
rect 3698 7848 3754 7857
rect 3698 7783 3754 7792
rect 2318 7304 2374 7313
rect 2318 7239 2374 7248
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 952 480 980 4111
rect 1582 2544 1638 2553
rect 1582 2479 1638 2488
rect 1596 480 1624 2479
rect 2332 480 2360 7239
rect 2962 4584 3018 4593
rect 2962 4519 3018 4528
rect 2976 480 3004 4519
rect 3712 480 3740 7783
rect 4342 3632 4398 3641
rect 4342 3567 4398 3576
rect 4356 480 4384 3567
rect 5000 480 5028 10095
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 7102 4040 7158 4049
rect 7102 3975 7158 3984
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6366 3088 6422 3097
rect 6366 3023 6422 3032
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5722 1864 5778 1873
rect 5722 1799 5778 1808
rect 5736 480 5764 1799
rect 6380 480 6408 3023
rect 7116 480 7144 3975
rect 8220 3534 8248 16215
rect 9784 13938 9812 19751
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9876 13410 9904 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10244 19310 10272 19858
rect 10232 19304 10284 19310
rect 10230 19272 10232 19281
rect 10284 19272 10286 19281
rect 10230 19207 10286 19216
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9954 16552 10010 16561
rect 9954 16487 10010 16496
rect 9968 14618 9996 16487
rect 10704 15881 10732 20742
rect 10888 19990 10916 21082
rect 10980 20602 11008 21304
rect 11060 21286 11112 21292
rect 11060 21072 11112 21078
rect 11060 21014 11112 21020
rect 11072 20602 11100 21014
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10888 19514 10916 19926
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 11164 17218 11192 23287
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11256 21690 11284 22034
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11256 21146 11284 21626
rect 11624 21434 11652 23559
rect 11624 21406 11836 21434
rect 11610 21312 11666 21321
rect 11610 21247 11666 21256
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11256 20466 11284 21082
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11256 19417 11284 20198
rect 11532 20058 11560 20538
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11242 19408 11298 19417
rect 11242 19343 11298 19352
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18426 11376 19110
rect 11520 18760 11572 18766
rect 11426 18728 11482 18737
rect 11520 18702 11572 18708
rect 11426 18663 11428 18672
rect 11480 18663 11482 18672
rect 11428 18634 11480 18640
rect 11532 18578 11560 18702
rect 11440 18550 11560 18578
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 11440 18222 11468 18550
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11428 18216 11480 18222
rect 11426 18184 11428 18193
rect 11480 18184 11482 18193
rect 11426 18119 11482 18128
rect 11164 17190 11376 17218
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 10874 16824 10930 16833
rect 10874 16759 10876 16768
rect 10928 16759 10930 16768
rect 10876 16730 10928 16736
rect 10874 16688 10930 16697
rect 11256 16658 11284 16934
rect 10874 16623 10930 16632
rect 11244 16652 11296 16658
rect 10690 15872 10746 15881
rect 10289 15804 10585 15824
rect 10690 15807 10746 15816
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10046 15328 10102 15337
rect 10046 15263 10102 15272
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10060 13530 10088 15263
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10138 14240 10194 14249
rect 10138 14175 10194 14184
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9876 13382 10088 13410
rect 9954 10024 10010 10033
rect 9954 9959 10010 9968
rect 9770 7712 9826 7721
rect 9770 7647 9826 7656
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 7760 480 7788 3470
rect 8390 3360 8446 3369
rect 8390 3295 8446 3304
rect 8404 480 8432 3295
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 1601 8800 2246
rect 8758 1592 8814 1601
rect 8758 1527 8814 1536
rect 9140 480 9168 7142
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9232 2310 9260 2450
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 1737 9260 2246
rect 9218 1728 9274 1737
rect 9218 1663 9274 1672
rect 9784 480 9812 7647
rect 9862 6896 9918 6905
rect 9862 6831 9864 6840
rect 9916 6831 9918 6840
rect 9864 6802 9916 6808
rect 9876 6458 9904 6802
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9968 3194 9996 9959
rect 10060 4049 10088 13382
rect 10152 12442 10180 14175
rect 10796 14113 10824 14758
rect 10888 14362 10916 16623
rect 11244 16594 11296 16600
rect 11256 16250 11284 16594
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10980 14940 11008 15302
rect 11060 14952 11112 14958
rect 10980 14912 11060 14940
rect 11060 14894 11112 14900
rect 11164 14498 11192 15302
rect 10980 14482 11192 14498
rect 10968 14476 11192 14482
rect 11020 14470 11192 14476
rect 10968 14418 11020 14424
rect 10888 14334 11008 14362
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10782 14104 10838 14113
rect 10782 14039 10838 14048
rect 10888 13938 10916 14214
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10784 13864 10836 13870
rect 10980 13818 11008 14334
rect 10784 13806 10836 13812
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 13670
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10796 12986 10824 13806
rect 10888 13790 11008 13818
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10782 10296 10838 10305
rect 10782 10231 10838 10240
rect 10796 9654 10824 10231
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10888 9110 10916 13790
rect 11072 13326 11100 14470
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12442 11100 13262
rect 11152 13184 11204 13190
rect 11204 13144 11284 13172
rect 11152 13126 11204 13132
rect 11256 12646 11284 13144
rect 11244 12640 11296 12646
rect 11242 12608 11244 12617
rect 11296 12608 11298 12617
rect 11242 12543 11298 12552
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10980 12209 11008 12310
rect 11152 12232 11204 12238
rect 10966 12200 11022 12209
rect 11152 12174 11204 12180
rect 10966 12135 11022 12144
rect 11060 12164 11112 12170
rect 10980 11898 11008 12135
rect 11060 12106 11112 12112
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11072 11830 11100 12106
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 11072 11665 11100 11766
rect 11058 11656 11114 11665
rect 11164 11626 11192 12174
rect 11058 11591 11114 11600
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9636 11008 9862
rect 10980 9608 11192 9636
rect 11164 9382 11192 9608
rect 11152 9376 11204 9382
rect 11150 9344 11152 9353
rect 11204 9344 11206 9353
rect 11150 9279 11206 9288
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10140 8424 10192 8430
rect 10704 8401 10732 8978
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10140 8366 10192 8372
rect 10690 8392 10746 8401
rect 10152 7886 10180 8366
rect 10690 8327 10746 8336
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8327
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10796 7886 10824 8910
rect 11256 8838 11284 10066
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10322 7304 10378 7313
rect 10322 7239 10324 7248
rect 10376 7239 10378 7248
rect 10324 7210 10376 7216
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6458 10364 6802
rect 10796 6458 10824 7822
rect 10888 7206 10916 8230
rect 10980 8106 11008 8298
rect 10980 8090 11100 8106
rect 10980 8084 11112 8090
rect 10980 8078 11060 8084
rect 11060 8026 11112 8032
rect 11256 7857 11284 8774
rect 11348 8294 11376 17190
rect 11426 15056 11482 15065
rect 11426 14991 11428 15000
rect 11480 14991 11482 15000
rect 11428 14962 11480 14968
rect 11532 14906 11560 18294
rect 11624 17202 11652 21247
rect 11702 18864 11758 18873
rect 11702 18799 11704 18808
rect 11756 18799 11758 18808
rect 11704 18770 11756 18776
rect 11716 18358 11744 18770
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17338 11744 17682
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11808 16674 11836 21406
rect 11900 20602 11928 27520
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 12070 23896 12126 23905
rect 12070 23831 12072 23840
rect 12124 23831 12126 23840
rect 12072 23802 12124 23808
rect 12084 23594 12112 23802
rect 12072 23588 12124 23594
rect 12072 23530 12124 23536
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11992 22137 12020 23054
rect 11978 22128 12034 22137
rect 11978 22063 12034 22072
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 17082 11928 17478
rect 11992 17241 12020 17614
rect 11978 17232 12034 17241
rect 11978 17167 12034 17176
rect 11980 17128 12032 17134
rect 11900 17076 11980 17082
rect 11900 17070 12032 17076
rect 11900 17054 12020 17070
rect 11624 16658 11836 16674
rect 11612 16652 11836 16658
rect 11664 16646 11836 16652
rect 11612 16594 11664 16600
rect 11624 15910 11652 16594
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16250 11744 16526
rect 11992 16522 12020 17054
rect 12176 16697 12204 24210
rect 12544 23905 12572 27520
rect 12806 24848 12862 24857
rect 12806 24783 12862 24792
rect 12820 24410 12848 24783
rect 12808 24404 12860 24410
rect 12808 24346 12860 24352
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12530 23896 12586 23905
rect 12636 23866 12664 24210
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 12530 23831 12586 23840
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 13004 23730 13032 24006
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 23497 12480 23598
rect 12532 23588 12584 23594
rect 12532 23530 12584 23536
rect 12438 23488 12494 23497
rect 12438 23423 12494 23432
rect 12452 23322 12480 23423
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12346 23216 12402 23225
rect 12346 23151 12402 23160
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12268 22234 12296 22374
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12268 21554 12296 22170
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12360 20097 12388 23151
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12452 22642 12480 23054
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 20777 12480 21286
rect 12438 20768 12494 20777
rect 12438 20703 12494 20712
rect 12346 20088 12402 20097
rect 12346 20023 12402 20032
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12268 18086 12296 18702
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12256 18080 12308 18086
rect 12254 18048 12256 18057
rect 12308 18048 12310 18057
rect 12254 17983 12310 17992
rect 12452 17762 12480 18294
rect 12360 17746 12480 17762
rect 12348 17740 12480 17746
rect 12400 17734 12480 17740
rect 12348 17682 12400 17688
rect 12544 17218 12572 23530
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12820 22098 12848 23462
rect 13004 23254 13032 23666
rect 13188 23633 13216 27520
rect 13726 24712 13782 24721
rect 13726 24647 13782 24656
rect 13740 24614 13768 24647
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13174 23624 13230 23633
rect 13174 23559 13230 23568
rect 12992 23248 13044 23254
rect 12992 23190 13044 23196
rect 13004 22438 13032 23190
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 22234 13032 22374
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 13280 22148 13308 24210
rect 13249 22120 13308 22148
rect 12808 22092 12860 22098
rect 13249 22080 13277 22120
rect 13249 22052 13308 22080
rect 12808 22034 12860 22040
rect 13280 22012 13308 22052
rect 13280 21984 13400 22012
rect 13174 21448 13230 21457
rect 13174 21383 13230 21392
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 21146 12756 21286
rect 13188 21146 13216 21383
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 13096 20262 13124 20946
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13188 20058 13216 21082
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13280 20466 13308 20878
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12820 19514 12848 19858
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12624 19236 12676 19242
rect 12624 19178 12676 19184
rect 12636 18698 12664 19178
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12728 18426 12756 18770
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12912 18290 12940 18566
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12912 17882 12940 18226
rect 13188 18222 13216 18566
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12622 17640 12678 17649
rect 12622 17575 12624 17584
rect 12676 17575 12678 17584
rect 12624 17546 12676 17552
rect 12636 17354 12664 17546
rect 12636 17326 12848 17354
rect 12544 17190 12756 17218
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12162 16688 12218 16697
rect 12162 16623 12218 16632
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11440 14878 11560 14906
rect 11336 8288 11388 8294
rect 11440 8265 11468 14878
rect 11518 13696 11574 13705
rect 11518 13631 11574 13640
rect 11532 10130 11560 13631
rect 11624 11558 11652 15846
rect 11900 14550 11928 15914
rect 11992 15570 12020 16458
rect 12360 16402 12388 17002
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12360 16374 12480 16402
rect 12452 16250 12480 16374
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12544 15910 12572 16662
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12176 15026 12204 15506
rect 12544 15162 12572 15846
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12360 14770 12388 14826
rect 12360 14742 12480 14770
rect 12254 14648 12310 14657
rect 12254 14583 12310 14592
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11900 14074 11928 14486
rect 12268 14074 12296 14583
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 13530 11928 13874
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11808 12986 11836 13398
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12918 11928 13466
rect 12360 13462 12388 14214
rect 12452 13802 12480 14742
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12072 13184 12124 13190
rect 12452 13172 12480 13398
rect 12072 13126 12124 13132
rect 12360 13144 12480 13172
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11704 10056 11756 10062
rect 11900 10033 11928 10066
rect 11704 9998 11756 10004
rect 11886 10024 11942 10033
rect 11716 9722 11744 9998
rect 11886 9959 11942 9968
rect 11900 9722 11928 9959
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11992 9466 12020 12650
rect 12084 10169 12112 13126
rect 12360 12442 12388 13144
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11898 12204 12174
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12176 11801 12204 11834
rect 12162 11792 12218 11801
rect 12268 11762 12296 12242
rect 12452 12102 12480 12718
rect 12544 12442 12572 14894
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13394 12664 13670
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12728 12322 12756 17190
rect 12820 17066 12848 17326
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 16114 12848 16390
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 13096 15978 13124 16050
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 14929 12940 15846
rect 13096 15706 13124 15914
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13188 15586 13216 17002
rect 13096 15558 13216 15586
rect 12992 14952 13044 14958
rect 12898 14920 12954 14929
rect 12992 14894 13044 14900
rect 12898 14855 12954 14864
rect 12912 12424 12940 14855
rect 13004 14618 13032 14894
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 13096 13954 13124 15558
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13188 14278 13216 14418
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 14074 13216 14214
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13096 13926 13216 13954
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12912 12396 13032 12424
rect 12728 12294 12848 12322
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12728 11898 12756 12174
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12162 11727 12218 11736
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12268 11393 12296 11698
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12254 11384 12310 11393
rect 12254 11319 12310 11328
rect 12636 11082 12664 11630
rect 12728 11354 12756 11834
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12070 10160 12126 10169
rect 12070 10095 12126 10104
rect 12254 10160 12310 10169
rect 12254 10095 12310 10104
rect 12268 9897 12296 10095
rect 12254 9888 12310 9897
rect 12254 9823 12310 9832
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 11532 9438 12020 9466
rect 11336 8230 11388 8236
rect 11426 8256 11482 8265
rect 11426 8191 11482 8200
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11242 7848 11298 7857
rect 11242 7783 11298 7792
rect 11440 7410 11468 7890
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 10876 7200 10928 7206
rect 11532 7154 11560 9438
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11610 9208 11666 9217
rect 11610 9143 11666 9152
rect 11624 7274 11652 9143
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 10876 7142 10928 7148
rect 11164 7126 11560 7154
rect 11058 7032 11114 7041
rect 11058 6967 11114 6976
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10690 4992 10746 5001
rect 10289 4924 10585 4944
rect 10690 4927 10746 4936
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10046 4040 10102 4049
rect 10046 3975 10102 3984
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10520 1465 10548 2246
rect 10506 1456 10562 1465
rect 10506 1391 10562 1400
rect 10704 1306 10732 4927
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 2689 10916 3470
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 10980 2825 11008 3062
rect 10966 2816 11022 2825
rect 10966 2751 11022 2760
rect 10874 2680 10930 2689
rect 11072 2666 11100 6967
rect 10980 2650 11100 2666
rect 10874 2615 10930 2624
rect 10968 2644 11100 2650
rect 11020 2638 11100 2644
rect 10968 2586 11020 2592
rect 10520 1278 10732 1306
rect 10520 480 10548 1278
rect 11164 480 11192 7126
rect 11716 6361 11744 9318
rect 12268 9110 12296 9658
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12346 9072 12402 9081
rect 12072 9036 12124 9042
rect 12346 9007 12402 9016
rect 12072 8978 12124 8984
rect 12084 8634 12112 8978
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11794 8256 11850 8265
rect 12360 8242 12388 9007
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12452 8401 12480 8502
rect 12438 8392 12494 8401
rect 12438 8327 12494 8336
rect 12360 8214 12480 8242
rect 11794 8191 11850 8200
rect 11808 7041 11836 8191
rect 11978 8120 12034 8129
rect 11978 8055 12034 8064
rect 12256 8084 12308 8090
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11900 7206 11928 7346
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11794 7032 11850 7041
rect 11900 7002 11928 7142
rect 11794 6967 11850 6976
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11900 6905 11928 6938
rect 11886 6896 11942 6905
rect 11886 6831 11942 6840
rect 11702 6352 11758 6361
rect 11702 6287 11758 6296
rect 11796 4616 11848 4622
rect 11794 4584 11796 4593
rect 11848 4584 11850 4593
rect 11794 4519 11850 4528
rect 11428 3936 11480 3942
rect 11888 3936 11940 3942
rect 11428 3878 11480 3884
rect 11886 3904 11888 3913
rect 11940 3904 11942 3913
rect 11440 3777 11468 3878
rect 11886 3839 11942 3848
rect 11426 3768 11482 3777
rect 11426 3703 11482 3712
rect 11992 3641 12020 8055
rect 12256 8026 12308 8032
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7478 12204 7822
rect 12268 7546 12296 8026
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12164 7472 12216 7478
rect 12452 7426 12480 8214
rect 12544 7721 12572 10406
rect 12636 9654 12664 11018
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12728 10130 12756 10474
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12728 9722 12756 10066
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12820 8906 12848 12294
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12912 9586 12940 10134
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12912 9178 12940 9522
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12808 8288 12860 8294
rect 12622 8256 12678 8265
rect 12808 8230 12860 8236
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12622 8191 12678 8200
rect 12530 7712 12586 7721
rect 12530 7647 12586 7656
rect 12164 7414 12216 7420
rect 12268 7398 12480 7426
rect 12070 6080 12126 6089
rect 12070 6015 12126 6024
rect 12084 5914 12112 6015
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 12268 3670 12296 7398
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12452 6769 12480 6870
rect 12532 6792 12584 6798
rect 12438 6760 12494 6769
rect 12532 6734 12584 6740
rect 12438 6695 12494 6704
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12256 3664 12308 3670
rect 11978 3632 12034 3641
rect 12256 3606 12308 3612
rect 11978 3567 12034 3576
rect 11426 3496 11482 3505
rect 11426 3431 11428 3440
rect 11480 3431 11482 3440
rect 11428 3402 11480 3408
rect 11886 3224 11942 3233
rect 11886 3159 11942 3168
rect 11426 2952 11482 2961
rect 11426 2887 11482 2896
rect 11440 2854 11468 2887
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 2009 11652 2246
rect 11610 2000 11666 2009
rect 11610 1935 11666 1944
rect 11900 480 11928 3159
rect 12268 3058 12296 3606
rect 12360 3602 12388 6598
rect 12452 6390 12480 6695
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12544 6322 12572 6734
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12636 6202 12664 8191
rect 12820 8090 12848 8230
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12912 8022 12940 8230
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 7546 12756 7754
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12728 6798 12756 7482
rect 12912 7002 12940 7958
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 6458 12756 6734
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12544 6174 12664 6202
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 3194 12388 3538
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12452 3074 12480 5306
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12360 3046 12480 3074
rect 12360 2990 12388 3046
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12544 480 12572 6174
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 3670 12664 4966
rect 12806 4720 12862 4729
rect 12806 4655 12808 4664
rect 12860 4655 12862 4664
rect 12808 4626 12860 4632
rect 12820 4214 12848 4626
rect 13004 4604 13032 12396
rect 13096 12102 13124 12718
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13096 11694 13124 12038
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13096 10606 13124 11630
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 13188 10452 13216 13926
rect 13280 13462 13308 14758
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13372 11762 13400 21984
rect 13464 21049 13492 24550
rect 13924 24449 13952 27520
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 14016 24614 14044 25298
rect 14568 24857 14596 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14554 24848 14610 24857
rect 14554 24783 14610 24792
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 13910 24440 13966 24449
rect 13910 24375 13966 24384
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13556 21350 13584 22034
rect 13544 21344 13596 21350
rect 13820 21344 13872 21350
rect 13544 21286 13596 21292
rect 13740 21292 13820 21298
rect 13740 21286 13872 21292
rect 13450 21040 13506 21049
rect 13450 20975 13506 20984
rect 13556 18850 13584 21286
rect 13740 21270 13860 21286
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13648 20466 13676 20810
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13648 19990 13676 20402
rect 13636 19984 13688 19990
rect 13636 19926 13688 19932
rect 13648 18970 13676 19926
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13556 18822 13676 18850
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13464 17678 13492 18226
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13450 17096 13506 17105
rect 13556 17082 13584 17682
rect 13506 17054 13584 17082
rect 13450 17031 13506 17040
rect 13464 16998 13492 17031
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13544 16992 13596 16998
rect 13648 16969 13676 18822
rect 13544 16934 13596 16940
rect 13634 16960 13690 16969
rect 13556 16658 13584 16934
rect 13634 16895 13690 16904
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13556 16250 13584 16594
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13648 16130 13676 16895
rect 13740 16289 13768 21270
rect 14016 21078 14044 24550
rect 14278 24304 14334 24313
rect 14278 24239 14334 24248
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14108 21570 14136 23258
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 14200 21690 14228 22442
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14108 21542 14228 21570
rect 14004 21072 14056 21078
rect 14004 21014 14056 21020
rect 14002 20904 14058 20913
rect 14200 20874 14228 21542
rect 14002 20839 14058 20848
rect 14188 20868 14240 20874
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13924 20398 13952 20742
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13910 20088 13966 20097
rect 13910 20023 13966 20032
rect 13818 19952 13874 19961
rect 13818 19887 13874 19896
rect 13832 19417 13860 19887
rect 13924 19786 13952 20023
rect 13912 19780 13964 19786
rect 13912 19722 13964 19728
rect 13818 19408 13874 19417
rect 13818 19343 13874 19352
rect 13818 19272 13874 19281
rect 13924 19242 13952 19722
rect 13818 19207 13874 19216
rect 13912 19236 13964 19242
rect 13832 19174 13860 19207
rect 13912 19178 13964 19184
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18290 13860 19110
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13726 16280 13782 16289
rect 13726 16215 13782 16224
rect 13464 16102 13676 16130
rect 13464 15178 13492 16102
rect 13832 16046 13860 16390
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13832 15688 13860 15982
rect 13648 15660 13860 15688
rect 13542 15600 13598 15609
rect 13542 15535 13598 15544
rect 13556 15366 13584 15535
rect 13544 15360 13596 15366
rect 13542 15328 13544 15337
rect 13596 15328 13598 15337
rect 13542 15263 13598 15272
rect 13464 15150 13584 15178
rect 13452 14272 13504 14278
rect 13450 14240 13452 14249
rect 13504 14240 13506 14249
rect 13450 14175 13506 14184
rect 13464 13938 13492 14175
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11898 13492 12106
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 10606 13308 10950
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 12912 4576 13032 4604
rect 13096 10424 13216 10452
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 2650 12664 3334
rect 12912 2972 12940 4576
rect 13096 4468 13124 10424
rect 13372 10198 13400 11494
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13450 9616 13506 9625
rect 13450 9551 13506 9560
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13372 7546 13400 7890
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13464 7426 13492 9551
rect 13372 7398 13492 7426
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13188 6866 13216 7278
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13188 6254 13216 6802
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13280 6390 13308 6734
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13004 4440 13124 4468
rect 13004 3466 13032 4440
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 13096 3369 13124 3878
rect 13188 3670 13216 5646
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4865 13308 4966
rect 13266 4856 13322 4865
rect 13266 4791 13322 4800
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3738 13308 3878
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13082 3360 13138 3369
rect 13082 3295 13138 3304
rect 13188 3126 13216 3606
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13280 2990 13308 3334
rect 13372 3097 13400 7398
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13464 7002 13492 7210
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13464 6225 13492 6258
rect 13450 6216 13506 6225
rect 13450 6151 13506 6160
rect 13556 4146 13584 15150
rect 13648 15026 13676 15660
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13832 15042 13860 15438
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13740 15014 13860 15042
rect 13740 14958 13768 15014
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13648 13258 13676 13738
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13634 11112 13690 11121
rect 13634 11047 13690 11056
rect 13648 9042 13676 11047
rect 13740 10538 13768 11494
rect 13832 11218 13860 12378
rect 13924 11778 13952 19178
rect 14016 18902 14044 20839
rect 14188 20810 14240 20816
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14094 19374 14150 19383
rect 14094 19309 14150 19318
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 14016 18426 14044 18838
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14002 14648 14058 14657
rect 14002 14583 14058 14592
rect 14016 14550 14044 14583
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 13530 14044 13670
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14016 12986 14044 13330
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14108 12594 14136 19309
rect 14200 18766 14228 19654
rect 14292 19310 14320 24239
rect 14372 23588 14424 23594
rect 14372 23530 14424 23536
rect 14384 22982 14412 23530
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22030 14412 22918
rect 14568 22778 14596 24686
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 14936 24313 14964 24618
rect 15304 24426 15332 27520
rect 15120 24410 15332 24426
rect 15948 24410 15976 27520
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16500 24886 16528 25298
rect 16028 24880 16080 24886
rect 16028 24822 16080 24828
rect 16488 24880 16540 24886
rect 16488 24822 16540 24828
rect 15108 24404 15332 24410
rect 15160 24398 15332 24404
rect 15936 24404 15988 24410
rect 15108 24346 15160 24352
rect 15936 24346 15988 24352
rect 14922 24304 14978 24313
rect 14922 24239 14978 24248
rect 15752 24268 15804 24274
rect 15752 24210 15804 24216
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14738 23896 14794 23905
rect 14738 23831 14794 23840
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14554 22536 14610 22545
rect 14554 22471 14610 22480
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 14370 21584 14426 21593
rect 14370 21519 14426 21528
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14200 18426 14228 18702
rect 14292 18465 14320 19110
rect 14278 18456 14334 18465
rect 14188 18420 14240 18426
rect 14278 18391 14334 18400
rect 14188 18362 14240 18368
rect 14200 17678 14228 18362
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14200 17338 14228 17614
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14200 15042 14228 15642
rect 14292 15144 14320 18294
rect 14384 18193 14412 21519
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14476 20058 14504 20946
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14476 18970 14504 19994
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14370 18184 14426 18193
rect 14370 18119 14426 18128
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14384 17066 14412 17682
rect 14476 17134 14504 18906
rect 14568 18426 14596 22471
rect 14660 22234 14688 22918
rect 14752 22545 14780 23831
rect 14844 23662 14872 24142
rect 15764 24070 15792 24210
rect 15934 24168 15990 24177
rect 15934 24103 15990 24112
rect 15752 24064 15804 24070
rect 15752 24006 15804 24012
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14844 23322 14872 23598
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 15580 23186 15608 23462
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15290 22672 15346 22681
rect 15580 22642 15608 23122
rect 15290 22607 15346 22616
rect 15568 22636 15620 22642
rect 14738 22536 14794 22545
rect 14738 22471 14794 22480
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15120 22234 15148 22374
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 14646 22128 14702 22137
rect 14646 22063 14648 22072
rect 14700 22063 14702 22072
rect 14830 22128 14886 22137
rect 15304 22098 15332 22607
rect 15568 22578 15620 22584
rect 14830 22063 14886 22072
rect 15292 22092 15344 22098
rect 14648 22034 14700 22040
rect 14660 21486 14688 22034
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14752 21554 14780 21966
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14752 21146 14780 21490
rect 14844 21350 14872 22063
rect 15292 22034 15344 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21690 15332 22034
rect 15580 22030 15608 22061
rect 15568 22024 15620 22030
rect 15566 21992 15568 22001
rect 15620 21992 15622 22001
rect 15566 21927 15622 21936
rect 15580 21690 15608 21927
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15474 21584 15530 21593
rect 15672 21554 15700 21830
rect 15474 21519 15530 21528
rect 15660 21548 15712 21554
rect 14832 21344 14884 21350
rect 15488 21298 15516 21519
rect 15660 21490 15712 21496
rect 14832 21286 14884 21292
rect 15396 21270 15516 21298
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 14660 19258 14688 21014
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14752 19446 14780 20198
rect 14844 19922 14872 20198
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14844 19378 14872 19858
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19514 15332 20538
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14660 19230 14872 19258
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14554 18320 14610 18329
rect 14554 18255 14610 18264
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14462 16824 14518 16833
rect 14462 16759 14464 16768
rect 14516 16759 14518 16768
rect 14464 16730 14516 16736
rect 14476 16114 14504 16730
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14292 15116 14504 15144
rect 14200 15026 14412 15042
rect 14188 15020 14412 15026
rect 14240 15014 14412 15020
rect 14188 14962 14240 14968
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14200 14074 14228 14350
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14200 13841 14228 14010
rect 14186 13832 14242 13841
rect 14186 13767 14242 13776
rect 14292 13326 14320 14826
rect 14384 13870 14412 15014
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14476 13569 14504 15116
rect 14462 13560 14518 13569
rect 14568 13546 14596 18255
rect 14660 17882 14688 19110
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14752 17814 14780 18770
rect 14740 17808 14792 17814
rect 14738 17776 14740 17785
rect 14792 17776 14794 17785
rect 14738 17711 14794 17720
rect 14648 17264 14700 17270
rect 14844 17218 14872 19230
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15014 18184 15070 18193
rect 15070 18154 15240 18170
rect 15070 18148 15252 18154
rect 15070 18142 15200 18148
rect 15014 18119 15070 18128
rect 15028 17882 15056 18119
rect 15200 18090 15252 18096
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 15120 17524 15148 18022
rect 15120 17496 15332 17524
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14648 17206 14700 17212
rect 14660 15706 14688 17206
rect 14752 17190 14872 17218
rect 14752 15745 14780 17190
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14844 16794 14872 17070
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16114 15332 17496
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 14830 16008 14886 16017
rect 14830 15943 14886 15952
rect 14738 15736 14794 15745
rect 14648 15700 14700 15706
rect 14738 15671 14794 15680
rect 14648 15642 14700 15648
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 14113 14688 14418
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14646 14104 14702 14113
rect 14646 14039 14648 14048
rect 14700 14039 14702 14048
rect 14648 14010 14700 14016
rect 14568 13518 14688 13546
rect 14462 13495 14518 13504
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12986 14320 13262
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14108 12566 14228 12594
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14016 11898 14044 12242
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13924 11750 14044 11778
rect 13910 11656 13966 11665
rect 13910 11591 13966 11600
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13726 10432 13782 10441
rect 13726 10367 13782 10376
rect 13740 10266 13768 10367
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13832 9518 13860 11018
rect 13924 9625 13952 11591
rect 14016 11286 14044 11750
rect 14108 11354 14136 12242
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14004 11280 14056 11286
rect 14200 11234 14228 12566
rect 14292 12238 14320 12922
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14004 11222 14056 11228
rect 14108 11206 14228 11234
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14016 10470 14044 11086
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13910 9616 13966 9625
rect 13910 9551 13966 9560
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3602 13584 4082
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13358 3088 13414 3097
rect 13358 3023 13414 3032
rect 13268 2984 13320 2990
rect 12912 2944 13216 2972
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12898 2408 12954 2417
rect 12898 2343 12900 2352
rect 12952 2343 12954 2352
rect 12900 2314 12952 2320
rect 13188 480 13216 2944
rect 13268 2926 13320 2932
rect 13648 2650 13676 8842
rect 13740 7857 13768 9318
rect 13832 9178 13860 9454
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13924 9110 13952 9454
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13726 7848 13782 7857
rect 13726 7783 13782 7792
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13740 6458 13768 6938
rect 13832 6497 13860 8978
rect 14002 8528 14058 8537
rect 14002 8463 14058 8472
rect 14016 8430 14044 8463
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14016 8090 14044 8366
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14016 7002 14044 7754
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14108 6746 14136 11206
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13924 6718 14136 6746
rect 13818 6488 13874 6497
rect 13728 6452 13780 6458
rect 13818 6423 13874 6432
rect 13728 6394 13780 6400
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13740 5778 13768 6190
rect 13832 5914 13860 6190
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5772 13780 5778
rect 13780 5732 13860 5760
rect 13728 5714 13780 5720
rect 13726 5672 13782 5681
rect 13726 5607 13782 5616
rect 13740 4826 13768 5607
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13832 4622 13860 5732
rect 13924 5370 13952 6718
rect 14094 6488 14150 6497
rect 14094 6423 14150 6432
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 14108 5001 14136 6423
rect 14200 6118 14228 10542
rect 14292 9602 14320 12038
rect 14476 11665 14504 13495
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14462 11656 14518 11665
rect 14462 11591 14518 11600
rect 14568 11506 14596 13398
rect 14660 13297 14688 13518
rect 14646 13288 14702 13297
rect 14752 13258 14780 14214
rect 14646 13223 14702 13232
rect 14740 13252 14792 13258
rect 14384 11478 14596 11506
rect 14384 10606 14412 11478
rect 14660 11370 14688 13223
rect 14740 13194 14792 13200
rect 14752 12782 14780 13194
rect 14844 12968 14872 15943
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 14634 15332 15506
rect 15120 14618 15332 14634
rect 15108 14612 15332 14618
rect 15160 14606 15332 14612
rect 15108 14554 15160 14560
rect 15396 14278 15424 21270
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15580 19922 15608 20810
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15672 19242 15700 19858
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15672 18970 15700 19178
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15580 18290 15608 18566
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15580 16726 15608 18226
rect 15672 17134 15700 18566
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15672 16726 15700 17070
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15580 16250 15608 16662
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15580 15434 15608 16186
rect 15658 15872 15714 15881
rect 15658 15807 15714 15816
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 15178 15608 15370
rect 15488 15162 15608 15178
rect 15476 15156 15608 15162
rect 15528 15150 15608 15156
rect 15476 15098 15528 15104
rect 15568 15088 15620 15094
rect 15566 15056 15568 15065
rect 15620 15056 15622 15065
rect 15566 14991 15622 15000
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15580 14074 15608 14991
rect 15568 14068 15620 14074
rect 15488 14028 15568 14056
rect 15106 13968 15162 13977
rect 15106 13903 15108 13912
rect 15160 13903 15162 13912
rect 15108 13874 15160 13880
rect 15488 13870 15516 14028
rect 15568 14010 15620 14016
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 13172 15148 13330
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15120 13144 15332 13172
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14844 12940 15148 12968
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14568 11342 14688 11370
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 9722 14412 10406
rect 14476 10266 14504 10950
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14292 9574 14412 9602
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 8566 14320 9318
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14292 8401 14320 8502
rect 14278 8392 14334 8401
rect 14278 8327 14334 8336
rect 14384 8129 14412 9574
rect 14370 8120 14426 8129
rect 14370 8055 14426 8064
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6254 14320 6734
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14094 4992 14150 5001
rect 14094 4927 14150 4936
rect 14200 4758 14228 5714
rect 14292 5370 14320 5850
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 14476 4146 14504 9998
rect 14568 5166 14596 11342
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14660 10810 14688 11154
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14752 10062 14780 12582
rect 14844 12322 14872 12650
rect 15120 12442 15148 12940
rect 15304 12442 15332 13144
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15396 12374 15424 13194
rect 15566 13152 15622 13161
rect 15566 13087 15622 13096
rect 15384 12368 15436 12374
rect 14844 12306 14964 12322
rect 15384 12310 15436 12316
rect 14844 12300 14976 12306
rect 14844 12294 14924 12300
rect 14844 11830 14872 12294
rect 14924 12242 14976 12248
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 12050 15332 12174
rect 15382 12064 15438 12073
rect 15304 12022 15382 12050
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11880 15332 12022
rect 15382 11999 15438 12008
rect 15028 11852 15332 11880
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14844 11354 14872 11766
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14660 8430 14688 9590
rect 14844 9586 14872 11154
rect 15028 11121 15056 11852
rect 15580 11830 15608 13087
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15292 11144 15344 11150
rect 15014 11112 15070 11121
rect 15292 11086 15344 11092
rect 15014 11047 15016 11056
rect 15068 11047 15070 11056
rect 15016 11018 15068 11024
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10792 15332 11086
rect 15028 10764 15332 10792
rect 15028 10470 15056 10764
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15028 10305 15056 10406
rect 15014 10296 15070 10305
rect 15014 10231 15070 10240
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 9930
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15396 9602 15424 11290
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15488 9926 15516 11154
rect 15672 10962 15700 15807
rect 15764 14550 15792 24006
rect 15948 23866 15976 24103
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15948 23594 15976 23802
rect 15936 23588 15988 23594
rect 15936 23530 15988 23536
rect 15934 22536 15990 22545
rect 15934 22471 15990 22480
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15856 20466 15884 21286
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15948 19825 15976 22471
rect 15934 19816 15990 19825
rect 15934 19751 15990 19760
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15856 14362 15884 18090
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15948 14521 15976 17614
rect 16040 15638 16068 24822
rect 16396 24608 16448 24614
rect 16592 24596 16620 27520
rect 16948 26852 17000 26858
rect 16948 26794 17000 26800
rect 16448 24568 16620 24596
rect 16396 24550 16448 24556
rect 16210 24440 16266 24449
rect 16210 24375 16212 24384
rect 16264 24375 16266 24384
rect 16212 24346 16264 24352
rect 16224 23662 16252 24346
rect 16672 24336 16724 24342
rect 16672 24278 16724 24284
rect 16684 23730 16712 24278
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16120 23588 16172 23594
rect 16120 23530 16172 23536
rect 16132 19553 16160 23530
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 16500 23338 16528 23462
rect 16500 23322 16620 23338
rect 16500 23316 16632 23322
rect 16500 23310 16580 23316
rect 16580 23258 16632 23264
rect 16592 22642 16620 23258
rect 16684 23050 16712 23666
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16500 22216 16528 22374
rect 16500 22188 16620 22216
rect 16592 22030 16620 22188
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16316 21350 16344 21830
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16118 19544 16174 19553
rect 16118 19479 16174 19488
rect 16316 19174 16344 21286
rect 16500 21010 16528 21966
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16500 20602 16528 20946
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 20058 16436 20198
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16500 19378 16528 20538
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16304 19168 16356 19174
rect 16488 19168 16540 19174
rect 16304 19110 16356 19116
rect 16408 19116 16488 19122
rect 16408 19110 16540 19116
rect 16224 18986 16252 19110
rect 16408 19094 16528 19110
rect 16408 18986 16436 19094
rect 16224 18958 16436 18986
rect 16592 18970 16620 20266
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16670 19408 16726 19417
rect 16670 19343 16726 19352
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16132 16697 16160 18566
rect 16224 17882 16252 18702
rect 16408 18290 16436 18770
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16118 16688 16174 16697
rect 16118 16623 16174 16632
rect 16118 16280 16174 16289
rect 16224 16250 16252 17818
rect 16118 16215 16174 16224
rect 16212 16244 16264 16250
rect 16132 16130 16160 16215
rect 16212 16186 16264 16192
rect 16132 16102 16252 16130
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16132 15706 16160 15846
rect 16224 15745 16252 16102
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16210 15736 16266 15745
rect 16120 15700 16172 15706
rect 16210 15671 16266 15680
rect 16120 15642 16172 15648
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 15934 14512 15990 14521
rect 15934 14447 15990 14456
rect 15856 14334 16160 14362
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15764 12238 15792 12378
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 12102 15792 12174
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15856 11778 15884 14214
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16040 12102 16068 13398
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15580 10934 15700 10962
rect 15764 11750 15884 11778
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 15120 9574 15424 9602
rect 15120 9518 15148 9574
rect 15108 9512 15160 9518
rect 15580 9489 15608 10934
rect 15658 10840 15714 10849
rect 15658 10775 15714 10784
rect 15108 9454 15160 9460
rect 15566 9480 15622 9489
rect 15566 9415 15622 9424
rect 14740 9376 14792 9382
rect 15568 9376 15620 9382
rect 14740 9318 14792 9324
rect 15382 9344 15438 9353
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14752 7993 14780 9318
rect 15672 9353 15700 10775
rect 15764 10130 15792 11750
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 11014 15976 11086
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10810 15976 10950
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 16040 10418 16068 12038
rect 15856 10390 16068 10418
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15568 9318 15620 9324
rect 15658 9344 15714 9353
rect 15382 9279 15438 9288
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8090 14872 8910
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14738 7984 14794 7993
rect 14738 7919 14794 7928
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7274 14688 7686
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 6798 14780 7142
rect 14844 6866 14872 8026
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 6882 15332 8774
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 15120 6854 15332 6882
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 15120 6730 15148 6854
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14568 4486 14596 4626
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 4282 14596 4422
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 3194 14228 3470
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14476 3126 14504 4082
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13648 2310 13676 2450
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13648 1873 13676 2246
rect 13634 1864 13690 1873
rect 13634 1799 13690 1808
rect 14554 1592 14610 1601
rect 14554 1527 14610 1536
rect 13912 604 13964 610
rect 13912 546 13964 552
rect 13924 480 13952 546
rect 14568 480 14596 1527
rect 14660 610 14688 6054
rect 15304 5914 15332 6734
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 4826 14780 5170
rect 14844 5001 14872 5510
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5166 15332 5646
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 14830 4992 14886 5001
rect 14830 4927 14886 4936
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 15304 4622 15332 5102
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 14738 4448 14794 4457
rect 14738 4383 14794 4392
rect 14752 3641 14780 4383
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15396 4146 15424 9279
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15488 8809 15516 8842
rect 15474 8800 15530 8809
rect 15474 8735 15530 8744
rect 15474 7984 15530 7993
rect 15474 7919 15530 7928
rect 15488 7546 15516 7919
rect 15580 7886 15608 9318
rect 15658 9279 15714 9288
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8906 15700 8978
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15672 8634 15700 8842
rect 15764 8838 15792 10066
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15580 7002 15608 7822
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15580 5846 15608 6394
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15580 5370 15608 5782
rect 15568 5364 15620 5370
rect 15488 5324 15568 5352
rect 15488 4146 15516 5324
rect 15568 5306 15620 5312
rect 15672 4282 15700 6870
rect 15764 6730 15792 7142
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15752 6112 15804 6118
rect 15750 6080 15752 6089
rect 15804 6080 15806 6089
rect 15750 6015 15806 6024
rect 15856 5930 15884 10390
rect 16132 10248 16160 14334
rect 16224 13462 16252 15671
rect 16316 15638 16344 16050
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16316 15026 16344 15574
rect 16408 15094 16436 18226
rect 16500 18086 16528 18634
rect 16592 18222 16620 18906
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16488 18080 16540 18086
rect 16540 18040 16620 18068
rect 16488 18022 16540 18028
rect 16592 17814 16620 18040
rect 16580 17808 16632 17814
rect 16580 17750 16632 17756
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16592 16794 16620 17002
rect 16580 16788 16632 16794
rect 16500 16748 16580 16776
rect 16500 16114 16528 16748
rect 16580 16730 16632 16736
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16578 15600 16634 15609
rect 16488 15564 16540 15570
rect 16578 15535 16634 15544
rect 16488 15506 16540 15512
rect 16500 15162 16528 15506
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16316 14618 16344 14962
rect 16486 14784 16542 14793
rect 16486 14719 16542 14728
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16500 13530 16528 14719
rect 16592 14618 16620 15535
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16592 14006 16620 14418
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16592 13326 16620 13942
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16592 11762 16620 12038
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16040 10220 16160 10248
rect 16040 10062 16068 10220
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16040 9518 16068 9998
rect 16224 9722 16252 9998
rect 16316 9897 16344 11494
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16302 9888 16358 9897
rect 16302 9823 16358 9832
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16040 9081 16068 9454
rect 16132 9178 16160 9522
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16026 9072 16082 9081
rect 16026 9007 16082 9016
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8294 15976 8910
rect 16132 8430 16160 9114
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15948 7886 15976 8230
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15764 5902 15884 5930
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15566 3904 15622 3913
rect 15566 3839 15622 3848
rect 15290 3768 15346 3777
rect 15290 3703 15346 3712
rect 15474 3768 15530 3777
rect 15474 3703 15530 3712
rect 14738 3632 14794 3641
rect 14738 3567 14794 3576
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2650 14964 2790
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14648 604 14700 610
rect 14648 546 14700 552
rect 15304 480 15332 3703
rect 15488 3602 15516 3703
rect 15580 3670 15608 3839
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15488 2990 15516 3402
rect 15566 3224 15622 3233
rect 15566 3159 15622 3168
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15580 2514 15608 3159
rect 15764 3097 15792 5902
rect 15842 4856 15898 4865
rect 15948 4826 15976 6054
rect 16040 4826 16068 6598
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 15842 4791 15898 4800
rect 15936 4820 15988 4826
rect 15750 3088 15806 3097
rect 15750 3023 15806 3032
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 1601 15792 2246
rect 15750 1592 15806 1601
rect 15750 1527 15806 1536
rect 15856 626 15884 4791
rect 15936 4762 15988 4768
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16040 3738 16068 4762
rect 16132 4622 16160 4966
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16132 4214 16160 4558
rect 16224 4554 16252 9386
rect 16316 9178 16344 9823
rect 16408 9761 16436 10406
rect 16394 9752 16450 9761
rect 16394 9687 16450 9696
rect 16500 9654 16528 11630
rect 16592 11286 16620 11698
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16684 10577 16712 19343
rect 16776 15450 16804 20198
rect 16868 19310 16896 22442
rect 16960 22114 16988 26794
rect 17328 25498 17356 27520
rect 17316 25492 17368 25498
rect 17316 25434 17368 25440
rect 17972 24614 18000 27520
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17408 24608 17460 24614
rect 17408 24550 17460 24556
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 17052 22234 17080 22578
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 16960 22086 17080 22114
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16960 19786 16988 20334
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16854 18184 16910 18193
rect 16854 18119 16856 18128
rect 16908 18119 16910 18128
rect 16856 18090 16908 18096
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16960 16998 16988 17750
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16794 16988 16934
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16776 15422 16988 15450
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16776 14958 16804 15302
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16868 14550 16896 14894
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16762 13968 16818 13977
rect 16762 13903 16818 13912
rect 16776 13802 16804 13903
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16776 13530 16804 13738
rect 16854 13560 16910 13569
rect 16764 13524 16816 13530
rect 16854 13495 16856 13504
rect 16764 13466 16816 13472
rect 16908 13495 16910 13504
rect 16856 13466 16908 13472
rect 16868 12782 16896 13466
rect 16960 13394 16988 15422
rect 17052 13462 17080 22086
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17236 20806 17264 21286
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17144 15638 17172 19450
rect 17236 19242 17264 20742
rect 17328 19394 17356 24550
rect 17420 19514 17448 24550
rect 18156 24410 18184 25230
rect 18708 24410 18736 27520
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19260 24614 19288 25298
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 17498 24168 17554 24177
rect 17498 24103 17554 24112
rect 17868 24132 17920 24138
rect 17512 21321 17540 24103
rect 17868 24074 17920 24080
rect 17590 23760 17646 23769
rect 17590 23695 17646 23704
rect 17498 21312 17554 21321
rect 17498 21247 17554 21256
rect 17604 20913 17632 23695
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17788 23361 17816 23462
rect 17774 23352 17830 23361
rect 17774 23287 17830 23296
rect 17880 23254 17908 24074
rect 18156 23662 18184 24346
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18616 23730 18644 24006
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18418 23624 18474 23633
rect 18418 23559 18474 23568
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17868 23248 17920 23254
rect 17868 23190 17920 23196
rect 17880 22778 17908 23190
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 18064 22234 18092 23462
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 18052 22228 18104 22234
rect 18052 22170 18104 22176
rect 18248 22030 18276 22510
rect 17776 22024 17828 22030
rect 17682 21992 17738 22001
rect 17776 21966 17828 21972
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 17682 21927 17684 21936
rect 17736 21927 17738 21936
rect 17684 21898 17736 21904
rect 17788 21146 17816 21966
rect 18248 21690 18276 21966
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17590 20904 17646 20913
rect 17590 20839 17646 20848
rect 17972 20618 18000 20946
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17880 20602 18000 20618
rect 17868 20596 18000 20602
rect 17920 20590 18000 20596
rect 17868 20538 17920 20544
rect 17880 19904 17908 20538
rect 18064 20058 18092 20742
rect 18156 20262 18184 20878
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17788 19876 17908 19904
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17328 19366 17632 19394
rect 17788 19378 17816 19876
rect 18064 19802 18092 19994
rect 17880 19774 18092 19802
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 17134 17356 19110
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 17420 16998 17448 19246
rect 17498 18320 17554 18329
rect 17498 18255 17554 18264
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17132 15632 17184 15638
rect 17132 15574 17184 15580
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17328 14822 17356 15574
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17222 14104 17278 14113
rect 17222 14039 17278 14048
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 17052 12442 17080 13398
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11558 16804 12242
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 11558 17172 12174
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 16670 10568 16726 10577
rect 16670 10503 16726 10512
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16488 9648 16540 9654
rect 16394 9616 16450 9625
rect 16488 9590 16540 9596
rect 16394 9551 16450 9560
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7410 16344 7686
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6458 16344 7346
rect 16408 7342 16436 9551
rect 16488 9036 16540 9042
rect 16540 8996 16620 9024
rect 16488 8978 16540 8984
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 7970 16528 8774
rect 16592 8090 16620 8996
rect 16684 8838 16712 9998
rect 16776 8974 16804 11494
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10674 16988 10950
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16868 10266 16896 10406
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16960 10198 16988 10610
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17052 10266 17080 10542
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 10192 17000 10198
rect 17144 10146 17172 11494
rect 16948 10134 17000 10140
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 17052 10118 17172 10146
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16684 8022 16712 8774
rect 16776 8362 16804 8910
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16672 8016 16724 8022
rect 16500 7942 16620 7970
rect 16672 7958 16724 7964
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16302 6352 16358 6361
rect 16408 6322 16436 6666
rect 16592 6497 16620 7942
rect 16776 7585 16804 8298
rect 16762 7576 16818 7585
rect 16762 7511 16818 7520
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16578 6488 16634 6497
rect 16578 6423 16634 6432
rect 16684 6322 16712 6734
rect 16302 6287 16358 6296
rect 16396 6316 16448 6322
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16224 3670 16252 4082
rect 16316 4078 16344 6287
rect 16396 6258 16448 6264
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16684 5574 16712 6258
rect 16762 6216 16818 6225
rect 16762 6151 16818 6160
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 5098 16712 5510
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16684 4826 16712 5034
rect 16776 4826 16804 6151
rect 16868 5817 16896 10066
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16960 7313 16988 8298
rect 16946 7304 17002 7313
rect 16946 7239 17002 7248
rect 16854 5808 16910 5817
rect 16854 5743 16910 5752
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17052 4758 17080 10118
rect 17236 9217 17264 14039
rect 17328 13705 17356 14758
rect 17314 13696 17370 13705
rect 17314 13631 17370 13640
rect 17222 9208 17278 9217
rect 17222 9143 17278 9152
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17328 8634 17356 9114
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17130 8392 17186 8401
rect 17130 8327 17186 8336
rect 17144 6866 17172 8327
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17236 7206 17264 7754
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 7041 17264 7142
rect 17222 7032 17278 7041
rect 17222 6967 17278 6976
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17144 5914 17172 6802
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17132 5704 17184 5710
rect 17236 5692 17264 6598
rect 17184 5664 17264 5692
rect 17132 5646 17184 5652
rect 17144 5166 17172 5646
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 17144 4486 17172 5102
rect 17314 4992 17370 5001
rect 17314 4927 17370 4936
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 17144 3670 17172 4422
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16868 3194 16896 3538
rect 16856 3188 16908 3194
rect 16776 3148 16856 3176
rect 16670 2680 16726 2689
rect 16670 2615 16672 2624
rect 16724 2615 16726 2624
rect 16672 2586 16724 2592
rect 16776 2446 16804 3148
rect 16856 3130 16908 3136
rect 16854 2816 16910 2825
rect 16854 2751 16910 2760
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16672 2304 16724 2310
rect 16670 2272 16672 2281
rect 16724 2272 16726 2281
rect 16670 2207 16726 2216
rect 16868 626 16896 2751
rect 15856 598 15976 626
rect 15948 480 15976 598
rect 16592 598 16896 626
rect 16592 480 16620 598
rect 17328 480 17356 4927
rect 17420 2854 17448 16934
rect 17512 16017 17540 18255
rect 17498 16008 17554 16017
rect 17498 15943 17554 15952
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17512 15609 17540 15846
rect 17498 15600 17554 15609
rect 17498 15535 17554 15544
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17512 12850 17540 14758
rect 17604 14113 17632 19366
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17880 18970 17908 19774
rect 18156 19378 18184 19790
rect 18248 19689 18276 21354
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18340 20058 18368 21286
rect 18432 20602 18460 23559
rect 18708 23526 18736 24210
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18604 21888 18656 21894
rect 18602 21856 18604 21865
rect 18656 21856 18658 21865
rect 18602 21791 18658 21800
rect 18616 21350 18644 21791
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18234 19680 18290 19689
rect 18234 19615 18290 19624
rect 18248 19394 18276 19615
rect 18340 19514 18368 19994
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18144 19372 18196 19378
rect 18248 19366 18460 19394
rect 18144 19314 18196 19320
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18306 18000 18566
rect 17880 18278 18000 18306
rect 17776 17740 17828 17746
rect 17880 17728 17908 18278
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17972 18057 18000 18090
rect 18052 18080 18104 18086
rect 17958 18048 18014 18057
rect 18052 18022 18104 18028
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17958 17983 18014 17992
rect 17972 17882 18000 17983
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17828 17700 17908 17728
rect 17958 17776 18014 17785
rect 17958 17711 17960 17720
rect 17776 17682 17828 17688
rect 18012 17711 18014 17720
rect 17960 17682 18012 17688
rect 17788 16794 17816 17682
rect 18064 17610 18092 18022
rect 18248 17785 18276 18022
rect 18234 17776 18290 17785
rect 18234 17711 18290 17720
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17202 18276 17478
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17696 14793 17724 16594
rect 17788 16046 17816 16730
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 15745 17816 15982
rect 17774 15736 17830 15745
rect 17774 15671 17830 15680
rect 17868 15700 17920 15706
rect 17972 15688 18000 16934
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17920 15660 18000 15688
rect 17868 15642 17920 15648
rect 18064 15042 18092 16730
rect 18248 16522 18276 17138
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18248 16250 18276 16458
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18156 15706 18184 15914
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18248 15434 18276 16186
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 17880 15014 18092 15042
rect 17880 14958 17908 15014
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 18052 14816 18104 14822
rect 17682 14784 17738 14793
rect 18052 14758 18104 14764
rect 17682 14719 17738 14728
rect 18064 14657 18092 14758
rect 18050 14648 18106 14657
rect 18050 14583 18106 14592
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17590 14104 17646 14113
rect 17590 14039 17646 14048
rect 17972 13870 18000 14214
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17866 13696 17922 13705
rect 17604 12889 17632 13670
rect 17866 13631 17922 13640
rect 17682 13016 17738 13025
rect 17880 12986 17908 13631
rect 17682 12951 17738 12960
rect 17868 12980 17920 12986
rect 17590 12880 17646 12889
rect 17500 12844 17552 12850
rect 17590 12815 17592 12824
rect 17500 12786 17552 12792
rect 17644 12815 17646 12824
rect 17592 12786 17644 12792
rect 17604 12755 17632 12786
rect 17696 12714 17724 12951
rect 17868 12922 17920 12928
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 18248 12617 18276 15098
rect 18340 13530 18368 17682
rect 18432 16590 18460 19366
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18524 18154 18552 18770
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18524 17814 18552 18090
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18616 17082 18644 21286
rect 18524 17054 18644 17082
rect 18708 17066 18736 23462
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22506 18920 22918
rect 18880 22500 18932 22506
rect 18880 22442 18932 22448
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18892 21554 18920 21830
rect 19260 21729 19288 24550
rect 19352 23866 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19444 24070 19472 24686
rect 19996 24614 20024 25298
rect 20088 24682 20116 27520
rect 20168 24744 20220 24750
rect 20168 24686 20220 24692
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19246 21720 19302 21729
rect 19246 21655 19302 21664
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18892 20942 18920 21490
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18892 20262 18920 20878
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18800 18465 18828 20198
rect 18892 20058 18920 20198
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18892 19446 18920 19994
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 19076 19174 19104 20266
rect 19168 19854 19196 20334
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19168 19378 19196 19790
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 18786 18456 18842 18465
rect 18786 18391 18842 18400
rect 18696 17060 18748 17066
rect 18524 16794 18552 17054
rect 18696 17002 18748 17008
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18524 15609 18552 16730
rect 18510 15600 18566 15609
rect 18510 15535 18566 15544
rect 18616 15162 18644 16934
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18512 14816 18564 14822
rect 18510 14784 18512 14793
rect 18564 14784 18566 14793
rect 18510 14719 18566 14728
rect 18616 14278 18644 14962
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18708 14090 18736 17002
rect 18616 14062 18736 14090
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18234 12608 18290 12617
rect 18234 12543 18290 12552
rect 17868 12368 17920 12374
rect 17960 12368 18012 12374
rect 17920 12328 17960 12356
rect 17868 12310 17920 12316
rect 17960 12310 18012 12316
rect 18142 12200 18198 12209
rect 18142 12135 18144 12144
rect 18196 12135 18198 12144
rect 18144 12106 18196 12112
rect 18236 12096 18288 12102
rect 18156 12044 18236 12050
rect 18156 12038 18288 12044
rect 18156 12022 18276 12038
rect 18050 11928 18106 11937
rect 18050 11863 18106 11872
rect 17774 11792 17830 11801
rect 17774 11727 17776 11736
rect 17828 11727 17830 11736
rect 17776 11698 17828 11704
rect 17868 11552 17920 11558
rect 17788 11512 17868 11540
rect 17590 11384 17646 11393
rect 17590 11319 17646 11328
rect 17604 10810 17632 11319
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17788 10606 17816 11512
rect 17868 11494 17920 11500
rect 18064 11393 18092 11863
rect 18050 11384 18106 11393
rect 18050 11319 18052 11328
rect 18104 11319 18106 11328
rect 18052 11290 18104 11296
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17880 9704 17908 11018
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17972 10441 18000 10542
rect 17958 10432 18014 10441
rect 17958 10367 18014 10376
rect 17972 10266 18000 10367
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17880 9676 18000 9704
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17500 8968 17552 8974
rect 17498 8936 17500 8945
rect 17552 8936 17554 8945
rect 17498 8871 17554 8880
rect 17512 8430 17540 8871
rect 17880 8634 17908 9522
rect 17972 9518 18000 9676
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17512 7886 17540 8366
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17512 7546 17540 7822
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17604 7449 17632 7890
rect 17590 7440 17646 7449
rect 17590 7375 17592 7384
rect 17644 7375 17646 7384
rect 17592 7346 17644 7352
rect 17604 7315 17632 7346
rect 17868 6928 17920 6934
rect 17498 6896 17554 6905
rect 17868 6870 17920 6876
rect 17498 6831 17500 6840
rect 17552 6831 17554 6840
rect 17500 6802 17552 6808
rect 17512 4690 17540 6802
rect 17682 6760 17738 6769
rect 17682 6695 17684 6704
rect 17736 6695 17738 6704
rect 17684 6666 17736 6672
rect 17880 6458 17908 6870
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17604 5030 17632 5714
rect 17682 5128 17738 5137
rect 17682 5063 17738 5072
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17696 4826 17724 5063
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17512 4214 17540 4626
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17420 1873 17448 2790
rect 17604 2582 17632 4422
rect 17696 4282 17724 4762
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17788 4282 17816 4694
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17972 3777 18000 9318
rect 18064 9178 18092 10950
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18064 8022 18092 8366
rect 18156 8265 18184 12022
rect 18340 11914 18368 13126
rect 18616 12374 18644 14062
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18248 11886 18368 11914
rect 18248 10810 18276 11886
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18340 11014 18368 11562
rect 18432 11121 18460 11630
rect 18418 11112 18474 11121
rect 18418 11047 18474 11056
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18340 10538 18368 10950
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18340 10033 18368 10474
rect 18326 10024 18382 10033
rect 18248 9982 18326 10010
rect 18248 9722 18276 9982
rect 18326 9959 18382 9968
rect 18326 9752 18382 9761
rect 18236 9716 18288 9722
rect 18326 9687 18382 9696
rect 18236 9658 18288 9664
rect 18340 9450 18368 9687
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18340 9178 18368 9386
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18142 8256 18198 8265
rect 18142 8191 18198 8200
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18340 6458 18368 6938
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18432 6202 18460 10746
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18524 9586 18552 9862
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18524 6322 18552 7686
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18432 6174 18552 6202
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18432 4622 18460 4966
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 17958 3768 18014 3777
rect 18432 3738 18460 4558
rect 17958 3703 18014 3712
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18050 3496 18106 3505
rect 18050 3431 18106 3440
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17880 3194 17908 3334
rect 17868 3188 17920 3194
rect 17788 3148 17868 3176
rect 17788 2922 17816 3148
rect 17868 3130 17920 3136
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17788 2650 17816 2858
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17788 2446 17816 2586
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17406 1864 17462 1873
rect 17406 1799 17462 1808
rect 18064 1442 18092 3431
rect 18156 3097 18184 3606
rect 18524 3505 18552 6174
rect 18616 4078 18644 8774
rect 18708 8401 18736 13466
rect 18800 12850 18828 18391
rect 18892 14929 18920 19110
rect 19076 18426 19104 19110
rect 19168 18902 19196 19314
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19260 18306 19288 21655
rect 19352 21146 19380 21898
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19444 21010 19472 23598
rect 19996 23594 20024 24550
rect 19984 23588 20036 23594
rect 19984 23530 20036 23536
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19536 23186 19564 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19982 23216 20038 23225
rect 19524 23180 19576 23186
rect 19982 23151 20038 23160
rect 19524 23122 19576 23128
rect 19536 22574 19564 23122
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19536 21962 19564 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19628 21690 19656 22034
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19522 21584 19578 21593
rect 19522 21519 19524 21528
rect 19576 21519 19578 21528
rect 19524 21490 19576 21496
rect 19628 21457 19656 21626
rect 19720 21554 19748 21966
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19614 21448 19670 21457
rect 19614 21383 19670 21392
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19522 21040 19578 21049
rect 19432 21004 19484 21010
rect 19522 20975 19578 20984
rect 19706 21040 19762 21049
rect 19706 20975 19708 20984
rect 19432 20946 19484 20952
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19242 19380 19654
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19352 18970 19380 19178
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19076 18278 19288 18306
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 18972 17536 19024 17542
rect 18970 17504 18972 17513
rect 19024 17504 19026 17513
rect 18970 17439 19026 17448
rect 18984 16726 19012 17439
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18878 14920 18934 14929
rect 18878 14855 18934 14864
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18970 13832 19026 13841
rect 18892 13394 18920 13806
rect 18970 13767 19026 13776
rect 18984 13734 19012 13767
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 13462 19012 13670
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18892 12866 18920 13330
rect 18984 12986 19012 13398
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18892 12850 19012 12866
rect 18788 12844 18840 12850
rect 18892 12844 19024 12850
rect 18892 12838 18972 12844
rect 18788 12786 18840 12792
rect 18972 12786 19024 12792
rect 18800 12306 18828 12786
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 18892 12374 18920 12650
rect 18970 12608 19026 12617
rect 18970 12543 19026 12552
rect 18880 12368 18932 12374
rect 18878 12336 18880 12345
rect 18932 12336 18934 12345
rect 18788 12300 18840 12306
rect 18878 12271 18934 12280
rect 18788 12242 18840 12248
rect 18892 12245 18920 12271
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18800 11558 18828 12106
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18694 8392 18750 8401
rect 18694 8327 18750 8336
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18708 7546 18736 7958
rect 18800 7886 18828 11494
rect 18878 7984 18934 7993
rect 18878 7919 18880 7928
rect 18932 7919 18934 7928
rect 18880 7890 18932 7896
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18708 6662 18736 7210
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 5137 18736 6598
rect 18892 6186 18920 7346
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18892 5914 18920 6122
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18786 5400 18842 5409
rect 18786 5335 18842 5344
rect 18800 5166 18828 5335
rect 18892 5234 18920 5850
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18788 5160 18840 5166
rect 18694 5128 18750 5137
rect 18788 5102 18840 5108
rect 18694 5063 18750 5072
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18800 4486 18828 4966
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18892 4282 18920 5170
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18616 3738 18644 4014
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18510 3496 18566 3505
rect 18510 3431 18566 3440
rect 18142 3088 18198 3097
rect 18142 3023 18144 3032
rect 18196 3023 18198 3032
rect 18144 2994 18196 3000
rect 18892 1737 18920 3946
rect 18878 1728 18934 1737
rect 18878 1663 18934 1672
rect 17972 1414 18092 1442
rect 18694 1456 18750 1465
rect 17972 480 18000 1414
rect 18694 1391 18750 1400
rect 18708 480 18736 1391
rect 18984 921 19012 12543
rect 19076 12073 19104 18278
rect 19340 18080 19392 18086
rect 19260 18040 19340 18068
rect 19260 17610 19288 18040
rect 19340 18022 19392 18028
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19248 16992 19300 16998
rect 19246 16960 19248 16969
rect 19300 16960 19302 16969
rect 19246 16895 19302 16904
rect 19352 16794 19380 17750
rect 19444 17134 19472 18294
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19444 16794 19472 17070
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19168 15910 19196 16594
rect 19246 16416 19302 16425
rect 19246 16351 19302 16360
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19168 13190 19196 15846
rect 19260 15706 19288 16351
rect 19248 15700 19300 15706
rect 19536 15688 19564 20975
rect 19760 20975 19762 20984
rect 19708 20946 19760 20952
rect 19996 20369 20024 23151
rect 20074 22400 20130 22409
rect 20074 22335 20130 22344
rect 20088 21146 20116 22335
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 19982 20360 20038 20369
rect 19982 20295 20038 20304
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 20074 20088 20130 20097
rect 20074 20023 20076 20032
rect 20128 20023 20130 20032
rect 20076 19994 20128 20000
rect 20180 19961 20208 24686
rect 20732 24410 20760 27520
rect 21376 24954 21404 27520
rect 21548 26648 21600 26654
rect 21548 26590 21600 26596
rect 21364 24948 21416 24954
rect 21364 24890 21416 24896
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20456 22438 20484 22918
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20364 21350 20392 21830
rect 20444 21616 20496 21622
rect 20442 21584 20444 21593
rect 20496 21584 20498 21593
rect 20442 21519 20498 21528
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20364 21146 20392 21286
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20350 21040 20406 21049
rect 20350 20975 20406 20984
rect 20364 20058 20392 20975
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20166 19952 20222 19961
rect 19708 19916 19760 19922
rect 20166 19887 20222 19896
rect 19708 19858 19760 19864
rect 19720 19310 19748 19858
rect 20180 19666 20208 19887
rect 20180 19638 20392 19666
rect 20166 19544 20222 19553
rect 20166 19479 20222 19488
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19996 18426 20024 18906
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17678 20024 18362
rect 20088 18358 20116 18566
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 20088 18222 20116 18294
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20180 17814 20208 19479
rect 20258 18728 20314 18737
rect 20258 18663 20314 18672
rect 20272 18290 20300 18663
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19996 17338 20024 17614
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19982 17232 20038 17241
rect 19982 17167 19984 17176
rect 20036 17167 20038 17176
rect 19984 17138 20036 17144
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19904 16153 19932 16390
rect 19890 16144 19946 16153
rect 19890 16079 19946 16088
rect 19996 15910 20024 16594
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19536 15660 19656 15688
rect 19248 15642 19300 15648
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19536 14822 19564 15506
rect 19628 15065 19656 15660
rect 19996 15638 20024 15846
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 20088 15502 20116 15982
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 19614 15056 19670 15065
rect 19614 14991 19670 15000
rect 19812 14890 19840 15438
rect 20088 15042 20116 15438
rect 19996 15014 20116 15042
rect 19996 14958 20024 15014
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19154 12608 19210 12617
rect 19154 12543 19210 12552
rect 19168 12442 19196 12543
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19156 12232 19208 12238
rect 19260 12220 19288 14214
rect 19352 14074 19380 14282
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19352 13546 19380 14010
rect 19444 13705 19472 14418
rect 19430 13696 19486 13705
rect 19430 13631 19486 13640
rect 19352 13518 19472 13546
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19352 12306 19380 12854
rect 19444 12646 19472 13518
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19208 12192 19288 12220
rect 19156 12174 19208 12180
rect 19062 12064 19118 12073
rect 19062 11999 19118 12008
rect 19168 11354 19196 12174
rect 19246 11656 19302 11665
rect 19246 11591 19302 11600
rect 19260 11354 19288 11591
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19260 11098 19288 11154
rect 19260 11070 19380 11098
rect 19246 10704 19302 10713
rect 19246 10639 19302 10648
rect 19260 10198 19288 10639
rect 19352 10266 19380 11070
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19444 10810 19472 10950
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19536 10674 19564 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19708 12912 19760 12918
rect 19706 12880 19708 12889
rect 19760 12880 19762 12889
rect 19706 12815 19762 12824
rect 19720 12782 19748 12815
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19892 12232 19944 12238
rect 19890 12200 19892 12209
rect 19944 12200 19946 12209
rect 19890 12135 19946 12144
rect 19904 11898 19932 12135
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19996 11558 20024 14418
rect 20074 14104 20130 14113
rect 20272 14074 20300 15506
rect 20074 14039 20076 14048
rect 20128 14039 20130 14048
rect 20260 14068 20312 14074
rect 20076 14010 20128 14016
rect 20260 14010 20312 14016
rect 20088 13802 20116 14010
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20180 12782 20208 13126
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20180 12617 20208 12718
rect 20166 12608 20222 12617
rect 20166 12543 20222 12552
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 20074 11520 20130 11529
rect 19622 11452 19918 11472
rect 20074 11455 20130 11464
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20088 11354 20116 11455
rect 20272 11354 20300 12242
rect 20364 11898 20392 19638
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20456 14006 20484 15642
rect 20548 15178 20576 24006
rect 20640 23338 20668 24142
rect 20916 23769 20944 24210
rect 21560 23866 21588 26590
rect 22008 24608 22060 24614
rect 22112 24596 22140 27520
rect 22756 25498 22784 27520
rect 23386 26616 23442 26625
rect 23386 26551 23442 26560
rect 23294 26072 23350 26081
rect 23294 26007 23350 26016
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22560 25356 22612 25362
rect 22560 25298 22612 25304
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22060 24568 22140 24596
rect 22008 24550 22060 24556
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 20902 23760 20958 23769
rect 20902 23695 20904 23704
rect 20956 23695 20958 23704
rect 20904 23666 20956 23672
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20640 23322 20760 23338
rect 20640 23316 20772 23322
rect 20640 23310 20720 23316
rect 20720 23258 20772 23264
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20640 21622 20668 23054
rect 20732 22234 20760 23258
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20824 21865 20852 23598
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20994 22944 21050 22953
rect 20916 22098 20944 22918
rect 20994 22879 21050 22888
rect 21008 22137 21036 22879
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 20994 22128 21050 22137
rect 20904 22092 20956 22098
rect 20994 22063 21050 22072
rect 20904 22034 20956 22040
rect 20810 21856 20866 21865
rect 20810 21791 20866 21800
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20916 21486 20944 22034
rect 20994 21720 21050 21729
rect 20994 21655 21050 21664
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 21008 21418 21036 21655
rect 20996 21412 21048 21418
rect 20996 21354 21048 21360
rect 21100 21026 21128 22714
rect 21284 22574 21312 23122
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21376 22778 21404 23054
rect 22204 22953 22232 24686
rect 22572 24614 22600 25298
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 22376 24268 22428 24274
rect 22376 24210 22428 24216
rect 22388 23118 22416 24210
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22652 23520 22704 23526
rect 22652 23462 22704 23468
rect 22480 23361 22508 23462
rect 22466 23352 22522 23361
rect 22466 23287 22522 23296
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 22190 22944 22246 22953
rect 22190 22879 22246 22888
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21454 22672 21510 22681
rect 21454 22607 21510 22616
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21180 22092 21232 22098
rect 21180 22034 21232 22040
rect 21192 21554 21220 22034
rect 21284 21894 21312 22510
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21362 21856 21418 21865
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21192 21146 21220 21490
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21100 20998 21220 21026
rect 21284 21010 21312 21830
rect 21362 21791 21418 21800
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 21086 20360 21142 20369
rect 20732 20058 20760 20334
rect 21086 20295 21142 20304
rect 21100 20262 21128 20295
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20732 19496 20760 19994
rect 20732 19468 20852 19496
rect 20718 19408 20774 19417
rect 20718 19343 20774 19352
rect 20732 18970 20760 19343
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20732 18222 20760 18906
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20824 17513 20852 19468
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20810 17504 20866 17513
rect 20810 17439 20866 17448
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20732 16794 20760 17138
rect 20916 17066 20944 17614
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20628 15972 20680 15978
rect 20732 15960 20760 16730
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20680 15932 20760 15960
rect 20628 15914 20680 15920
rect 20640 15706 20668 15914
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20916 15570 20944 16390
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20548 15150 20760 15178
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20442 13560 20498 13569
rect 20442 13495 20498 13504
rect 20456 13025 20484 13495
rect 20732 13326 20760 15150
rect 20824 14550 20852 15302
rect 20916 15162 20944 15506
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 21008 14482 21036 16934
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20824 13734 20852 14214
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20824 13258 20852 13670
rect 21008 13530 21036 14418
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21100 13410 21128 20198
rect 21192 18834 21220 20998
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21284 20602 21312 20946
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21284 20330 21312 20538
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21376 20058 21404 21791
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21284 19174 21312 19858
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 19009 21312 19110
rect 21270 19000 21326 19009
rect 21468 18970 21496 22607
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22572 22166 22600 22374
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21914 21448 21970 21457
rect 22020 21434 22048 21558
rect 22572 21554 22600 21830
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22020 21406 22140 21434
rect 21914 21383 21970 21392
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21744 20466 21772 20946
rect 21928 20534 21956 21383
rect 22112 21350 22140 21406
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22020 21185 22048 21286
rect 22006 21176 22062 21185
rect 22006 21111 22062 21120
rect 22376 20800 22428 20806
rect 22296 20748 22376 20754
rect 22296 20742 22428 20748
rect 22296 20726 22416 20742
rect 22006 20632 22062 20641
rect 22006 20567 22008 20576
rect 22060 20567 22062 20576
rect 22008 20538 22060 20544
rect 21916 20528 21968 20534
rect 21916 20470 21968 20476
rect 21732 20460 21784 20466
rect 21732 20402 21784 20408
rect 21546 20360 21602 20369
rect 21546 20295 21602 20304
rect 21270 18935 21326 18944
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21192 18329 21220 18770
rect 21178 18320 21234 18329
rect 21178 18255 21234 18264
rect 21270 17776 21326 17785
rect 21270 17711 21272 17720
rect 21324 17711 21326 17720
rect 21272 17682 21324 17688
rect 21284 17338 21312 17682
rect 21560 17678 21588 20295
rect 21822 18320 21878 18329
rect 21822 18255 21824 18264
rect 21876 18255 21878 18264
rect 21824 18226 21876 18232
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21928 17270 21956 20470
rect 22296 20330 22324 20726
rect 22572 20466 22600 21490
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22112 19718 22140 20198
rect 22296 19854 22324 20266
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22100 19712 22152 19718
rect 22098 19680 22100 19689
rect 22152 19680 22154 19689
rect 22098 19615 22154 19624
rect 22006 19272 22062 19281
rect 22006 19207 22062 19216
rect 22100 19236 22152 19242
rect 22020 19174 22048 19207
rect 22100 19178 22152 19184
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22112 17882 22140 19178
rect 22296 18766 22324 19790
rect 22388 19514 22416 19858
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22664 19378 22692 23462
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 22848 22574 22876 23122
rect 22836 22568 22888 22574
rect 22834 22536 22836 22545
rect 22888 22536 22890 22545
rect 22834 22471 22890 22480
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22756 20806 22784 21830
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22572 18970 22600 19314
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22756 19174 22784 19246
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 22100 17128 22152 17134
rect 21454 17096 21510 17105
rect 22100 17070 22152 17076
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 21454 17031 21456 17040
rect 21508 17031 21510 17040
rect 21456 17002 21508 17008
rect 22112 16998 22140 17070
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21192 16425 21220 16594
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21178 16416 21234 16425
rect 21178 16351 21234 16360
rect 21192 16017 21220 16351
rect 21178 16008 21234 16017
rect 21284 15978 21312 16458
rect 21178 15943 21234 15952
rect 21272 15972 21324 15978
rect 21272 15914 21324 15920
rect 21284 14618 21312 15914
rect 21468 15910 21496 16526
rect 21744 15910 21772 16662
rect 22204 16454 22232 17070
rect 22296 16794 22324 18702
rect 22388 18426 22416 18770
rect 22650 18728 22706 18737
rect 22650 18663 22706 18672
rect 22664 18426 22692 18663
rect 22756 18426 22784 19110
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22480 17542 22508 18158
rect 22558 17912 22614 17921
rect 22558 17847 22614 17856
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 17377 22508 17478
rect 22466 17368 22522 17377
rect 22466 17303 22522 17312
rect 22572 17202 22600 17847
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22374 17096 22430 17105
rect 22374 17031 22430 17040
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21468 15094 21496 15846
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21560 14890 21588 15846
rect 22020 15706 22048 16390
rect 22284 16040 22336 16046
rect 22282 16008 22284 16017
rect 22336 16008 22338 16017
rect 22282 15943 22338 15952
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21730 15464 21786 15473
rect 21730 15399 21786 15408
rect 21548 14884 21600 14890
rect 21548 14826 21600 14832
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21560 14414 21588 14826
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 14074 21588 14350
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21178 13968 21234 13977
rect 21178 13903 21234 13912
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 21008 13382 21128 13410
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20442 13016 20498 13025
rect 20442 12951 20498 12960
rect 20536 12980 20588 12986
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20364 11694 20392 11834
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 10713 19932 11086
rect 19890 10704 19946 10713
rect 19524 10668 19576 10674
rect 19890 10639 19946 10648
rect 19524 10610 19576 10616
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19340 10260 19392 10266
rect 19996 10248 20024 11154
rect 20088 10810 20116 11290
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 19340 10202 19392 10208
rect 19904 10220 20024 10248
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19628 9722 19656 10066
rect 19904 9926 19932 10220
rect 20352 10192 20404 10198
rect 20350 10160 20352 10169
rect 20404 10160 20406 10169
rect 20350 10095 20406 10104
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19628 9586 19656 9658
rect 19904 9625 19932 9862
rect 19890 9616 19946 9625
rect 19616 9580 19668 9586
rect 19890 9551 19946 9560
rect 19616 9522 19668 9528
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19430 8936 19486 8945
rect 19536 8906 19564 9386
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19430 8871 19486 8880
rect 19524 8900 19576 8906
rect 19444 8634 19472 8871
rect 19524 8842 19576 8848
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19812 8634 19840 8842
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19154 7984 19210 7993
rect 19154 7919 19210 7928
rect 19616 7948 19668 7954
rect 19168 7342 19196 7919
rect 19616 7890 19668 7896
rect 19628 7857 19656 7890
rect 19800 7880 19852 7886
rect 19614 7848 19670 7857
rect 19614 7783 19670 7792
rect 19798 7848 19800 7857
rect 19852 7848 19854 7857
rect 19996 7818 20024 9046
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20272 8294 20300 8774
rect 20260 8288 20312 8294
rect 20074 8256 20130 8265
rect 20260 8230 20312 8236
rect 20074 8191 20130 8200
rect 19798 7783 19854 7792
rect 19984 7812 20036 7818
rect 19628 7546 19656 7783
rect 19984 7754 20036 7760
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19522 7304 19578 7313
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19076 4758 19104 7142
rect 19168 7002 19196 7278
rect 19522 7239 19578 7248
rect 19536 7002 19564 7239
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 6225 19288 6598
rect 19246 6216 19302 6225
rect 19246 6151 19302 6160
rect 19352 5914 19380 6802
rect 19536 6474 19564 6938
rect 20088 6866 20116 8191
rect 20272 7886 20300 8230
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20272 7206 20300 7822
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 6934 20300 7142
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20074 6488 20130 6497
rect 19536 6458 19656 6474
rect 19536 6452 19668 6458
rect 19536 6446 19616 6452
rect 20074 6423 20130 6432
rect 19616 6394 19668 6400
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19522 5672 19578 5681
rect 19522 5607 19578 5616
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19444 4282 19472 4558
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19168 3194 19196 3334
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19168 2514 19196 3130
rect 19340 2984 19392 2990
rect 19260 2932 19340 2938
rect 19260 2926 19392 2932
rect 19260 2910 19380 2926
rect 19260 2582 19288 2910
rect 19338 2816 19394 2825
rect 19338 2751 19394 2760
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 18970 912 19026 921
rect 18970 847 19026 856
rect 19352 480 19380 2751
rect 19536 1442 19564 5607
rect 19720 5370 19748 5714
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19996 5234 20024 6190
rect 20088 5817 20116 6423
rect 20180 6118 20208 6734
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20074 5808 20130 5817
rect 20074 5743 20130 5752
rect 20180 5574 20208 6054
rect 20364 5778 20392 9114
rect 20456 8022 20484 12951
rect 20536 12922 20588 12928
rect 20548 12238 20576 12922
rect 20916 12753 20944 13330
rect 20902 12744 20958 12753
rect 20720 12708 20772 12714
rect 20640 12668 20720 12696
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20548 11082 20576 12174
rect 20640 11898 20668 12668
rect 20902 12679 20958 12688
rect 20720 12650 20772 12656
rect 20718 12608 20774 12617
rect 20718 12543 20774 12552
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20732 11354 20760 12543
rect 20902 11656 20958 11665
rect 20902 11591 20904 11600
rect 20956 11591 20958 11600
rect 20904 11562 20956 11568
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20824 11354 20852 11494
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20548 10606 20576 11018
rect 20732 10810 20760 11086
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20548 9926 20576 10542
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9722 20576 9862
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20548 9194 20576 9658
rect 20732 9654 20760 10746
rect 21008 10248 21036 13382
rect 21086 12472 21142 12481
rect 21086 12407 21088 12416
rect 21140 12407 21142 12416
rect 21088 12378 21140 12384
rect 21100 11762 21128 12378
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21008 10220 21128 10248
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 20810 10024 20866 10033
rect 20810 9959 20866 9968
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20824 9382 20852 9959
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20548 9166 20852 9194
rect 20824 9042 20852 9166
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20444 8016 20496 8022
rect 20444 7958 20496 7964
rect 20548 7546 20576 8978
rect 20628 8424 20680 8430
rect 20626 8392 20628 8401
rect 20680 8392 20682 8401
rect 20626 8327 20682 8336
rect 20916 8022 20944 9862
rect 21008 8634 21036 10066
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20904 8016 20956 8022
rect 20904 7958 20956 7964
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20916 7410 20944 7958
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 21008 6254 21036 8570
rect 21100 8129 21128 10220
rect 21192 9761 21220 13903
rect 21652 13530 21680 14554
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21548 12776 21600 12782
rect 21546 12744 21548 12753
rect 21600 12744 21602 12753
rect 21546 12679 21602 12688
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21468 12306 21496 12582
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21468 11898 21496 12242
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21362 11792 21418 11801
rect 21362 11727 21418 11736
rect 21376 11354 21404 11727
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21376 10810 21404 11290
rect 21744 10810 21772 15399
rect 21822 14920 21878 14929
rect 21822 14855 21878 14864
rect 21836 14346 21864 14855
rect 22190 14512 22246 14521
rect 22190 14447 22246 14456
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21836 14006 21864 14282
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 22006 13832 22062 13841
rect 22006 13767 22062 13776
rect 22100 13796 22152 13802
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21928 12714 21956 13262
rect 21916 12708 21968 12714
rect 21916 12650 21968 12656
rect 22020 11898 22048 13767
rect 22100 13738 22152 13744
rect 22112 13190 22140 13738
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 21822 10976 21878 10985
rect 21822 10911 21878 10920
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21270 10568 21326 10577
rect 21270 10503 21326 10512
rect 21284 10130 21312 10503
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21178 9752 21234 9761
rect 21178 9687 21234 9696
rect 21284 9178 21312 10066
rect 21376 9722 21404 10746
rect 21836 10266 21864 10911
rect 22112 10266 22140 13126
rect 22204 12374 22232 14447
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22296 12782 22324 13126
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22388 12646 22416 17031
rect 22558 16960 22614 16969
rect 22558 16895 22614 16904
rect 22466 15056 22522 15065
rect 22466 14991 22468 15000
rect 22520 14991 22522 15000
rect 22468 14962 22520 14968
rect 22572 14618 22600 16895
rect 22650 16688 22706 16697
rect 22650 16623 22652 16632
rect 22704 16623 22706 16632
rect 22652 16594 22704 16600
rect 22756 16538 22784 18158
rect 22664 16510 22784 16538
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22572 13938 22600 14214
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22572 13818 22600 13874
rect 22480 13790 22600 13818
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22480 12481 22508 13790
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22572 13394 22600 13670
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22466 12472 22522 12481
rect 22572 12442 22600 13330
rect 22664 13258 22692 16510
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22756 13802 22784 14282
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22466 12407 22522 12416
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22192 12368 22244 12374
rect 22192 12310 22244 12316
rect 22190 12200 22246 12209
rect 22190 12135 22246 12144
rect 22204 12102 22232 12135
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 10606 22232 12038
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22296 11354 22324 11494
rect 22480 11354 22508 11698
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21928 9586 21956 9862
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21744 8566 21772 8978
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21086 8120 21142 8129
rect 21086 8055 21142 8064
rect 21100 7449 21128 8055
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 21284 7721 21312 7890
rect 21744 7886 21772 8502
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21270 7712 21326 7721
rect 21270 7647 21326 7656
rect 21284 7546 21312 7647
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21086 7440 21142 7449
rect 21744 7410 21772 7822
rect 21836 7546 21864 9318
rect 21928 8362 21956 9522
rect 22296 8537 22324 11290
rect 22664 8922 22692 13194
rect 22744 11280 22796 11286
rect 22744 11222 22796 11228
rect 22756 10742 22784 11222
rect 22744 10736 22796 10742
rect 22742 10704 22744 10713
rect 22796 10704 22798 10713
rect 22742 10639 22798 10648
rect 22756 10130 22784 10639
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22572 8894 22692 8922
rect 22282 8528 22338 8537
rect 22282 8463 22338 8472
rect 22282 8392 22338 8401
rect 21916 8356 21968 8362
rect 22282 8327 22338 8336
rect 21916 8298 21968 8304
rect 22190 8120 22246 8129
rect 22296 8090 22324 8327
rect 22190 8055 22246 8064
rect 22284 8084 22336 8090
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21086 7375 21142 7384
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21192 7002 21220 7346
rect 21836 7274 21864 7482
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 20996 6248 21048 6254
rect 20718 6216 20774 6225
rect 20996 6190 21048 6196
rect 21100 6186 21128 6802
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21284 6662 21312 6734
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21284 6390 21312 6598
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 20718 6151 20774 6160
rect 21088 6180 21140 6186
rect 20732 5914 20760 6151
rect 21088 6122 21140 6128
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19706 4584 19762 4593
rect 19706 4519 19762 4528
rect 19720 4146 19748 4519
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19614 3632 19670 3641
rect 19614 3567 19616 3576
rect 19668 3567 19670 3576
rect 19616 3538 19668 3544
rect 19628 3194 19656 3538
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 20088 2825 20116 5510
rect 20180 5098 20208 5510
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 20180 4622 20208 5034
rect 20916 4690 20944 5510
rect 21100 5273 21128 6122
rect 21468 5914 21496 6190
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21652 5710 21680 6122
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21086 5264 21142 5273
rect 21086 5199 21142 5208
rect 21376 4826 21404 5646
rect 21652 5370 21680 5646
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 21640 5364 21692 5370
rect 21640 5306 21692 5312
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21086 4720 21142 4729
rect 20904 4684 20956 4690
rect 21086 4655 21142 4664
rect 20904 4626 20956 4632
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20916 4282 20944 4626
rect 21100 4622 21128 4655
rect 22112 4622 22140 5510
rect 22204 5370 22232 8055
rect 22284 8026 22336 8032
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22296 5574 22324 6598
rect 22466 5808 22522 5817
rect 22466 5743 22468 5752
rect 22520 5743 22522 5752
rect 22468 5714 22520 5720
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22480 5370 22508 5714
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22572 4826 22600 8894
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22664 8430 22692 8774
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20272 3398 20300 4082
rect 21822 4040 21878 4049
rect 21822 3975 21824 3984
rect 21876 3975 21878 3984
rect 22006 4040 22062 4049
rect 22006 3975 22062 3984
rect 21824 3946 21876 3952
rect 22020 3942 22048 3975
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 20364 3738 20392 3878
rect 22112 3754 22140 4558
rect 22572 4010 22600 4762
rect 22664 4185 22692 4966
rect 22650 4176 22706 4185
rect 22650 4111 22706 4120
rect 22560 4004 22612 4010
rect 22560 3946 22612 3952
rect 22572 3777 22600 3946
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 21928 3726 22140 3754
rect 21928 3618 21956 3726
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 21744 3590 21956 3618
rect 22008 3596 22060 3602
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20272 2922 20300 3334
rect 20364 3058 20392 3538
rect 21744 3534 21772 3590
rect 22008 3538 22060 3544
rect 21732 3528 21784 3534
rect 20442 3496 20498 3505
rect 21732 3470 21784 3476
rect 20442 3431 20498 3440
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20364 2961 20392 2994
rect 20350 2952 20406 2961
rect 20260 2916 20312 2922
rect 20350 2887 20406 2896
rect 20260 2858 20312 2864
rect 20074 2816 20130 2825
rect 19622 2748 19918 2768
rect 20074 2751 20130 2760
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20272 2650 20300 2858
rect 20456 2650 20484 3431
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21560 3097 21588 3334
rect 21546 3088 21602 3097
rect 21546 3023 21602 3032
rect 21744 2990 21772 3470
rect 22020 3194 22048 3538
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 21914 3088 21970 3097
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 21836 2650 21864 3062
rect 21914 3023 21970 3032
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21928 2582 21956 3023
rect 21916 2576 21968 2582
rect 20902 2544 20958 2553
rect 21916 2518 21968 2524
rect 20902 2479 20904 2488
rect 20956 2479 20958 2488
rect 20904 2450 20956 2456
rect 22020 2446 22048 3130
rect 22112 2650 22140 3726
rect 22558 3768 22614 3777
rect 22558 3703 22614 3712
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22388 3194 22416 3334
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22098 2408 22154 2417
rect 22098 2343 22154 2352
rect 20718 2000 20774 2009
rect 20718 1935 20774 1944
rect 19536 1414 20116 1442
rect 20088 480 20116 1414
rect 20732 480 20760 1935
rect 21362 1592 21418 1601
rect 21362 1527 21418 1536
rect 21376 480 21404 1527
rect 22112 480 22140 2343
rect 22756 480 22784 7142
rect 22848 4282 22876 19314
rect 23032 18222 23060 20198
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22940 17134 22968 17614
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22940 16250 22968 16526
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22940 16046 22968 16186
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 23032 15892 23060 18022
rect 22940 15864 23060 15892
rect 22940 13433 22968 15864
rect 23020 15564 23072 15570
rect 23020 15506 23072 15512
rect 23032 15094 23060 15506
rect 23020 15088 23072 15094
rect 23020 15030 23072 15036
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 23032 13870 23060 14486
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22926 13424 22982 13433
rect 22926 13359 22982 13368
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22940 12986 22968 13262
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22940 12442 22968 12718
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22940 11558 22968 11630
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 22940 6118 22968 11494
rect 23032 10985 23060 13806
rect 23124 12850 23152 24550
rect 23308 23866 23336 26007
rect 23400 24410 23428 26551
rect 23492 25226 23520 27520
rect 23768 26858 23796 27639
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25502 27520 25558 28000
rect 26146 27520 26202 28000
rect 26882 27520 26938 28000
rect 27526 27520 27582 28000
rect 23756 26852 23808 26858
rect 23756 26794 23808 26800
rect 23662 25392 23718 25401
rect 23662 25327 23718 25336
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23676 24410 23704 25327
rect 24136 24426 24164 27520
rect 24780 27282 24808 27520
rect 24688 27254 24808 27282
rect 24688 25430 24716 27254
rect 24766 27160 24822 27169
rect 24766 27095 24822 27104
rect 24780 26654 24808 27095
rect 24768 26648 24820 26654
rect 24768 26590 24820 26596
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24216 25356 24268 25362
rect 24216 25298 24268 25304
rect 24228 24614 24256 25298
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24780 24857 24808 25094
rect 24766 24848 24822 24857
rect 24766 24783 24822 24792
rect 24584 24744 24636 24750
rect 25516 24721 25544 27520
rect 26160 25294 26188 27520
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 24584 24686 24636 24692
rect 25502 24712 25558 24721
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 24044 24398 24164 24426
rect 23754 24304 23810 24313
rect 23480 24268 23532 24274
rect 23754 24239 23810 24248
rect 23480 24210 23532 24216
rect 23492 23866 23520 24210
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23478 23760 23534 23769
rect 23478 23695 23534 23704
rect 23492 23338 23520 23695
rect 23400 23322 23520 23338
rect 23388 23316 23520 23322
rect 23440 23310 23520 23316
rect 23388 23258 23440 23264
rect 23768 23089 23796 24239
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 23754 23080 23810 23089
rect 23754 23015 23810 23024
rect 23754 22944 23810 22953
rect 23754 22879 23810 22888
rect 23294 22808 23350 22817
rect 23294 22743 23350 22752
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23216 17814 23244 18906
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23216 17338 23244 17750
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23308 17082 23336 22743
rect 23664 20392 23716 20398
rect 23662 20360 23664 20369
rect 23716 20360 23718 20369
rect 23662 20295 23718 20304
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23492 19417 23520 19722
rect 23676 19553 23704 20198
rect 23662 19544 23718 19553
rect 23662 19479 23718 19488
rect 23478 19408 23534 19417
rect 23478 19343 23534 19352
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23570 17640 23626 17649
rect 23570 17575 23626 17584
rect 23216 17054 23336 17082
rect 23216 16114 23244 17054
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 23110 12336 23166 12345
rect 23110 12271 23112 12280
rect 23164 12271 23166 12280
rect 23112 12242 23164 12248
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 23018 10976 23074 10985
rect 23018 10911 23074 10920
rect 23124 10266 23152 11222
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23032 8809 23060 9318
rect 23124 9178 23152 10202
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23018 8800 23074 8809
rect 23018 8735 23074 8744
rect 23216 8514 23244 16050
rect 23308 15994 23336 16934
rect 23478 16824 23534 16833
rect 23478 16759 23534 16768
rect 23492 16266 23520 16759
rect 23584 16522 23612 17575
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23400 16238 23520 16266
rect 23584 16250 23612 16458
rect 23676 16289 23704 19246
rect 23662 16280 23718 16289
rect 23572 16244 23624 16250
rect 23400 16182 23428 16238
rect 23662 16215 23718 16224
rect 23572 16186 23624 16192
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23308 15966 23704 15994
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23308 14414 23336 15302
rect 23492 15178 23520 15370
rect 23400 15162 23520 15178
rect 23388 15156 23520 15162
rect 23440 15150 23520 15156
rect 23388 15098 23440 15104
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23308 13938 23336 14350
rect 23400 14074 23428 14554
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23388 14068 23440 14074
rect 23440 14028 23520 14056
rect 23388 14010 23440 14016
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23308 13530 23336 13874
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12782 23428 13126
rect 23492 12850 23520 14028
rect 23584 13326 23612 14214
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23676 13002 23704 15966
rect 23768 14550 23796 22879
rect 23848 22432 23900 22438
rect 23952 22386 23980 23122
rect 24044 22681 24072 24398
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24136 23526 24164 24210
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 24030 22672 24086 22681
rect 24030 22607 24086 22616
rect 23900 22380 23980 22386
rect 23848 22374 23980 22380
rect 23860 22358 23980 22374
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23860 22001 23888 22034
rect 23846 21992 23902 22001
rect 23846 21927 23902 21936
rect 23860 21690 23888 21927
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23952 21570 23980 22358
rect 23860 21542 23980 21570
rect 23860 15978 23888 21542
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23952 16794 23980 21422
rect 24030 21176 24086 21185
rect 24030 21111 24032 21120
rect 24084 21111 24086 21120
rect 24032 21082 24084 21088
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 24044 20641 24072 20878
rect 24030 20632 24086 20641
rect 24030 20567 24086 20576
rect 24044 20210 24072 20567
rect 24136 20505 24164 23462
rect 24228 22642 24256 24550
rect 24596 24177 24624 24686
rect 25502 24647 25558 24656
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24582 24168 24638 24177
rect 24582 24103 24638 24112
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24688 22522 24716 24006
rect 24780 23225 24808 24550
rect 25870 24304 25926 24313
rect 25870 24239 25926 24248
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 24766 23216 24822 23225
rect 24766 23151 24822 23160
rect 24872 23066 24900 23462
rect 25226 23352 25282 23361
rect 25226 23287 25282 23296
rect 25240 23254 25268 23287
rect 25228 23248 25280 23254
rect 25228 23190 25280 23196
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 24228 22494 24716 22522
rect 24780 23038 24900 23066
rect 24228 21457 24256 22494
rect 24400 22432 24452 22438
rect 24398 22400 24400 22409
rect 24452 22400 24454 22409
rect 24780 22386 24808 23038
rect 25056 22778 25084 23122
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 25056 22658 25084 22714
rect 25056 22630 25176 22658
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 24398 22335 24454 22344
rect 24596 22358 24808 22386
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24596 21962 24624 22358
rect 24872 22250 24900 22374
rect 24688 22222 24900 22250
rect 24952 22228 25004 22234
rect 24688 21978 24716 22222
rect 24952 22170 25004 22176
rect 24766 22128 24822 22137
rect 24964 22114 24992 22170
rect 25056 22137 25084 22510
rect 25148 22234 25176 22630
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 24766 22063 24768 22072
rect 24820 22063 24822 22072
rect 24872 22086 24992 22114
rect 25042 22128 25098 22137
rect 24768 22034 24820 22040
rect 24584 21956 24636 21962
rect 24688 21950 24808 21978
rect 24584 21898 24636 21904
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24214 21448 24270 21457
rect 24214 21383 24270 21392
rect 24492 21412 24544 21418
rect 24492 21354 24544 21360
rect 24504 21049 24532 21354
rect 24688 21049 24716 21830
rect 24490 21040 24546 21049
rect 24490 20975 24546 20984
rect 24674 21040 24730 21049
rect 24674 20975 24730 20984
rect 24216 20936 24268 20942
rect 24780 20890 24808 21950
rect 24216 20878 24268 20884
rect 24228 20806 24256 20878
rect 24688 20862 24808 20890
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24122 20496 24178 20505
rect 24122 20431 24178 20440
rect 24044 20182 24164 20210
rect 24136 20058 24164 20182
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24044 19378 24072 19994
rect 24228 19922 24256 20742
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24584 20392 24636 20398
rect 24688 20369 24716 20862
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24584 20334 24636 20340
rect 24674 20360 24730 20369
rect 24216 19916 24268 19922
rect 24216 19858 24268 19864
rect 24596 19854 24624 20334
rect 24674 20295 24730 20304
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 24044 18834 24072 19314
rect 24124 19168 24176 19174
rect 24124 19110 24176 19116
rect 24136 18873 24164 19110
rect 24122 18864 24178 18873
rect 24032 18828 24084 18834
rect 24122 18799 24178 18808
rect 24032 18770 24084 18776
rect 24044 18290 24072 18770
rect 24216 18692 24268 18698
rect 24216 18634 24268 18640
rect 24122 18456 24178 18465
rect 24122 18391 24124 18400
rect 24176 18391 24178 18400
rect 24124 18362 24176 18368
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24044 17066 24072 17818
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23938 16552 23994 16561
rect 23938 16487 23994 16496
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23846 14648 23902 14657
rect 23846 14583 23902 14592
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23768 14074 23796 14486
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23860 13161 23888 14583
rect 23952 14482 23980 16487
rect 24044 16114 24072 17002
rect 24136 16726 24164 17002
rect 24228 16794 24256 18634
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18170 24716 19450
rect 24780 19145 24808 20742
rect 24766 19136 24822 19145
rect 24766 19071 24822 19080
rect 24688 18142 24808 18170
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24780 16969 24808 18142
rect 24766 16960 24822 16969
rect 24766 16895 24822 16904
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24124 16720 24176 16726
rect 24124 16662 24176 16668
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 24228 16250 24256 16526
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24216 15972 24268 15978
rect 24216 15914 24268 15920
rect 24122 15736 24178 15745
rect 24122 15671 24178 15680
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23846 13152 23902 13161
rect 23846 13087 23902 13096
rect 23676 12974 23888 13002
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23308 11218 23336 12310
rect 23400 12238 23428 12718
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23400 11626 23428 12174
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23400 11286 23428 11562
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23492 10826 23520 12106
rect 23032 8486 23244 8514
rect 23308 10798 23520 10826
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 23032 5409 23060 8486
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 23216 7750 23244 8366
rect 23308 8265 23336 10798
rect 23478 9616 23534 9625
rect 23478 9551 23534 9560
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23400 9194 23428 9454
rect 23492 9382 23520 9551
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23400 9166 23520 9194
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23400 8362 23428 8978
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23294 8256 23350 8265
rect 23294 8191 23350 8200
rect 23400 7970 23428 8298
rect 23492 8129 23520 9166
rect 23478 8120 23534 8129
rect 23478 8055 23534 8064
rect 23400 7942 23520 7970
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23216 7342 23244 7686
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 23124 6458 23152 6734
rect 23216 6662 23244 7278
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 5914 23152 6394
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 23124 5681 23152 5714
rect 23110 5672 23166 5681
rect 23110 5607 23166 5616
rect 23018 5400 23074 5409
rect 23124 5370 23152 5607
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23018 5335 23074 5344
rect 23112 5364 23164 5370
rect 23032 4865 23060 5335
rect 23112 5306 23164 5312
rect 23216 5234 23244 5510
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 23018 4856 23074 4865
rect 23018 4791 23074 4800
rect 23020 4684 23072 4690
rect 23020 4626 23072 4632
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 23032 3942 23060 4626
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23032 3466 23060 3878
rect 23308 3670 23336 7822
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23296 3664 23348 3670
rect 23296 3606 23348 3612
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23124 3194 23152 3470
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23400 2922 23428 7142
rect 23492 4282 23520 7942
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23584 4078 23612 12582
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23492 3194 23520 3878
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23388 2916 23440 2922
rect 23388 2858 23440 2864
rect 23478 2816 23534 2825
rect 23478 2751 23534 2760
rect 23492 480 23520 2751
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2318 0 2374 480
rect 2962 0 3018 480
rect 3698 0 3754 480
rect 4342 0 4398 480
rect 4986 0 5042 480
rect 5722 0 5778 480
rect 6366 0 6422 480
rect 7102 0 7158 480
rect 7746 0 7802 480
rect 8390 0 8446 480
rect 9126 0 9182 480
rect 9770 0 9826 480
rect 10506 0 10562 480
rect 11150 0 11206 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13174 0 13230 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15290 0 15346 480
rect 15934 0 15990 480
rect 16578 0 16634 480
rect 17314 0 17370 480
rect 17958 0 18014 480
rect 18694 0 18750 480
rect 19338 0 19394 480
rect 20074 0 20130 480
rect 20718 0 20774 480
rect 21362 0 21418 480
rect 22098 0 22154 480
rect 22742 0 22798 480
rect 23478 0 23534 480
rect 23676 377 23704 12854
rect 23756 12708 23808 12714
rect 23756 12650 23808 12656
rect 23768 12481 23796 12650
rect 23754 12472 23810 12481
rect 23754 12407 23810 12416
rect 23768 12102 23796 12407
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23768 11354 23796 12038
rect 23860 11937 23888 12974
rect 23952 12889 23980 13806
rect 24136 13569 24164 15671
rect 24122 13560 24178 13569
rect 24122 13495 24178 13504
rect 24032 13456 24084 13462
rect 24032 13398 24084 13404
rect 24122 13424 24178 13433
rect 24044 12986 24072 13398
rect 24122 13359 24178 13368
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 23938 12880 23994 12889
rect 23938 12815 23994 12824
rect 23846 11928 23902 11937
rect 23846 11863 23902 11872
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23860 10198 23888 11630
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 23860 9586 23888 10134
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23846 8936 23902 8945
rect 23846 8871 23902 8880
rect 23860 8537 23888 8871
rect 23952 8634 23980 12815
rect 24136 12170 24164 13359
rect 24228 12646 24256 15914
rect 24412 15706 24440 16050
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 14958 24716 15642
rect 24780 15366 24808 15846
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24766 15192 24822 15201
rect 24766 15127 24822 15136
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24400 14884 24452 14890
rect 24400 14826 24452 14832
rect 24412 14346 24440 14826
rect 24400 14340 24452 14346
rect 24400 14282 24452 14288
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12730 24808 15127
rect 24872 13716 24900 22086
rect 25424 22098 25452 23462
rect 25502 23080 25558 23089
rect 25502 23015 25558 23024
rect 25042 22063 25098 22072
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 25148 21622 25176 22034
rect 25136 21616 25188 21622
rect 25134 21584 25136 21593
rect 25188 21584 25190 21593
rect 25134 21519 25190 21528
rect 25516 21486 25544 23015
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25042 21176 25098 21185
rect 25042 21111 25098 21120
rect 24952 20868 25004 20874
rect 24952 20810 25004 20816
rect 24964 20398 24992 20810
rect 25056 20602 25084 21111
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25240 20602 25268 20946
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24964 20058 24992 20334
rect 25240 20233 25268 20538
rect 25410 20496 25466 20505
rect 25410 20431 25412 20440
rect 25464 20431 25466 20440
rect 25412 20402 25464 20408
rect 25226 20224 25282 20233
rect 25226 20159 25282 20168
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 25320 19984 25372 19990
rect 25320 19926 25372 19932
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 24964 19514 24992 19858
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 25228 19304 25280 19310
rect 25226 19272 25228 19281
rect 25280 19272 25282 19281
rect 25226 19207 25282 19216
rect 25240 18970 25268 19207
rect 25332 19174 25360 19926
rect 25700 19689 25728 21286
rect 25686 19680 25742 19689
rect 25686 19615 25742 19624
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 25044 18896 25096 18902
rect 25044 18838 25096 18844
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24964 18426 24992 18702
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25056 18086 25084 18838
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17921 25084 18022
rect 25042 17912 25098 17921
rect 25148 17882 25176 18702
rect 25228 18216 25280 18222
rect 25226 18184 25228 18193
rect 25280 18184 25282 18193
rect 25226 18119 25282 18128
rect 25332 17898 25360 19110
rect 25516 19009 25544 19178
rect 25502 19000 25558 19009
rect 25502 18935 25558 18944
rect 25594 18864 25650 18873
rect 25594 18799 25650 18808
rect 25412 18080 25464 18086
rect 25410 18048 25412 18057
rect 25464 18048 25466 18057
rect 25410 17983 25466 17992
rect 25042 17847 25098 17856
rect 25136 17876 25188 17882
rect 25332 17870 25452 17898
rect 25136 17818 25188 17824
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 25240 17252 25268 17682
rect 25320 17536 25372 17542
rect 25318 17504 25320 17513
rect 25372 17504 25374 17513
rect 25318 17439 25374 17448
rect 25320 17264 25372 17270
rect 25240 17232 25320 17252
rect 25372 17232 25374 17241
rect 25240 17224 25318 17232
rect 25318 17167 25374 17176
rect 25424 17105 25452 17870
rect 25410 17096 25466 17105
rect 25410 17031 25466 17040
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 24964 16182 24992 16730
rect 25056 16658 25084 16934
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 25056 15706 25084 16390
rect 25608 16114 25636 18799
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24964 14618 24992 15506
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25056 14890 25084 15438
rect 25148 15162 25176 15438
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 25056 14074 25084 14826
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 25148 13954 25176 14214
rect 25056 13926 25176 13954
rect 25240 13938 25268 14350
rect 25608 14074 25636 14418
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25228 13932 25280 13938
rect 25056 13870 25084 13926
rect 25228 13874 25280 13880
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25044 13864 25096 13870
rect 25042 13832 25044 13841
rect 25096 13832 25098 13841
rect 25042 13767 25098 13776
rect 24872 13688 25084 13716
rect 24596 12702 24808 12730
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24596 12209 24624 12702
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24582 12200 24638 12209
rect 24124 12164 24176 12170
rect 24582 12135 24638 12144
rect 24124 12106 24176 12112
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24136 11529 24164 11698
rect 24216 11552 24268 11558
rect 24122 11520 24178 11529
rect 24216 11494 24268 11500
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24122 11455 24178 11464
rect 24228 10606 24256 11494
rect 24596 11082 24624 11494
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24216 10600 24268 10606
rect 24122 10568 24178 10577
rect 24216 10542 24268 10548
rect 24122 10503 24178 10512
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23846 8528 23902 8537
rect 23846 8463 23902 8472
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 23768 7002 23796 7890
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23768 6458 23796 6938
rect 23860 6769 23888 8463
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 23846 6760 23902 6769
rect 23846 6695 23902 6704
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23754 6352 23810 6361
rect 23754 6287 23810 6296
rect 23768 6186 23796 6287
rect 23756 6180 23808 6186
rect 23756 6122 23808 6128
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 23768 4486 23796 5034
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 4214 23796 4422
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23860 4146 23888 6598
rect 23952 6322 23980 7210
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23768 1465 23796 4014
rect 23860 3738 23888 4082
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 23860 3194 23888 3538
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23952 2394 23980 5578
rect 24044 3516 24072 10406
rect 24136 9897 24164 10503
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24122 9888 24178 9897
rect 24122 9823 24178 9832
rect 24228 9722 24256 10406
rect 24320 10266 24348 10610
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 24124 8560 24176 8566
rect 24124 8502 24176 8508
rect 24136 5930 24164 8502
rect 24228 8265 24256 9318
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24214 8256 24270 8265
rect 24214 8191 24270 8200
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24228 6458 24256 6802
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24136 5902 24256 5930
rect 24124 5840 24176 5846
rect 24124 5782 24176 5788
rect 24136 4486 24164 5782
rect 24124 4480 24176 4486
rect 24122 4448 24124 4457
rect 24176 4448 24178 4457
rect 24122 4383 24178 4392
rect 24122 4176 24178 4185
rect 24122 4111 24178 4120
rect 24136 3618 24164 4111
rect 24228 4010 24256 5902
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 4826 24716 12582
rect 24860 12368 24912 12374
rect 24766 12336 24822 12345
rect 24860 12310 24912 12316
rect 24766 12271 24822 12280
rect 24780 11762 24808 12271
rect 24872 11898 24900 12310
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24872 11354 24900 11834
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24766 9480 24822 9489
rect 24766 9415 24822 9424
rect 24780 7993 24808 9415
rect 25056 8616 25084 13688
rect 25318 13288 25374 13297
rect 25318 13223 25374 13232
rect 25228 13184 25280 13190
rect 25228 13126 25280 13132
rect 25240 12374 25268 13126
rect 25228 12368 25280 12374
rect 25228 12310 25280 12316
rect 25332 12220 25360 13223
rect 25608 12442 25636 13874
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25240 12192 25360 12220
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25148 9178 25176 9522
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 24964 8588 25084 8616
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24872 8090 24900 8298
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24766 7984 24822 7993
rect 24766 7919 24822 7928
rect 24766 7440 24822 7449
rect 24766 7375 24822 7384
rect 24780 6633 24808 7375
rect 24766 6624 24822 6633
rect 24766 6559 24822 6568
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24768 5296 24820 5302
rect 24766 5264 24768 5273
rect 24820 5264 24822 5273
rect 24766 5199 24822 5208
rect 24872 5030 24900 5714
rect 24860 5024 24912 5030
rect 24780 4972 24860 4978
rect 24780 4966 24912 4972
rect 24780 4950 24900 4966
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24228 3738 24256 3946
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24136 3590 24256 3618
rect 24044 3488 24164 3516
rect 24136 2514 24164 3488
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24228 2394 24256 3590
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3470
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24780 3074 24808 4950
rect 24858 4856 24914 4865
rect 24858 4791 24914 4800
rect 24688 3046 24808 3074
rect 24582 2952 24638 2961
rect 24582 2887 24638 2896
rect 24596 2553 24624 2887
rect 24688 2582 24716 3046
rect 24872 2990 24900 4791
rect 24964 3398 24992 8588
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 25056 7954 25084 8434
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 25056 7546 25084 7890
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 25148 5642 25176 6258
rect 25136 5636 25188 5642
rect 25136 5578 25188 5584
rect 25148 5370 25176 5578
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 25056 4622 25084 5238
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 25044 4616 25096 4622
rect 25044 4558 25096 4564
rect 25056 4282 25084 4558
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24676 2576 24728 2582
rect 24582 2544 24638 2553
rect 24676 2518 24728 2524
rect 25148 2514 25176 5170
rect 25240 4078 25268 12192
rect 25884 11354 25912 24239
rect 26896 23633 26924 27520
rect 26882 23624 26938 23633
rect 26882 23559 26938 23568
rect 27540 20097 27568 27520
rect 27526 20088 27582 20097
rect 27526 20023 27582 20032
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 25976 19514 26004 19790
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26056 15360 26108 15366
rect 26056 15302 26108 15308
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25780 11212 25832 11218
rect 25780 11154 25832 11160
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25332 10674 25360 10950
rect 25792 10810 25820 11154
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25424 8430 25452 9318
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 25332 4865 25360 6054
rect 25318 4856 25374 4865
rect 25424 4826 25452 6734
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25318 4791 25374 4800
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25228 4072 25280 4078
rect 25332 4049 25360 4626
rect 25424 4214 25452 4762
rect 25412 4208 25464 4214
rect 25412 4150 25464 4156
rect 25228 4014 25280 4020
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 25332 3738 25360 3975
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 24582 2479 24638 2488
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 23952 2366 24164 2394
rect 24228 2366 24808 2394
rect 23754 1456 23810 1465
rect 23754 1391 23810 1400
rect 24136 480 24164 2366
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24780 480 24808 2366
rect 25516 480 25544 5510
rect 26068 4321 26096 15302
rect 26160 15178 26188 15506
rect 26160 15162 26280 15178
rect 26160 15156 26292 15162
rect 26160 15150 26240 15156
rect 26240 15098 26292 15104
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26160 10130 26188 10406
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 26054 4312 26110 4321
rect 26054 4247 26110 4256
rect 26148 4004 26200 4010
rect 26148 3946 26200 3952
rect 26160 480 26188 3946
rect 26884 3120 26936 3126
rect 26884 3062 26936 3068
rect 26896 480 26924 3062
rect 27528 2372 27580 2378
rect 27528 2314 27580 2320
rect 27540 480 27568 2314
rect 23662 368 23718 377
rect 23662 303 23718 312
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25502 0 25558 480
rect 26146 0 26202 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 23754 27648 23810 27704
rect 938 24384 994 24440
rect 386 11600 442 11656
rect 3698 23704 3754 23760
rect 2962 21936 3018 21992
rect 4066 20984 4122 21040
rect 1582 18128 1638 18184
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5998 24792 6054 24848
rect 5998 24384 6054 24440
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 4986 22616 5042 22672
rect 6090 23704 6146 23760
rect 5998 22480 6054 22536
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 7746 23840 7802 23896
rect 9126 24112 9182 24168
rect 7102 23432 7158 23488
rect 6366 23160 6422 23216
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10138 23432 10194 23488
rect 9770 21664 9826 21720
rect 6090 21528 6146 21584
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 11610 23568 11666 23624
rect 11150 23432 11206 23488
rect 11150 23296 11206 23352
rect 10690 23024 10746 23080
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10230 21392 10286 21448
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 9402 20712 9458 20768
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 9770 20460 9826 20496
rect 9770 20440 9772 20460
rect 9772 20440 9824 20460
rect 9824 20440 9826 20460
rect 9770 19760 9826 19816
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4342 18808 4398 18864
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 8206 16224 8262 16280
rect 4066 15408 4122 15464
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 1398 10104 1454 10160
rect 4986 10104 5042 10160
rect 294 8064 350 8120
rect 3698 7792 3754 7848
rect 2318 7248 2374 7304
rect 938 4120 994 4176
rect 1582 2488 1638 2544
rect 2962 4528 3018 4584
rect 4342 3576 4398 3632
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 7102 3984 7158 4040
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6366 3032 6422 3088
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5722 1808 5778 1864
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10230 19252 10232 19272
rect 10232 19252 10284 19272
rect 10284 19252 10286 19272
rect 10230 19216 10286 19252
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 9954 16496 10010 16552
rect 11610 21256 11666 21312
rect 11242 19352 11298 19408
rect 11426 18692 11482 18728
rect 11426 18672 11428 18692
rect 11428 18672 11480 18692
rect 11480 18672 11482 18692
rect 11426 18164 11428 18184
rect 11428 18164 11480 18184
rect 11480 18164 11482 18184
rect 11426 18128 11482 18164
rect 10874 16788 10930 16824
rect 10874 16768 10876 16788
rect 10876 16768 10928 16788
rect 10928 16768 10930 16788
rect 10874 16632 10930 16688
rect 10690 15816 10746 15872
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10046 15272 10102 15328
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10138 14184 10194 14240
rect 9954 9968 10010 10024
rect 9770 7656 9826 7712
rect 8390 3304 8446 3360
rect 8758 1536 8814 1592
rect 9218 1672 9274 1728
rect 9862 6860 9918 6896
rect 9862 6840 9864 6860
rect 9864 6840 9916 6860
rect 9916 6840 9918 6860
rect 10782 14048 10838 14104
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10782 10240 10838 10296
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 11242 12588 11244 12608
rect 11244 12588 11296 12608
rect 11296 12588 11298 12608
rect 11242 12552 11298 12588
rect 10966 12144 11022 12200
rect 11058 11600 11114 11656
rect 11150 9324 11152 9344
rect 11152 9324 11204 9344
rect 11204 9324 11206 9344
rect 11150 9288 11206 9324
rect 10690 8336 10746 8392
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10322 7268 10378 7304
rect 10322 7248 10324 7268
rect 10324 7248 10376 7268
rect 10376 7248 10378 7268
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 11426 15020 11482 15056
rect 11426 15000 11428 15020
rect 11428 15000 11480 15020
rect 11480 15000 11482 15020
rect 11702 18828 11758 18864
rect 11702 18808 11704 18828
rect 11704 18808 11756 18828
rect 11756 18808 11758 18828
rect 12070 23860 12126 23896
rect 12070 23840 12072 23860
rect 12072 23840 12124 23860
rect 12124 23840 12126 23860
rect 11978 22072 12034 22128
rect 11978 17176 12034 17232
rect 12806 24792 12862 24848
rect 12530 23840 12586 23896
rect 12438 23432 12494 23488
rect 12346 23160 12402 23216
rect 12438 20712 12494 20768
rect 12346 20032 12402 20088
rect 12254 18028 12256 18048
rect 12256 18028 12308 18048
rect 12308 18028 12310 18048
rect 12254 17992 12310 18028
rect 13726 24656 13782 24712
rect 13174 23568 13230 23624
rect 13174 21392 13230 21448
rect 12622 17604 12678 17640
rect 12622 17584 12624 17604
rect 12624 17584 12676 17604
rect 12676 17584 12678 17604
rect 12162 16632 12218 16688
rect 11518 13640 11574 13696
rect 12254 14592 12310 14648
rect 11886 9968 11942 10024
rect 12162 11736 12218 11792
rect 12898 14864 12954 14920
rect 12254 11328 12310 11384
rect 12070 10104 12126 10160
rect 12254 10104 12310 10160
rect 12254 9832 12310 9888
rect 11426 8200 11482 8256
rect 11242 7792 11298 7848
rect 11610 9152 11666 9208
rect 11058 6976 11114 7032
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10690 4936 10746 4992
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10046 3984 10102 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10506 1400 10562 1456
rect 10966 2760 11022 2816
rect 10874 2624 10930 2680
rect 12346 9016 12402 9072
rect 11794 8200 11850 8256
rect 12438 8336 12494 8392
rect 11978 8064 12034 8120
rect 11794 6976 11850 7032
rect 11886 6840 11942 6896
rect 11702 6296 11758 6352
rect 11794 4564 11796 4584
rect 11796 4564 11848 4584
rect 11848 4564 11850 4584
rect 11794 4528 11850 4564
rect 11886 3884 11888 3904
rect 11888 3884 11940 3904
rect 11940 3884 11942 3904
rect 11886 3848 11942 3884
rect 11426 3712 11482 3768
rect 12622 8200 12678 8256
rect 12530 7656 12586 7712
rect 12070 6024 12126 6080
rect 12438 6704 12494 6760
rect 11978 3576 12034 3632
rect 11426 3460 11482 3496
rect 11426 3440 11428 3460
rect 11428 3440 11480 3460
rect 11480 3440 11482 3460
rect 11886 3168 11942 3224
rect 11426 2896 11482 2952
rect 11610 1944 11666 2000
rect 12806 4684 12862 4720
rect 12806 4664 12808 4684
rect 12808 4664 12860 4684
rect 12860 4664 12862 4684
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14554 24792 14610 24848
rect 13910 24384 13966 24440
rect 13450 20984 13506 21040
rect 13450 17040 13506 17096
rect 13634 16904 13690 16960
rect 14278 24248 14334 24304
rect 14002 20848 14058 20904
rect 13910 20032 13966 20088
rect 13818 19896 13874 19952
rect 13818 19352 13874 19408
rect 13818 19216 13874 19272
rect 13726 16224 13782 16280
rect 13542 15544 13598 15600
rect 13542 15308 13544 15328
rect 13544 15308 13596 15328
rect 13596 15308 13598 15328
rect 13542 15272 13598 15308
rect 13450 14220 13452 14240
rect 13452 14220 13504 14240
rect 13504 14220 13506 14240
rect 13450 14184 13506 14220
rect 13450 9560 13506 9616
rect 13266 4800 13322 4856
rect 13082 3304 13138 3360
rect 13450 6160 13506 6216
rect 13634 11056 13690 11112
rect 14094 19318 14150 19374
rect 14002 14592 14058 14648
rect 14922 24248 14978 24304
rect 14738 23840 14794 23896
rect 14554 22480 14610 22536
rect 14370 21528 14426 21584
rect 14278 18400 14334 18456
rect 14370 18128 14426 18184
rect 15934 24112 15990 24168
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15290 22616 15346 22672
rect 14738 22480 14794 22536
rect 14646 22092 14702 22128
rect 14646 22072 14648 22092
rect 14648 22072 14700 22092
rect 14700 22072 14702 22092
rect 14830 22072 14886 22128
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15566 21972 15568 21992
rect 15568 21972 15620 21992
rect 15620 21972 15622 21992
rect 15566 21936 15622 21972
rect 15474 21528 15530 21584
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14554 18264 14610 18320
rect 14462 16788 14518 16824
rect 14462 16768 14464 16788
rect 14464 16768 14516 16788
rect 14516 16768 14518 16788
rect 14186 13776 14242 13832
rect 14462 13504 14518 13560
rect 14738 17756 14740 17776
rect 14740 17756 14792 17776
rect 14792 17756 14794 17776
rect 14738 17720 14794 17756
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15014 18128 15070 18184
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14830 15952 14886 16008
rect 14738 15680 14794 15736
rect 14646 14068 14702 14104
rect 14646 14048 14648 14068
rect 14648 14048 14700 14068
rect 14700 14048 14702 14068
rect 13910 11600 13966 11656
rect 13726 10376 13782 10432
rect 13910 9560 13966 9616
rect 13358 3032 13414 3088
rect 12898 2372 12954 2408
rect 12898 2352 12900 2372
rect 12900 2352 12952 2372
rect 12952 2352 12954 2372
rect 13726 7792 13782 7848
rect 14002 8472 14058 8528
rect 13818 6432 13874 6488
rect 13726 5616 13782 5672
rect 14094 6432 14150 6488
rect 14462 11600 14518 11656
rect 14646 13232 14702 13288
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15658 15816 15714 15872
rect 15566 15036 15568 15056
rect 15568 15036 15620 15056
rect 15620 15036 15622 15056
rect 15566 15000 15622 15036
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15106 13932 15162 13968
rect 15106 13912 15108 13932
rect 15108 13912 15160 13932
rect 15160 13912 15162 13932
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14278 8336 14334 8392
rect 14370 8064 14426 8120
rect 14094 4936 14150 4992
rect 15566 13096 15622 13152
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15382 12008 15438 12064
rect 15014 11076 15070 11112
rect 15014 11056 15016 11076
rect 15016 11056 15068 11076
rect 15068 11056 15070 11076
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15014 10240 15070 10296
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15934 22480 15990 22536
rect 15934 19760 15990 19816
rect 16210 24404 16266 24440
rect 16210 24384 16212 24404
rect 16212 24384 16264 24404
rect 16264 24384 16266 24404
rect 16118 19488 16174 19544
rect 16670 19352 16726 19408
rect 16118 16632 16174 16688
rect 16118 16224 16174 16280
rect 16210 15680 16266 15736
rect 15934 14456 15990 14512
rect 15658 10784 15714 10840
rect 15566 9424 15622 9480
rect 15382 9288 15438 9344
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14738 7928 14794 7984
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 13634 1808 13690 1864
rect 14554 1536 14610 1592
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14830 4936 14886 4992
rect 14738 4392 14794 4448
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15474 8744 15530 8800
rect 15474 7928 15530 7984
rect 15658 9288 15714 9344
rect 15750 6060 15752 6080
rect 15752 6060 15804 6080
rect 15804 6060 15806 6080
rect 15750 6024 15806 6060
rect 16578 15544 16634 15600
rect 16486 14728 16542 14784
rect 16302 9832 16358 9888
rect 16026 9016 16082 9072
rect 15566 3848 15622 3904
rect 15290 3712 15346 3768
rect 15474 3712 15530 3768
rect 14738 3576 14794 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15566 3168 15622 3224
rect 15842 4800 15898 4856
rect 15750 3032 15806 3088
rect 15750 1536 15806 1592
rect 16394 9696 16450 9752
rect 16854 18148 16910 18184
rect 16854 18128 16856 18148
rect 16856 18128 16908 18148
rect 16908 18128 16910 18148
rect 16762 13912 16818 13968
rect 16854 13524 16910 13560
rect 16854 13504 16856 13524
rect 16856 13504 16908 13524
rect 16908 13504 16910 13524
rect 17498 24112 17554 24168
rect 17590 23704 17646 23760
rect 17498 21256 17554 21312
rect 17774 23296 17830 23352
rect 18418 23568 18474 23624
rect 17682 21956 17738 21992
rect 17682 21936 17684 21956
rect 17684 21936 17736 21956
rect 17736 21936 17738 21956
rect 17590 20848 17646 20904
rect 17498 18264 17554 18320
rect 17222 14048 17278 14104
rect 16670 10512 16726 10568
rect 16394 9560 16450 9616
rect 16302 6296 16358 6352
rect 16762 7520 16818 7576
rect 16578 6432 16634 6488
rect 16762 6160 16818 6216
rect 16946 7248 17002 7304
rect 16854 5752 16910 5808
rect 17314 13640 17370 13696
rect 17222 9152 17278 9208
rect 17130 8336 17186 8392
rect 17222 6976 17278 7032
rect 17314 4936 17370 4992
rect 16670 2644 16726 2680
rect 16670 2624 16672 2644
rect 16672 2624 16724 2644
rect 16724 2624 16726 2644
rect 16854 2760 16910 2816
rect 16670 2252 16672 2272
rect 16672 2252 16724 2272
rect 16724 2252 16726 2272
rect 16670 2216 16726 2252
rect 17498 15952 17554 16008
rect 17498 15544 17554 15600
rect 18602 21836 18604 21856
rect 18604 21836 18656 21856
rect 18656 21836 18658 21856
rect 18602 21800 18658 21836
rect 18234 19624 18290 19680
rect 17958 17992 18014 18048
rect 17958 17740 18014 17776
rect 17958 17720 17960 17740
rect 17960 17720 18012 17740
rect 18012 17720 18014 17740
rect 18234 17720 18290 17776
rect 17774 15680 17830 15736
rect 17682 14728 17738 14784
rect 18050 14592 18106 14648
rect 17590 14048 17646 14104
rect 17866 13640 17922 13696
rect 17682 12960 17738 13016
rect 17590 12844 17646 12880
rect 17590 12824 17592 12844
rect 17592 12824 17644 12844
rect 17644 12824 17646 12844
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19246 21664 19302 21720
rect 18786 18400 18842 18456
rect 18510 15544 18566 15600
rect 18510 14764 18512 14784
rect 18512 14764 18564 14784
rect 18564 14764 18566 14784
rect 18510 14728 18566 14764
rect 18234 12552 18290 12608
rect 18142 12164 18198 12200
rect 18142 12144 18144 12164
rect 18144 12144 18196 12164
rect 18196 12144 18198 12164
rect 18050 11872 18106 11928
rect 17774 11756 17830 11792
rect 17774 11736 17776 11756
rect 17776 11736 17828 11756
rect 17828 11736 17830 11756
rect 17590 11328 17646 11384
rect 18050 11348 18106 11384
rect 18050 11328 18052 11348
rect 18052 11328 18104 11348
rect 18104 11328 18106 11348
rect 17958 10376 18014 10432
rect 17498 8916 17500 8936
rect 17500 8916 17552 8936
rect 17552 8916 17554 8936
rect 17498 8880 17554 8916
rect 17590 7404 17646 7440
rect 17590 7384 17592 7404
rect 17592 7384 17644 7404
rect 17644 7384 17646 7404
rect 17498 6860 17554 6896
rect 17498 6840 17500 6860
rect 17500 6840 17552 6860
rect 17552 6840 17554 6860
rect 17682 6724 17738 6760
rect 17682 6704 17684 6724
rect 17684 6704 17736 6724
rect 17736 6704 17738 6724
rect 17682 5072 17738 5128
rect 18418 11056 18474 11112
rect 18326 9968 18382 10024
rect 18326 9696 18382 9752
rect 18142 8200 18198 8256
rect 17958 3712 18014 3768
rect 18050 3440 18106 3496
rect 17406 1808 17462 1864
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19982 23160 20038 23216
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19522 21548 19578 21584
rect 19522 21528 19524 21548
rect 19524 21528 19576 21548
rect 19576 21528 19578 21548
rect 19614 21392 19670 21448
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19522 20984 19578 21040
rect 19706 21004 19762 21040
rect 19706 20984 19708 21004
rect 19708 20984 19760 21004
rect 19760 20984 19762 21004
rect 18970 17484 18972 17504
rect 18972 17484 19024 17504
rect 19024 17484 19026 17504
rect 18970 17448 19026 17484
rect 18878 14864 18934 14920
rect 18970 13776 19026 13832
rect 18970 12552 19026 12608
rect 18878 12316 18880 12336
rect 18880 12316 18932 12336
rect 18932 12316 18934 12336
rect 18878 12280 18934 12316
rect 18694 8336 18750 8392
rect 18878 7948 18934 7984
rect 18878 7928 18880 7948
rect 18880 7928 18932 7948
rect 18932 7928 18934 7948
rect 18786 5344 18842 5400
rect 18694 5072 18750 5128
rect 18510 3440 18566 3496
rect 18142 3052 18198 3088
rect 18142 3032 18144 3052
rect 18144 3032 18196 3052
rect 18196 3032 18198 3052
rect 18878 1672 18934 1728
rect 18694 1400 18750 1456
rect 19246 16940 19248 16960
rect 19248 16940 19300 16960
rect 19300 16940 19302 16960
rect 19246 16904 19302 16940
rect 19246 16360 19302 16416
rect 20074 22344 20130 22400
rect 19982 20304 20038 20360
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 20074 20052 20130 20088
rect 20074 20032 20076 20052
rect 20076 20032 20128 20052
rect 20128 20032 20130 20052
rect 20442 21564 20444 21584
rect 20444 21564 20496 21584
rect 20496 21564 20498 21584
rect 20442 21528 20498 21564
rect 20350 20984 20406 21040
rect 20166 19896 20222 19952
rect 20166 19488 20222 19544
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20258 18672 20314 18728
rect 19982 17196 20038 17232
rect 19982 17176 19984 17196
rect 19984 17176 20036 17196
rect 20036 17176 20038 17196
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19890 16088 19946 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19614 15000 19670 15056
rect 19154 12552 19210 12608
rect 19430 13640 19486 13696
rect 19062 12008 19118 12064
rect 19246 11600 19302 11656
rect 19246 10648 19302 10704
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19706 12860 19708 12880
rect 19708 12860 19760 12880
rect 19760 12860 19762 12880
rect 19706 12824 19762 12860
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19890 12180 19892 12200
rect 19892 12180 19944 12200
rect 19944 12180 19946 12200
rect 19890 12144 19946 12180
rect 20074 14068 20130 14104
rect 20074 14048 20076 14068
rect 20076 14048 20128 14068
rect 20128 14048 20130 14068
rect 20166 12552 20222 12608
rect 20074 11464 20130 11520
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 23386 26560 23442 26616
rect 23294 26016 23350 26072
rect 20902 23724 20958 23760
rect 20902 23704 20904 23724
rect 20904 23704 20956 23724
rect 20956 23704 20958 23724
rect 20994 22888 21050 22944
rect 20994 22072 21050 22128
rect 20810 21800 20866 21856
rect 20994 21664 21050 21720
rect 22466 23296 22522 23352
rect 22190 22888 22246 22944
rect 21454 22616 21510 22672
rect 21362 21800 21418 21856
rect 21086 20304 21142 20360
rect 20718 19352 20774 19408
rect 20810 17448 20866 17504
rect 20442 13504 20498 13560
rect 21270 18944 21326 19000
rect 21914 21392 21970 21448
rect 22006 21120 22062 21176
rect 22006 20596 22062 20632
rect 22006 20576 22008 20596
rect 22008 20576 22060 20596
rect 22060 20576 22062 20596
rect 21546 20304 21602 20360
rect 21178 18264 21234 18320
rect 21270 17740 21326 17776
rect 21270 17720 21272 17740
rect 21272 17720 21324 17740
rect 21324 17720 21326 17740
rect 21822 18284 21878 18320
rect 21822 18264 21824 18284
rect 21824 18264 21876 18284
rect 21876 18264 21878 18284
rect 22098 19660 22100 19680
rect 22100 19660 22152 19680
rect 22152 19660 22154 19680
rect 22098 19624 22154 19660
rect 22006 19216 22062 19272
rect 22834 22516 22836 22536
rect 22836 22516 22888 22536
rect 22888 22516 22890 22536
rect 22834 22480 22890 22516
rect 21454 17060 21510 17096
rect 21454 17040 21456 17060
rect 21456 17040 21508 17060
rect 21508 17040 21510 17060
rect 21178 16360 21234 16416
rect 21178 15952 21234 16008
rect 22650 18672 22706 18728
rect 22558 17856 22614 17912
rect 22466 17312 22522 17368
rect 22374 17040 22430 17096
rect 22282 15988 22284 16008
rect 22284 15988 22336 16008
rect 22336 15988 22338 16008
rect 22282 15952 22338 15988
rect 21730 15408 21786 15464
rect 21178 13912 21234 13968
rect 20442 12960 20498 13016
rect 19890 10648 19946 10704
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 20350 10140 20352 10160
rect 20352 10140 20404 10160
rect 20404 10140 20406 10160
rect 20350 10104 20406 10140
rect 19890 9560 19946 9616
rect 19430 8880 19486 8936
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19154 7928 19210 7984
rect 19614 7792 19670 7848
rect 19798 7828 19800 7848
rect 19800 7828 19852 7848
rect 19852 7828 19854 7848
rect 19798 7792 19854 7828
rect 20074 8200 20130 8256
rect 19522 7248 19578 7304
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19246 6160 19302 6216
rect 20074 6432 20130 6488
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19522 5616 19578 5672
rect 19338 2760 19394 2816
rect 18970 856 19026 912
rect 20074 5752 20130 5808
rect 20902 12688 20958 12744
rect 20718 12552 20774 12608
rect 20902 11620 20958 11656
rect 20902 11600 20904 11620
rect 20904 11600 20956 11620
rect 20956 11600 20958 11620
rect 21086 12436 21142 12472
rect 21086 12416 21088 12436
rect 21088 12416 21140 12436
rect 21140 12416 21142 12436
rect 20810 9968 20866 10024
rect 20626 8372 20628 8392
rect 20628 8372 20680 8392
rect 20680 8372 20682 8392
rect 20626 8336 20682 8372
rect 21546 12724 21548 12744
rect 21548 12724 21600 12744
rect 21600 12724 21602 12744
rect 21546 12688 21602 12724
rect 21362 11736 21418 11792
rect 21822 14864 21878 14920
rect 22190 14456 22246 14512
rect 22006 13776 22062 13832
rect 21822 10920 21878 10976
rect 21270 10512 21326 10568
rect 21178 9696 21234 9752
rect 22558 16904 22614 16960
rect 22466 15020 22522 15056
rect 22466 15000 22468 15020
rect 22468 15000 22520 15020
rect 22520 15000 22522 15020
rect 22650 16652 22706 16688
rect 22650 16632 22652 16652
rect 22652 16632 22704 16652
rect 22704 16632 22706 16652
rect 22466 12416 22522 12472
rect 22190 12144 22246 12200
rect 21086 8064 21142 8120
rect 21270 7656 21326 7712
rect 21086 7384 21142 7440
rect 22742 10684 22744 10704
rect 22744 10684 22796 10704
rect 22796 10684 22798 10704
rect 22742 10648 22798 10684
rect 22282 8472 22338 8528
rect 22282 8336 22338 8392
rect 22190 8064 22246 8120
rect 20718 6160 20774 6216
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19706 4528 19762 4584
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19614 3596 19670 3632
rect 19614 3576 19616 3596
rect 19616 3576 19668 3596
rect 19668 3576 19670 3596
rect 21086 5208 21142 5264
rect 21086 4664 21142 4720
rect 22466 5772 22522 5808
rect 22466 5752 22468 5772
rect 22468 5752 22520 5772
rect 22520 5752 22522 5772
rect 21822 4004 21878 4040
rect 21822 3984 21824 4004
rect 21824 3984 21876 4004
rect 21876 3984 21878 4004
rect 22006 3984 22062 4040
rect 22650 4120 22706 4176
rect 20442 3440 20498 3496
rect 20350 2896 20406 2952
rect 20074 2760 20130 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 21546 3032 21602 3088
rect 21914 3032 21970 3088
rect 20902 2508 20958 2544
rect 20902 2488 20904 2508
rect 20904 2488 20956 2508
rect 20956 2488 20958 2508
rect 22558 3712 22614 3768
rect 22098 2352 22154 2408
rect 20718 1944 20774 2000
rect 21362 1536 21418 1592
rect 22926 13368 22982 13424
rect 23662 25336 23718 25392
rect 24766 27104 24822 27160
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24792 24822 24848
rect 23754 24248 23810 24304
rect 23478 23704 23534 23760
rect 23754 23024 23810 23080
rect 23754 22888 23810 22944
rect 23294 22752 23350 22808
rect 23662 20340 23664 20360
rect 23664 20340 23716 20360
rect 23716 20340 23718 20360
rect 23662 20304 23718 20340
rect 23662 19488 23718 19544
rect 23478 19352 23534 19408
rect 23570 17584 23626 17640
rect 23110 12300 23166 12336
rect 23110 12280 23112 12300
rect 23112 12280 23164 12300
rect 23164 12280 23166 12300
rect 23018 10920 23074 10976
rect 23018 8744 23074 8800
rect 23478 16768 23534 16824
rect 23662 16224 23718 16280
rect 24030 22616 24086 22672
rect 23846 21936 23902 21992
rect 24030 21140 24086 21176
rect 24030 21120 24032 21140
rect 24032 21120 24084 21140
rect 24084 21120 24086 21140
rect 24030 20576 24086 20632
rect 25502 24656 25558 24712
rect 24582 24112 24638 24168
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25870 24248 25926 24304
rect 24766 23160 24822 23216
rect 25226 23296 25282 23352
rect 24398 22380 24400 22400
rect 24400 22380 24452 22400
rect 24452 22380 24454 22400
rect 24398 22344 24454 22380
rect 24766 22092 24822 22128
rect 24766 22072 24768 22092
rect 24768 22072 24820 22092
rect 24820 22072 24822 22092
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24214 21392 24270 21448
rect 24490 20984 24546 21040
rect 24674 20984 24730 21040
rect 24122 20440 24178 20496
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24674 20304 24730 20360
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24122 18808 24178 18864
rect 24122 18420 24178 18456
rect 24122 18400 24124 18420
rect 24124 18400 24176 18420
rect 24176 18400 24178 18420
rect 23938 16496 23994 16552
rect 23846 14592 23902 14648
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24766 19080 24822 19136
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 16904 24822 16960
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24122 15680 24178 15736
rect 23846 13096 23902 13152
rect 23478 9560 23534 9616
rect 23294 8200 23350 8256
rect 23478 8064 23534 8120
rect 23110 5616 23166 5672
rect 23018 5344 23074 5400
rect 23018 4800 23074 4856
rect 23478 2760 23534 2816
rect 23754 12416 23810 12472
rect 24122 13504 24178 13560
rect 24122 13368 24178 13424
rect 23938 12824 23994 12880
rect 23846 11872 23902 11928
rect 23846 8880 23902 8936
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24766 15136 24822 15192
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 25042 22072 25098 22128
rect 25502 23024 25558 23080
rect 25134 21564 25136 21584
rect 25136 21564 25188 21584
rect 25188 21564 25190 21584
rect 25134 21528 25190 21564
rect 25042 21120 25098 21176
rect 25410 20460 25466 20496
rect 25410 20440 25412 20460
rect 25412 20440 25464 20460
rect 25464 20440 25466 20460
rect 25226 20168 25282 20224
rect 25226 19252 25228 19272
rect 25228 19252 25280 19272
rect 25280 19252 25282 19272
rect 25226 19216 25282 19252
rect 25686 19624 25742 19680
rect 25042 17856 25098 17912
rect 25226 18164 25228 18184
rect 25228 18164 25280 18184
rect 25280 18164 25282 18184
rect 25226 18128 25282 18164
rect 25502 18944 25558 19000
rect 25594 18808 25650 18864
rect 25410 18028 25412 18048
rect 25412 18028 25464 18048
rect 25464 18028 25466 18048
rect 25410 17992 25466 18028
rect 25318 17484 25320 17504
rect 25320 17484 25372 17504
rect 25372 17484 25374 17504
rect 25318 17448 25374 17484
rect 25318 17212 25320 17232
rect 25320 17212 25372 17232
rect 25372 17212 25374 17232
rect 25318 17176 25374 17212
rect 25410 17040 25466 17096
rect 25042 13812 25044 13832
rect 25044 13812 25096 13832
rect 25096 13812 25098 13832
rect 25042 13776 25098 13812
rect 24582 12144 24638 12200
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24122 11464 24178 11520
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24122 10512 24178 10568
rect 23846 8472 23902 8528
rect 23846 6704 23902 6760
rect 23754 6296 23810 6352
rect 24122 9832 24178 9888
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24214 8200 24270 8256
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24122 4428 24124 4448
rect 24124 4428 24176 4448
rect 24176 4428 24178 4448
rect 24122 4392 24178 4428
rect 24122 4120 24178 4176
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24766 12280 24822 12336
rect 24766 9424 24822 9480
rect 25318 13232 25374 13288
rect 24766 7928 24822 7984
rect 24766 7384 24822 7440
rect 24766 6568 24822 6624
rect 24766 5244 24768 5264
rect 24768 5244 24820 5264
rect 24820 5244 24822 5264
rect 24766 5208 24822 5244
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24858 4800 24914 4856
rect 24582 2896 24638 2952
rect 24582 2488 24638 2544
rect 26882 23568 26938 23624
rect 27526 20032 27582 20088
rect 25318 4800 25374 4856
rect 25318 3984 25374 4040
rect 23754 1400 23810 1456
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 26054 4256 26110 4312
rect 23662 312 23718 368
<< metal3 >>
rect 23749 27706 23815 27709
rect 27520 27706 28000 27736
rect 23749 27704 28000 27706
rect 23749 27648 23754 27704
rect 23810 27648 28000 27704
rect 23749 27646 28000 27648
rect 23749 27643 23815 27646
rect 27520 27616 28000 27646
rect 24761 27162 24827 27165
rect 27520 27162 28000 27192
rect 24761 27160 28000 27162
rect 24761 27104 24766 27160
rect 24822 27104 28000 27160
rect 24761 27102 28000 27104
rect 24761 27099 24827 27102
rect 27520 27072 28000 27102
rect 23381 26618 23447 26621
rect 27520 26618 28000 26648
rect 23381 26616 28000 26618
rect 23381 26560 23386 26616
rect 23442 26560 28000 26616
rect 23381 26558 28000 26560
rect 23381 26555 23447 26558
rect 27520 26528 28000 26558
rect 23289 26074 23355 26077
rect 27520 26074 28000 26104
rect 23289 26072 28000 26074
rect 23289 26016 23294 26072
rect 23350 26016 28000 26072
rect 23289 26014 28000 26016
rect 23289 26011 23355 26014
rect 27520 25984 28000 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 23657 25394 23723 25397
rect 27520 25394 28000 25424
rect 23657 25392 28000 25394
rect 23657 25336 23662 25392
rect 23718 25336 28000 25392
rect 23657 25334 28000 25336
rect 23657 25331 23723 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 5993 24850 6059 24853
rect 12801 24850 12867 24853
rect 14549 24850 14615 24853
rect 5993 24848 12634 24850
rect 5993 24792 5998 24848
rect 6054 24792 12634 24848
rect 5993 24790 12634 24792
rect 5993 24787 6059 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 933 24442 999 24445
rect 5993 24442 6059 24445
rect 933 24440 6059 24442
rect 933 24384 938 24440
rect 994 24384 5998 24440
rect 6054 24384 6059 24440
rect 933 24382 6059 24384
rect 933 24379 999 24382
rect 5993 24379 6059 24382
rect 12574 24306 12634 24790
rect 12801 24848 14615 24850
rect 12801 24792 12806 24848
rect 12862 24792 14554 24848
rect 14610 24792 14615 24848
rect 12801 24790 14615 24792
rect 12801 24787 12867 24790
rect 14549 24787 14615 24790
rect 24761 24850 24827 24853
rect 27520 24850 28000 24880
rect 24761 24848 28000 24850
rect 24761 24792 24766 24848
rect 24822 24792 28000 24848
rect 24761 24790 28000 24792
rect 24761 24787 24827 24790
rect 27520 24760 28000 24790
rect 13721 24714 13787 24717
rect 25497 24714 25563 24717
rect 13721 24712 25563 24714
rect 13721 24656 13726 24712
rect 13782 24656 25502 24712
rect 25558 24656 25563 24712
rect 13721 24654 25563 24656
rect 13721 24651 13787 24654
rect 25497 24651 25563 24654
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 13905 24442 13971 24445
rect 16205 24442 16271 24445
rect 13905 24440 16271 24442
rect 13905 24384 13910 24440
rect 13966 24384 16210 24440
rect 16266 24384 16271 24440
rect 13905 24382 16271 24384
rect 13905 24379 13971 24382
rect 16205 24379 16271 24382
rect 14273 24306 14339 24309
rect 12574 24304 14339 24306
rect 12574 24248 14278 24304
rect 14334 24248 14339 24304
rect 12574 24246 14339 24248
rect 14273 24243 14339 24246
rect 14917 24306 14983 24309
rect 23749 24306 23815 24309
rect 14917 24304 23815 24306
rect 14917 24248 14922 24304
rect 14978 24248 23754 24304
rect 23810 24248 23815 24304
rect 14917 24246 23815 24248
rect 14917 24243 14983 24246
rect 23749 24243 23815 24246
rect 25865 24306 25931 24309
rect 27520 24306 28000 24336
rect 25865 24304 28000 24306
rect 25865 24248 25870 24304
rect 25926 24248 28000 24304
rect 25865 24246 28000 24248
rect 25865 24243 25931 24246
rect 27520 24216 28000 24246
rect 9121 24170 9187 24173
rect 15929 24170 15995 24173
rect 9121 24168 15995 24170
rect 9121 24112 9126 24168
rect 9182 24112 15934 24168
rect 15990 24112 15995 24168
rect 9121 24110 15995 24112
rect 9121 24107 9187 24110
rect 15929 24107 15995 24110
rect 17493 24170 17559 24173
rect 24577 24170 24643 24173
rect 17493 24168 24643 24170
rect 17493 24112 17498 24168
rect 17554 24112 24582 24168
rect 24638 24112 24643 24168
rect 17493 24110 24643 24112
rect 17493 24107 17559 24110
rect 24577 24107 24643 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 7741 23898 7807 23901
rect 12065 23898 12131 23901
rect 7741 23896 12131 23898
rect 7741 23840 7746 23896
rect 7802 23840 12070 23896
rect 12126 23840 12131 23896
rect 7741 23838 12131 23840
rect 7741 23835 7807 23838
rect 12065 23835 12131 23838
rect 12525 23898 12591 23901
rect 14733 23898 14799 23901
rect 12525 23896 14799 23898
rect 12525 23840 12530 23896
rect 12586 23840 14738 23896
rect 14794 23840 14799 23896
rect 12525 23838 14799 23840
rect 12525 23835 12591 23838
rect 14733 23835 14799 23838
rect 3693 23762 3759 23765
rect 6085 23762 6151 23765
rect 3693 23760 6151 23762
rect 3693 23704 3698 23760
rect 3754 23704 6090 23760
rect 6146 23704 6151 23760
rect 3693 23702 6151 23704
rect 3693 23699 3759 23702
rect 6085 23699 6151 23702
rect 17585 23762 17651 23765
rect 20897 23762 20963 23765
rect 17585 23760 20963 23762
rect 17585 23704 17590 23760
rect 17646 23704 20902 23760
rect 20958 23704 20963 23760
rect 17585 23702 20963 23704
rect 17585 23699 17651 23702
rect 20897 23699 20963 23702
rect 23473 23762 23539 23765
rect 27520 23762 28000 23792
rect 23473 23760 28000 23762
rect 23473 23704 23478 23760
rect 23534 23704 28000 23760
rect 23473 23702 28000 23704
rect 23473 23699 23539 23702
rect 27520 23672 28000 23702
rect 11605 23626 11671 23629
rect 13169 23626 13235 23629
rect 11605 23624 13235 23626
rect 11605 23568 11610 23624
rect 11666 23568 13174 23624
rect 13230 23568 13235 23624
rect 11605 23566 13235 23568
rect 11605 23563 11671 23566
rect 13169 23563 13235 23566
rect 18413 23626 18479 23629
rect 26877 23626 26943 23629
rect 18413 23624 26943 23626
rect 18413 23568 18418 23624
rect 18474 23568 26882 23624
rect 26938 23568 26943 23624
rect 18413 23566 26943 23568
rect 18413 23563 18479 23566
rect 26877 23563 26943 23566
rect 7097 23490 7163 23493
rect 10133 23490 10199 23493
rect 7097 23488 10199 23490
rect 7097 23432 7102 23488
rect 7158 23432 10138 23488
rect 10194 23432 10199 23488
rect 7097 23430 10199 23432
rect 7097 23427 7163 23430
rect 10133 23427 10199 23430
rect 11145 23490 11211 23493
rect 12433 23490 12499 23493
rect 11145 23488 12499 23490
rect 11145 23432 11150 23488
rect 11206 23432 12438 23488
rect 12494 23432 12499 23488
rect 11145 23430 12499 23432
rect 11145 23427 11211 23430
rect 12433 23427 12499 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 11145 23354 11211 23357
rect 17769 23354 17835 23357
rect 11145 23352 17835 23354
rect 11145 23296 11150 23352
rect 11206 23296 17774 23352
rect 17830 23296 17835 23352
rect 11145 23294 17835 23296
rect 11145 23291 11211 23294
rect 17769 23291 17835 23294
rect 22461 23354 22527 23357
rect 25221 23354 25287 23357
rect 22461 23352 25287 23354
rect 22461 23296 22466 23352
rect 22522 23296 25226 23352
rect 25282 23296 25287 23352
rect 22461 23294 25287 23296
rect 22461 23291 22527 23294
rect 25221 23291 25287 23294
rect 6361 23218 6427 23221
rect 12341 23218 12407 23221
rect 19977 23218 20043 23221
rect 6361 23216 12407 23218
rect 6361 23160 6366 23216
rect 6422 23160 12346 23216
rect 12402 23160 12407 23216
rect 6361 23158 12407 23160
rect 6361 23155 6427 23158
rect 12341 23155 12407 23158
rect 14598 23216 20043 23218
rect 14598 23160 19982 23216
rect 20038 23160 20043 23216
rect 14598 23158 20043 23160
rect 10685 23082 10751 23085
rect 14598 23082 14658 23158
rect 19977 23155 20043 23158
rect 24761 23218 24827 23221
rect 27520 23218 28000 23248
rect 24761 23216 28000 23218
rect 24761 23160 24766 23216
rect 24822 23160 28000 23216
rect 24761 23158 28000 23160
rect 24761 23155 24827 23158
rect 27520 23128 28000 23158
rect 10685 23080 14658 23082
rect 10685 23024 10690 23080
rect 10746 23024 14658 23080
rect 10685 23022 14658 23024
rect 23749 23082 23815 23085
rect 25497 23082 25563 23085
rect 23749 23080 25563 23082
rect 23749 23024 23754 23080
rect 23810 23024 25502 23080
rect 25558 23024 25563 23080
rect 23749 23022 25563 23024
rect 10685 23019 10751 23022
rect 23749 23019 23815 23022
rect 25497 23019 25563 23022
rect 20989 22946 21055 22949
rect 22185 22946 22251 22949
rect 23749 22946 23815 22949
rect 20989 22944 23815 22946
rect 20989 22888 20994 22944
rect 21050 22888 22190 22944
rect 22246 22888 23754 22944
rect 23810 22888 23815 22944
rect 20989 22886 23815 22888
rect 20989 22883 21055 22886
rect 22185 22883 22251 22886
rect 23749 22883 23815 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 23289 22810 23355 22813
rect 15702 22808 23355 22810
rect 15702 22752 23294 22808
rect 23350 22752 23355 22808
rect 15702 22750 23355 22752
rect 4981 22674 5047 22677
rect 14222 22674 14228 22676
rect 4981 22672 14228 22674
rect 4981 22616 4986 22672
rect 5042 22616 14228 22672
rect 4981 22614 14228 22616
rect 4981 22611 5047 22614
rect 14222 22612 14228 22614
rect 14292 22674 14298 22676
rect 15285 22674 15351 22677
rect 14292 22672 15351 22674
rect 14292 22616 15290 22672
rect 15346 22616 15351 22672
rect 14292 22614 15351 22616
rect 14292 22612 14298 22614
rect 15285 22611 15351 22614
rect 5993 22538 6059 22541
rect 14549 22538 14615 22541
rect 5993 22536 14615 22538
rect 5993 22480 5998 22536
rect 6054 22480 14554 22536
rect 14610 22480 14615 22536
rect 5993 22478 14615 22480
rect 5993 22475 6059 22478
rect 14549 22475 14615 22478
rect 14733 22538 14799 22541
rect 15702 22538 15762 22750
rect 23289 22747 23355 22750
rect 21449 22674 21515 22677
rect 24025 22674 24091 22677
rect 21449 22672 24091 22674
rect 21449 22616 21454 22672
rect 21510 22616 24030 22672
rect 24086 22616 24091 22672
rect 21449 22614 24091 22616
rect 21449 22611 21515 22614
rect 24025 22611 24091 22614
rect 14733 22536 15762 22538
rect 14733 22480 14738 22536
rect 14794 22480 15762 22536
rect 14733 22478 15762 22480
rect 15929 22538 15995 22541
rect 22829 22538 22895 22541
rect 27520 22538 28000 22568
rect 15929 22536 22895 22538
rect 15929 22480 15934 22536
rect 15990 22480 22834 22536
rect 22890 22480 22895 22536
rect 15929 22478 22895 22480
rect 14733 22475 14799 22478
rect 15929 22475 15995 22478
rect 22829 22475 22895 22478
rect 23844 22478 28000 22538
rect 20069 22402 20135 22405
rect 23844 22402 23904 22478
rect 27520 22448 28000 22478
rect 20069 22400 23904 22402
rect 20069 22344 20074 22400
rect 20130 22344 23904 22400
rect 20069 22342 23904 22344
rect 20069 22339 20135 22342
rect 23974 22340 23980 22404
rect 24044 22402 24050 22404
rect 24393 22402 24459 22405
rect 24044 22400 24459 22402
rect 24044 22344 24398 22400
rect 24454 22344 24459 22400
rect 24044 22342 24459 22344
rect 24044 22340 24050 22342
rect 24393 22339 24459 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 11973 22130 12039 22133
rect 14641 22130 14707 22133
rect 11973 22128 14707 22130
rect 11973 22072 11978 22128
rect 12034 22072 14646 22128
rect 14702 22072 14707 22128
rect 11973 22070 14707 22072
rect 11973 22067 12039 22070
rect 14641 22067 14707 22070
rect 14825 22130 14891 22133
rect 20989 22130 21055 22133
rect 14825 22128 21055 22130
rect 14825 22072 14830 22128
rect 14886 22072 20994 22128
rect 21050 22072 21055 22128
rect 14825 22070 21055 22072
rect 14825 22067 14891 22070
rect 20989 22067 21055 22070
rect 24761 22130 24827 22133
rect 25037 22130 25103 22133
rect 24761 22128 25103 22130
rect 24761 22072 24766 22128
rect 24822 22072 25042 22128
rect 25098 22072 25103 22128
rect 24761 22070 25103 22072
rect 24761 22067 24827 22070
rect 25037 22067 25103 22070
rect 2957 21994 3023 21997
rect 15561 21994 15627 21997
rect 2957 21992 15627 21994
rect 2957 21936 2962 21992
rect 3018 21936 15566 21992
rect 15622 21936 15627 21992
rect 2957 21934 15627 21936
rect 2957 21931 3023 21934
rect 15561 21931 15627 21934
rect 17677 21994 17743 21997
rect 23841 21994 23907 21997
rect 27520 21994 28000 22024
rect 17677 21992 23907 21994
rect 17677 21936 17682 21992
rect 17738 21936 23846 21992
rect 23902 21936 23907 21992
rect 17677 21934 23907 21936
rect 17677 21931 17743 21934
rect 23841 21931 23907 21934
rect 23982 21934 28000 21994
rect 18597 21858 18663 21861
rect 20805 21858 20871 21861
rect 18597 21856 20871 21858
rect 18597 21800 18602 21856
rect 18658 21800 20810 21856
rect 20866 21800 20871 21856
rect 18597 21798 20871 21800
rect 18597 21795 18663 21798
rect 20805 21795 20871 21798
rect 21357 21858 21423 21861
rect 23982 21858 24042 21934
rect 27520 21904 28000 21934
rect 21357 21856 24042 21858
rect 21357 21800 21362 21856
rect 21418 21800 24042 21856
rect 21357 21798 24042 21800
rect 21357 21795 21423 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 9765 21722 9831 21725
rect 19241 21722 19307 21725
rect 20989 21722 21055 21725
rect 9765 21720 14842 21722
rect 9765 21664 9770 21720
rect 9826 21664 14842 21720
rect 9765 21662 14842 21664
rect 9765 21659 9831 21662
rect 6085 21586 6151 21589
rect 14365 21586 14431 21589
rect 6085 21584 14431 21586
rect 6085 21528 6090 21584
rect 6146 21528 14370 21584
rect 14426 21528 14431 21584
rect 6085 21526 14431 21528
rect 14782 21586 14842 21662
rect 19241 21720 21055 21722
rect 19241 21664 19246 21720
rect 19302 21664 20994 21720
rect 21050 21664 21055 21720
rect 19241 21662 21055 21664
rect 19241 21659 19307 21662
rect 20989 21659 21055 21662
rect 15469 21586 15535 21589
rect 19517 21586 19583 21589
rect 14782 21584 19583 21586
rect 14782 21528 15474 21584
rect 15530 21528 19522 21584
rect 19578 21528 19583 21584
rect 14782 21526 19583 21528
rect 6085 21523 6151 21526
rect 14365 21523 14431 21526
rect 15469 21523 15535 21526
rect 19517 21523 19583 21526
rect 20437 21586 20503 21589
rect 25129 21586 25195 21589
rect 20437 21584 25195 21586
rect 20437 21528 20442 21584
rect 20498 21528 25134 21584
rect 25190 21528 25195 21584
rect 20437 21526 25195 21528
rect 20437 21523 20503 21526
rect 25129 21523 25195 21526
rect 10225 21450 10291 21453
rect 13169 21450 13235 21453
rect 10225 21448 13235 21450
rect 10225 21392 10230 21448
rect 10286 21392 13174 21448
rect 13230 21392 13235 21448
rect 10225 21390 13235 21392
rect 10225 21387 10291 21390
rect 13169 21387 13235 21390
rect 19609 21450 19675 21453
rect 21909 21450 21975 21453
rect 19609 21448 21975 21450
rect 19609 21392 19614 21448
rect 19670 21392 21914 21448
rect 21970 21392 21975 21448
rect 19609 21390 21975 21392
rect 19609 21387 19675 21390
rect 21909 21387 21975 21390
rect 24209 21450 24275 21453
rect 27520 21450 28000 21480
rect 24209 21448 28000 21450
rect 24209 21392 24214 21448
rect 24270 21392 28000 21448
rect 24209 21390 28000 21392
rect 24209 21387 24275 21390
rect 27520 21360 28000 21390
rect 11605 21314 11671 21317
rect 17493 21314 17559 21317
rect 11605 21312 17559 21314
rect 11605 21256 11610 21312
rect 11666 21256 17498 21312
rect 17554 21256 17559 21312
rect 11605 21254 17559 21256
rect 11605 21251 11671 21254
rect 17493 21251 17559 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 22001 21178 22067 21181
rect 24025 21178 24091 21181
rect 25037 21178 25103 21181
rect 22001 21176 25103 21178
rect 22001 21120 22006 21176
rect 22062 21120 24030 21176
rect 24086 21120 25042 21176
rect 25098 21120 25103 21176
rect 22001 21118 25103 21120
rect 22001 21115 22067 21118
rect 24025 21115 24091 21118
rect 25037 21115 25103 21118
rect 0 21042 480 21072
rect 4061 21042 4127 21045
rect 0 21040 4127 21042
rect 0 20984 4066 21040
rect 4122 20984 4127 21040
rect 0 20982 4127 20984
rect 0 20952 480 20982
rect 4061 20979 4127 20982
rect 13445 21042 13511 21045
rect 19517 21042 19583 21045
rect 13445 21040 19583 21042
rect 13445 20984 13450 21040
rect 13506 20984 19522 21040
rect 19578 20984 19583 21040
rect 13445 20982 19583 20984
rect 13445 20979 13511 20982
rect 19517 20979 19583 20982
rect 19701 21042 19767 21045
rect 20345 21042 20411 21045
rect 24485 21042 24551 21045
rect 19701 21040 24551 21042
rect 19701 20984 19706 21040
rect 19762 20984 20350 21040
rect 20406 20984 24490 21040
rect 24546 20984 24551 21040
rect 19701 20982 24551 20984
rect 19701 20979 19767 20982
rect 20345 20979 20411 20982
rect 24485 20979 24551 20982
rect 24669 21042 24735 21045
rect 24669 21040 24778 21042
rect 24669 20984 24674 21040
rect 24730 20984 24778 21040
rect 24669 20979 24778 20984
rect 13997 20906 14063 20909
rect 17585 20906 17651 20909
rect 13997 20904 17651 20906
rect 13997 20848 14002 20904
rect 14058 20848 17590 20904
rect 17646 20848 17651 20904
rect 13997 20846 17651 20848
rect 24718 20906 24778 20979
rect 27520 20906 28000 20936
rect 24718 20846 28000 20906
rect 13997 20843 14063 20846
rect 17585 20843 17651 20846
rect 27520 20816 28000 20846
rect 9397 20770 9463 20773
rect 12433 20770 12499 20773
rect 9397 20768 12499 20770
rect 9397 20712 9402 20768
rect 9458 20712 12438 20768
rect 12494 20712 12499 20768
rect 9397 20710 12499 20712
rect 9397 20707 9463 20710
rect 12433 20707 12499 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 22001 20634 22067 20637
rect 24025 20634 24091 20637
rect 22001 20632 24091 20634
rect 22001 20576 22006 20632
rect 22062 20576 24030 20632
rect 24086 20576 24091 20632
rect 22001 20574 24091 20576
rect 22001 20571 22067 20574
rect 24025 20571 24091 20574
rect 9765 20498 9831 20501
rect 24117 20498 24183 20501
rect 25405 20498 25471 20501
rect 9765 20496 24042 20498
rect 9765 20440 9770 20496
rect 9826 20440 24042 20496
rect 9765 20438 24042 20440
rect 9765 20435 9831 20438
rect 19977 20362 20043 20365
rect 21081 20362 21147 20365
rect 19977 20360 21147 20362
rect 19977 20304 19982 20360
rect 20038 20304 21086 20360
rect 21142 20304 21147 20360
rect 19977 20302 21147 20304
rect 19977 20299 20043 20302
rect 21081 20299 21147 20302
rect 21541 20362 21607 20365
rect 23657 20362 23723 20365
rect 21541 20360 23723 20362
rect 21541 20304 21546 20360
rect 21602 20304 23662 20360
rect 23718 20304 23723 20360
rect 21541 20302 23723 20304
rect 21541 20299 21607 20302
rect 23657 20299 23723 20302
rect 23982 20226 24042 20438
rect 24117 20496 25471 20498
rect 24117 20440 24122 20496
rect 24178 20440 25410 20496
rect 25466 20440 25471 20496
rect 24117 20438 25471 20440
rect 24117 20435 24183 20438
rect 25405 20435 25471 20438
rect 24669 20362 24735 20365
rect 27520 20362 28000 20392
rect 24669 20360 28000 20362
rect 24669 20304 24674 20360
rect 24730 20304 28000 20360
rect 24669 20302 28000 20304
rect 24669 20299 24735 20302
rect 27520 20272 28000 20302
rect 25221 20226 25287 20229
rect 23982 20224 25287 20226
rect 23982 20168 25226 20224
rect 25282 20168 25287 20224
rect 23982 20166 25287 20168
rect 25221 20163 25287 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 12341 20090 12407 20093
rect 13905 20090 13971 20093
rect 12341 20088 13971 20090
rect 12341 20032 12346 20088
rect 12402 20032 13910 20088
rect 13966 20032 13971 20088
rect 12341 20030 13971 20032
rect 12341 20027 12407 20030
rect 13905 20027 13971 20030
rect 20069 20090 20135 20093
rect 27521 20090 27587 20093
rect 20069 20088 27587 20090
rect 20069 20032 20074 20088
rect 20130 20032 27526 20088
rect 27582 20032 27587 20088
rect 20069 20030 27587 20032
rect 20069 20027 20135 20030
rect 27521 20027 27587 20030
rect 13813 19954 13879 19957
rect 20161 19954 20227 19957
rect 13813 19952 20227 19954
rect 13813 19896 13818 19952
rect 13874 19896 20166 19952
rect 20222 19896 20227 19952
rect 13813 19894 20227 19896
rect 13813 19891 13879 19894
rect 20161 19891 20227 19894
rect 9765 19818 9831 19821
rect 15929 19818 15995 19821
rect 9765 19816 15995 19818
rect 9765 19760 9770 19816
rect 9826 19760 15934 19816
rect 15990 19760 15995 19816
rect 9765 19758 15995 19760
rect 9765 19755 9831 19758
rect 15929 19755 15995 19758
rect 18229 19682 18295 19685
rect 22093 19682 22159 19685
rect 18229 19680 22159 19682
rect 18229 19624 18234 19680
rect 18290 19624 22098 19680
rect 22154 19624 22159 19680
rect 18229 19622 22159 19624
rect 18229 19619 18295 19622
rect 22093 19619 22159 19622
rect 25681 19682 25747 19685
rect 27520 19682 28000 19712
rect 25681 19680 28000 19682
rect 25681 19624 25686 19680
rect 25742 19624 28000 19680
rect 25681 19622 28000 19624
rect 25681 19619 25747 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19622
rect 24277 19551 24597 19552
rect 16113 19546 16179 19549
rect 20161 19546 20227 19549
rect 23657 19546 23723 19549
rect 16113 19544 16866 19546
rect 16113 19488 16118 19544
rect 16174 19488 16866 19544
rect 16113 19486 16866 19488
rect 16113 19483 16179 19486
rect 11237 19410 11303 19413
rect 13813 19410 13879 19413
rect 11237 19408 13879 19410
rect 11237 19352 11242 19408
rect 11298 19352 13818 19408
rect 13874 19352 13879 19408
rect 11237 19350 13879 19352
rect 11237 19347 11303 19350
rect 13813 19347 13879 19350
rect 14089 19376 14155 19379
rect 14222 19376 14228 19412
rect 14089 19374 14228 19376
rect 14089 19318 14094 19374
rect 14150 19348 14228 19374
rect 14292 19348 14298 19412
rect 16665 19410 16731 19413
rect 16806 19410 16866 19486
rect 20161 19544 23723 19546
rect 20161 19488 20166 19544
rect 20222 19488 23662 19544
rect 23718 19488 23723 19544
rect 20161 19486 23723 19488
rect 20161 19483 20227 19486
rect 23657 19483 23723 19486
rect 16665 19408 16866 19410
rect 16665 19352 16670 19408
rect 16726 19352 16866 19408
rect 16665 19350 16866 19352
rect 20713 19410 20779 19413
rect 23473 19410 23539 19413
rect 20713 19408 23539 19410
rect 20713 19352 20718 19408
rect 20774 19352 23478 19408
rect 23534 19352 23539 19408
rect 20713 19350 23539 19352
rect 14150 19318 14290 19348
rect 16665 19347 16731 19350
rect 20713 19347 20779 19350
rect 23473 19347 23539 19350
rect 14089 19316 14290 19318
rect 14089 19313 14155 19316
rect 10225 19274 10291 19277
rect 13813 19274 13879 19277
rect 10225 19272 13879 19274
rect 10225 19216 10230 19272
rect 10286 19216 13818 19272
rect 13874 19216 13879 19272
rect 10225 19214 13879 19216
rect 10225 19211 10291 19214
rect 13813 19211 13879 19214
rect 22001 19274 22067 19277
rect 25221 19274 25287 19277
rect 22001 19272 25287 19274
rect 22001 19216 22006 19272
rect 22062 19216 25226 19272
rect 25282 19216 25287 19272
rect 22001 19214 25287 19216
rect 22001 19211 22067 19214
rect 25221 19211 25287 19214
rect 24761 19138 24827 19141
rect 27520 19138 28000 19168
rect 24761 19136 28000 19138
rect 24761 19080 24766 19136
rect 24822 19080 28000 19136
rect 24761 19078 28000 19080
rect 24761 19075 24827 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 21265 19002 21331 19005
rect 25497 19002 25563 19005
rect 21265 19000 25563 19002
rect 21265 18944 21270 19000
rect 21326 18944 25502 19000
rect 25558 18944 25563 19000
rect 21265 18942 25563 18944
rect 21265 18939 21331 18942
rect 25497 18939 25563 18942
rect 4337 18866 4403 18869
rect 11697 18866 11763 18869
rect 4337 18864 11763 18866
rect 4337 18808 4342 18864
rect 4398 18808 11702 18864
rect 11758 18808 11763 18864
rect 4337 18806 11763 18808
rect 4337 18803 4403 18806
rect 11697 18803 11763 18806
rect 24117 18866 24183 18869
rect 25589 18866 25655 18869
rect 24117 18864 25655 18866
rect 24117 18808 24122 18864
rect 24178 18808 25594 18864
rect 25650 18808 25655 18864
rect 24117 18806 25655 18808
rect 24117 18803 24183 18806
rect 25589 18803 25655 18806
rect 11421 18730 11487 18733
rect 20253 18730 20319 18733
rect 11421 18728 20319 18730
rect 11421 18672 11426 18728
rect 11482 18672 20258 18728
rect 20314 18672 20319 18728
rect 11421 18670 20319 18672
rect 11421 18667 11487 18670
rect 20253 18667 20319 18670
rect 22645 18730 22711 18733
rect 22645 18728 24778 18730
rect 22645 18672 22650 18728
rect 22706 18672 24778 18728
rect 22645 18670 24778 18672
rect 22645 18667 22711 18670
rect 24718 18594 24778 18670
rect 27520 18594 28000 18624
rect 24718 18534 28000 18594
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 27520 18504 28000 18534
rect 24277 18463 24597 18464
rect 14273 18458 14339 18461
rect 18781 18458 18847 18461
rect 24117 18458 24183 18461
rect 14273 18456 14474 18458
rect 14273 18400 14278 18456
rect 14334 18400 14474 18456
rect 14273 18398 14474 18400
rect 14273 18395 14339 18398
rect 14414 18322 14474 18398
rect 18781 18456 24183 18458
rect 18781 18400 18786 18456
rect 18842 18400 24122 18456
rect 24178 18400 24183 18456
rect 18781 18398 24183 18400
rect 18781 18395 18847 18398
rect 24117 18395 24183 18398
rect 14549 18322 14615 18325
rect 14414 18320 14615 18322
rect 14414 18264 14554 18320
rect 14610 18264 14615 18320
rect 14414 18262 14615 18264
rect 14549 18259 14615 18262
rect 17493 18322 17559 18325
rect 21173 18322 21239 18325
rect 21817 18322 21883 18325
rect 17493 18320 21883 18322
rect 17493 18264 17498 18320
rect 17554 18264 21178 18320
rect 21234 18264 21822 18320
rect 21878 18264 21883 18320
rect 17493 18262 21883 18264
rect 17493 18259 17559 18262
rect 21173 18259 21239 18262
rect 21817 18259 21883 18262
rect 1577 18186 1643 18189
rect 11421 18186 11487 18189
rect 1577 18184 11487 18186
rect 1577 18128 1582 18184
rect 1638 18128 11426 18184
rect 11482 18128 11487 18184
rect 1577 18126 11487 18128
rect 1577 18123 1643 18126
rect 11421 18123 11487 18126
rect 14365 18186 14431 18189
rect 15009 18186 15075 18189
rect 14365 18184 15075 18186
rect 14365 18128 14370 18184
rect 14426 18128 15014 18184
rect 15070 18128 15075 18184
rect 14365 18126 15075 18128
rect 14365 18123 14431 18126
rect 15009 18123 15075 18126
rect 16849 18186 16915 18189
rect 25221 18186 25287 18189
rect 16849 18184 25287 18186
rect 16849 18128 16854 18184
rect 16910 18128 25226 18184
rect 25282 18128 25287 18184
rect 16849 18126 25287 18128
rect 16849 18123 16915 18126
rect 25221 18123 25287 18126
rect 12249 18050 12315 18053
rect 17953 18050 18019 18053
rect 12249 18048 18019 18050
rect 12249 17992 12254 18048
rect 12310 17992 17958 18048
rect 18014 17992 18019 18048
rect 12249 17990 18019 17992
rect 12249 17987 12315 17990
rect 17953 17987 18019 17990
rect 25405 18050 25471 18053
rect 27520 18050 28000 18080
rect 25405 18048 28000 18050
rect 25405 17992 25410 18048
rect 25466 17992 28000 18048
rect 25405 17990 28000 17992
rect 25405 17987 25471 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 22553 17914 22619 17917
rect 25037 17914 25103 17917
rect 22553 17912 25103 17914
rect 22553 17856 22558 17912
rect 22614 17856 25042 17912
rect 25098 17856 25103 17912
rect 22553 17854 25103 17856
rect 22553 17851 22619 17854
rect 25037 17851 25103 17854
rect 14733 17778 14799 17781
rect 17953 17778 18019 17781
rect 14733 17776 18019 17778
rect 14733 17720 14738 17776
rect 14794 17720 17958 17776
rect 18014 17720 18019 17776
rect 14733 17718 18019 17720
rect 14733 17715 14799 17718
rect 17953 17715 18019 17718
rect 18229 17778 18295 17781
rect 21265 17778 21331 17781
rect 18229 17776 21331 17778
rect 18229 17720 18234 17776
rect 18290 17720 21270 17776
rect 21326 17720 21331 17776
rect 18229 17718 21331 17720
rect 18229 17715 18295 17718
rect 21265 17715 21331 17718
rect 12617 17642 12683 17645
rect 23565 17642 23631 17645
rect 12617 17640 23631 17642
rect 12617 17584 12622 17640
rect 12678 17584 23570 17640
rect 23626 17584 23631 17640
rect 12617 17582 23631 17584
rect 12617 17579 12683 17582
rect 23565 17579 23631 17582
rect 18965 17506 19031 17509
rect 20805 17506 20871 17509
rect 18965 17504 20871 17506
rect 18965 17448 18970 17504
rect 19026 17448 20810 17504
rect 20866 17448 20871 17504
rect 18965 17446 20871 17448
rect 18965 17443 19031 17446
rect 20805 17443 20871 17446
rect 25313 17506 25379 17509
rect 27520 17506 28000 17536
rect 25313 17504 28000 17506
rect 25313 17448 25318 17504
rect 25374 17448 28000 17504
rect 25313 17446 28000 17448
rect 25313 17443 25379 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 22461 17370 22527 17373
rect 17174 17368 22527 17370
rect 17174 17312 22466 17368
rect 22522 17312 22527 17368
rect 17174 17310 22527 17312
rect 11973 17234 12039 17237
rect 17174 17234 17234 17310
rect 22461 17307 22527 17310
rect 11973 17232 17234 17234
rect 11973 17176 11978 17232
rect 12034 17176 17234 17232
rect 11973 17174 17234 17176
rect 19977 17234 20043 17237
rect 25313 17234 25379 17237
rect 19977 17232 25379 17234
rect 19977 17176 19982 17232
rect 20038 17176 25318 17232
rect 25374 17176 25379 17232
rect 19977 17174 25379 17176
rect 11973 17171 12039 17174
rect 19977 17171 20043 17174
rect 25313 17171 25379 17174
rect 13445 17098 13511 17101
rect 21449 17098 21515 17101
rect 22369 17098 22435 17101
rect 25405 17098 25471 17101
rect 13445 17096 20132 17098
rect 13445 17040 13450 17096
rect 13506 17040 20132 17096
rect 13445 17038 20132 17040
rect 13445 17035 13511 17038
rect 13629 16962 13695 16965
rect 19241 16962 19307 16965
rect 13629 16960 19307 16962
rect 13629 16904 13634 16960
rect 13690 16904 19246 16960
rect 19302 16904 19307 16960
rect 13629 16902 19307 16904
rect 20072 16962 20132 17038
rect 21449 17096 25471 17098
rect 21449 17040 21454 17096
rect 21510 17040 22374 17096
rect 22430 17040 25410 17096
rect 25466 17040 25471 17096
rect 21449 17038 25471 17040
rect 21449 17035 21515 17038
rect 22369 17035 22435 17038
rect 25405 17035 25471 17038
rect 22553 16962 22619 16965
rect 24761 16962 24827 16965
rect 20072 16960 24827 16962
rect 20072 16904 22558 16960
rect 22614 16904 24766 16960
rect 24822 16904 24827 16960
rect 20072 16902 24827 16904
rect 13629 16899 13695 16902
rect 19241 16899 19307 16902
rect 22553 16899 22619 16902
rect 24761 16899 24827 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 10869 16826 10935 16829
rect 14457 16826 14523 16829
rect 10869 16824 14523 16826
rect 10869 16768 10874 16824
rect 10930 16768 14462 16824
rect 14518 16768 14523 16824
rect 10869 16766 14523 16768
rect 10869 16763 10935 16766
rect 14457 16763 14523 16766
rect 23473 16826 23539 16829
rect 27520 16826 28000 16856
rect 23473 16824 28000 16826
rect 23473 16768 23478 16824
rect 23534 16768 28000 16824
rect 23473 16766 28000 16768
rect 23473 16763 23539 16766
rect 27520 16736 28000 16766
rect 10869 16690 10935 16693
rect 12157 16690 12223 16693
rect 10869 16688 12223 16690
rect 10869 16632 10874 16688
rect 10930 16632 12162 16688
rect 12218 16632 12223 16688
rect 10869 16630 12223 16632
rect 10869 16627 10935 16630
rect 12157 16627 12223 16630
rect 16113 16690 16179 16693
rect 22645 16690 22711 16693
rect 16113 16688 22711 16690
rect 16113 16632 16118 16688
rect 16174 16632 22650 16688
rect 22706 16632 22711 16688
rect 16113 16630 22711 16632
rect 16113 16627 16179 16630
rect 22645 16627 22711 16630
rect 9949 16554 10015 16557
rect 23933 16554 23999 16557
rect 9949 16552 23999 16554
rect 9949 16496 9954 16552
rect 10010 16496 23938 16552
rect 23994 16496 23999 16552
rect 9949 16494 23999 16496
rect 9949 16491 10015 16494
rect 23933 16491 23999 16494
rect 19241 16418 19307 16421
rect 21173 16418 21239 16421
rect 19241 16416 21239 16418
rect 19241 16360 19246 16416
rect 19302 16360 21178 16416
rect 21234 16360 21239 16416
rect 19241 16358 21239 16360
rect 19241 16355 19307 16358
rect 21173 16355 21239 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 8201 16282 8267 16285
rect 13721 16282 13787 16285
rect 8201 16280 13787 16282
rect 8201 16224 8206 16280
rect 8262 16224 13726 16280
rect 13782 16224 13787 16280
rect 8201 16222 13787 16224
rect 8201 16219 8267 16222
rect 13721 16219 13787 16222
rect 16113 16282 16179 16285
rect 23657 16282 23723 16285
rect 27520 16282 28000 16312
rect 16113 16280 23723 16282
rect 16113 16224 16118 16280
rect 16174 16224 23662 16280
rect 23718 16224 23723 16280
rect 16113 16222 23723 16224
rect 16113 16219 16179 16222
rect 23657 16219 23723 16222
rect 24902 16222 28000 16282
rect 19885 16146 19951 16149
rect 24902 16146 24962 16222
rect 27520 16192 28000 16222
rect 19885 16144 24962 16146
rect 19885 16088 19890 16144
rect 19946 16088 24962 16144
rect 19885 16086 24962 16088
rect 19885 16083 19951 16086
rect 14825 16010 14891 16013
rect 17493 16010 17559 16013
rect 14825 16008 17559 16010
rect 14825 15952 14830 16008
rect 14886 15952 17498 16008
rect 17554 15952 17559 16008
rect 14825 15950 17559 15952
rect 14825 15947 14891 15950
rect 17493 15947 17559 15950
rect 21173 16010 21239 16013
rect 22277 16010 22343 16013
rect 21173 16008 22343 16010
rect 21173 15952 21178 16008
rect 21234 15952 22282 16008
rect 22338 15952 22343 16008
rect 21173 15950 22343 15952
rect 21173 15947 21239 15950
rect 22277 15947 22343 15950
rect 10685 15874 10751 15877
rect 15653 15874 15719 15877
rect 10685 15872 15719 15874
rect 10685 15816 10690 15872
rect 10746 15816 15658 15872
rect 15714 15816 15719 15872
rect 10685 15814 15719 15816
rect 10685 15811 10751 15814
rect 15653 15811 15719 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 14733 15738 14799 15741
rect 16205 15738 16271 15741
rect 17769 15738 17835 15741
rect 14733 15736 16271 15738
rect 14733 15680 14738 15736
rect 14794 15680 16210 15736
rect 16266 15680 16271 15736
rect 14733 15678 16271 15680
rect 14733 15675 14799 15678
rect 16205 15675 16271 15678
rect 17358 15736 17835 15738
rect 17358 15680 17774 15736
rect 17830 15680 17835 15736
rect 17358 15678 17835 15680
rect 13537 15602 13603 15605
rect 16573 15602 16639 15605
rect 17358 15602 17418 15678
rect 17769 15675 17835 15678
rect 24117 15738 24183 15741
rect 27520 15738 28000 15768
rect 24117 15736 28000 15738
rect 24117 15680 24122 15736
rect 24178 15680 28000 15736
rect 24117 15678 28000 15680
rect 24117 15675 24183 15678
rect 27520 15648 28000 15678
rect 13537 15600 17418 15602
rect 13537 15544 13542 15600
rect 13598 15544 16578 15600
rect 16634 15544 17418 15600
rect 13537 15542 17418 15544
rect 17493 15602 17559 15605
rect 18505 15602 18571 15605
rect 17493 15600 18571 15602
rect 17493 15544 17498 15600
rect 17554 15544 18510 15600
rect 18566 15544 18571 15600
rect 17493 15542 18571 15544
rect 13537 15539 13603 15542
rect 16573 15539 16639 15542
rect 17493 15539 17559 15542
rect 18505 15539 18571 15542
rect 4061 15466 4127 15469
rect 21725 15466 21791 15469
rect 4061 15464 21791 15466
rect 4061 15408 4066 15464
rect 4122 15408 21730 15464
rect 21786 15408 21791 15464
rect 4061 15406 21791 15408
rect 4061 15403 4127 15406
rect 21725 15403 21791 15406
rect 10041 15330 10107 15333
rect 13537 15330 13603 15333
rect 10041 15328 13603 15330
rect 10041 15272 10046 15328
rect 10102 15272 13542 15328
rect 13598 15272 13603 15328
rect 10041 15270 13603 15272
rect 10041 15267 10107 15270
rect 13537 15267 13603 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 24761 15194 24827 15197
rect 27520 15194 28000 15224
rect 24761 15192 28000 15194
rect 24761 15136 24766 15192
rect 24822 15136 28000 15192
rect 24761 15134 28000 15136
rect 24761 15131 24827 15134
rect 27520 15104 28000 15134
rect 11421 15058 11487 15061
rect 15561 15058 15627 15061
rect 11421 15056 15627 15058
rect 11421 15000 11426 15056
rect 11482 15000 15566 15056
rect 15622 15000 15627 15056
rect 11421 14998 15627 15000
rect 11421 14995 11487 14998
rect 15561 14995 15627 14998
rect 19609 15058 19675 15061
rect 22461 15058 22527 15061
rect 19609 15056 22527 15058
rect 19609 15000 19614 15056
rect 19670 15000 22466 15056
rect 22522 15000 22527 15056
rect 19609 14998 22527 15000
rect 19609 14995 19675 14998
rect 22461 14995 22527 14998
rect 12893 14922 12959 14925
rect 18873 14922 18939 14925
rect 21817 14922 21883 14925
rect 12893 14920 21883 14922
rect 12893 14864 12898 14920
rect 12954 14864 18878 14920
rect 18934 14864 21822 14920
rect 21878 14864 21883 14920
rect 12893 14862 21883 14864
rect 12893 14859 12959 14862
rect 18873 14859 18939 14862
rect 21817 14859 21883 14862
rect 16481 14786 16547 14789
rect 17677 14786 17743 14789
rect 18505 14786 18571 14789
rect 16481 14784 18571 14786
rect 16481 14728 16486 14784
rect 16542 14728 17682 14784
rect 17738 14728 18510 14784
rect 18566 14728 18571 14784
rect 16481 14726 18571 14728
rect 16481 14723 16547 14726
rect 17677 14723 17743 14726
rect 18505 14723 18571 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 12249 14650 12315 14653
rect 13997 14650 14063 14653
rect 18045 14650 18111 14653
rect 12249 14648 18111 14650
rect 12249 14592 12254 14648
rect 12310 14592 14002 14648
rect 14058 14592 18050 14648
rect 18106 14592 18111 14648
rect 12249 14590 18111 14592
rect 12249 14587 12315 14590
rect 13997 14587 14063 14590
rect 18045 14587 18111 14590
rect 23841 14650 23907 14653
rect 27520 14650 28000 14680
rect 23841 14648 28000 14650
rect 23841 14592 23846 14648
rect 23902 14592 28000 14648
rect 23841 14590 28000 14592
rect 23841 14587 23907 14590
rect 27520 14560 28000 14590
rect 15929 14514 15995 14517
rect 22185 14514 22251 14517
rect 15929 14512 22251 14514
rect 15929 14456 15934 14512
rect 15990 14456 22190 14512
rect 22246 14456 22251 14512
rect 15929 14454 22251 14456
rect 15929 14451 15995 14454
rect 22185 14451 22251 14454
rect 10133 14242 10199 14245
rect 13445 14242 13511 14245
rect 10133 14240 13511 14242
rect 10133 14184 10138 14240
rect 10194 14184 13450 14240
rect 13506 14184 13511 14240
rect 10133 14182 13511 14184
rect 10133 14179 10199 14182
rect 13445 14179 13511 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 10777 14106 10843 14109
rect 14641 14106 14707 14109
rect 10777 14104 14707 14106
rect 10777 14048 10782 14104
rect 10838 14048 14646 14104
rect 14702 14048 14707 14104
rect 10777 14046 14707 14048
rect 10777 14043 10843 14046
rect 14641 14043 14707 14046
rect 17217 14106 17283 14109
rect 17585 14106 17651 14109
rect 20069 14106 20135 14109
rect 17217 14104 20135 14106
rect 17217 14048 17222 14104
rect 17278 14048 17590 14104
rect 17646 14048 20074 14104
rect 20130 14048 20135 14104
rect 17217 14046 20135 14048
rect 17217 14043 17283 14046
rect 17585 14043 17651 14046
rect 20069 14043 20135 14046
rect 15101 13970 15167 13973
rect 16757 13970 16823 13973
rect 15101 13968 16823 13970
rect 15101 13912 15106 13968
rect 15162 13912 16762 13968
rect 16818 13912 16823 13968
rect 15101 13910 16823 13912
rect 15101 13907 15167 13910
rect 16757 13907 16823 13910
rect 21173 13970 21239 13973
rect 27520 13970 28000 14000
rect 21173 13968 28000 13970
rect 21173 13912 21178 13968
rect 21234 13912 28000 13968
rect 21173 13910 28000 13912
rect 21173 13907 21239 13910
rect 27520 13880 28000 13910
rect 14181 13834 14247 13837
rect 18965 13834 19031 13837
rect 14181 13832 19031 13834
rect 14181 13776 14186 13832
rect 14242 13776 18970 13832
rect 19026 13776 19031 13832
rect 14181 13774 19031 13776
rect 14181 13771 14247 13774
rect 18965 13771 19031 13774
rect 22001 13834 22067 13837
rect 25037 13834 25103 13837
rect 22001 13832 25103 13834
rect 22001 13776 22006 13832
rect 22062 13776 25042 13832
rect 25098 13776 25103 13832
rect 22001 13774 25103 13776
rect 22001 13771 22067 13774
rect 25037 13771 25103 13774
rect 11513 13698 11579 13701
rect 17309 13698 17375 13701
rect 11513 13696 17375 13698
rect 11513 13640 11518 13696
rect 11574 13640 17314 13696
rect 17370 13640 17375 13696
rect 11513 13638 17375 13640
rect 11513 13635 11579 13638
rect 17309 13635 17375 13638
rect 17861 13698 17927 13701
rect 19425 13698 19491 13701
rect 17861 13696 19491 13698
rect 17861 13640 17866 13696
rect 17922 13640 19430 13696
rect 19486 13640 19491 13696
rect 17861 13638 19491 13640
rect 17861 13635 17927 13638
rect 19425 13635 19491 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 14457 13562 14523 13565
rect 16849 13562 16915 13565
rect 14457 13560 16915 13562
rect 14457 13504 14462 13560
rect 14518 13504 16854 13560
rect 16910 13504 16915 13560
rect 14457 13502 16915 13504
rect 14457 13499 14523 13502
rect 16849 13499 16915 13502
rect 20437 13562 20503 13565
rect 24117 13562 24183 13565
rect 20437 13560 24183 13562
rect 20437 13504 20442 13560
rect 20498 13504 24122 13560
rect 24178 13504 24183 13560
rect 20437 13502 24183 13504
rect 20437 13499 20503 13502
rect 24117 13499 24183 13502
rect 22921 13426 22987 13429
rect 22878 13424 22987 13426
rect 22878 13368 22926 13424
rect 22982 13368 22987 13424
rect 22878 13363 22987 13368
rect 24117 13426 24183 13429
rect 27520 13426 28000 13456
rect 24117 13424 28000 13426
rect 24117 13368 24122 13424
rect 24178 13368 28000 13424
rect 24117 13366 28000 13368
rect 24117 13363 24183 13366
rect 14641 13290 14707 13293
rect 22878 13290 22938 13363
rect 27520 13336 28000 13366
rect 25313 13290 25379 13293
rect 14641 13288 25379 13290
rect 14641 13232 14646 13288
rect 14702 13232 25318 13288
rect 25374 13232 25379 13288
rect 14641 13230 25379 13232
rect 14641 13227 14707 13230
rect 25313 13227 25379 13230
rect 15561 13154 15627 13157
rect 23841 13154 23907 13157
rect 15561 13152 23907 13154
rect 15561 13096 15566 13152
rect 15622 13096 23846 13152
rect 23902 13096 23907 13152
rect 15561 13094 23907 13096
rect 15561 13091 15627 13094
rect 23841 13091 23907 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 17677 13018 17743 13021
rect 20437 13018 20503 13021
rect 17677 13016 20503 13018
rect 17677 12960 17682 13016
rect 17738 12960 20442 13016
rect 20498 12960 20503 13016
rect 17677 12958 20503 12960
rect 17677 12955 17743 12958
rect 20437 12955 20503 12958
rect 17585 12882 17651 12885
rect 19701 12882 19767 12885
rect 17585 12880 19767 12882
rect 17585 12824 17590 12880
rect 17646 12824 19706 12880
rect 19762 12824 19767 12880
rect 17585 12822 19767 12824
rect 17585 12819 17651 12822
rect 19701 12819 19767 12822
rect 23933 12882 23999 12885
rect 27520 12882 28000 12912
rect 23933 12880 28000 12882
rect 23933 12824 23938 12880
rect 23994 12824 28000 12880
rect 23933 12822 28000 12824
rect 23933 12819 23999 12822
rect 27520 12792 28000 12822
rect 20897 12746 20963 12749
rect 21541 12746 21607 12749
rect 19382 12744 21607 12746
rect 19382 12688 20902 12744
rect 20958 12688 21546 12744
rect 21602 12688 21607 12744
rect 19382 12686 21607 12688
rect 11237 12610 11303 12613
rect 18229 12610 18295 12613
rect 18965 12610 19031 12613
rect 11237 12608 19031 12610
rect 11237 12552 11242 12608
rect 11298 12552 18234 12608
rect 18290 12552 18970 12608
rect 19026 12552 19031 12608
rect 11237 12550 19031 12552
rect 11237 12547 11303 12550
rect 18229 12547 18295 12550
rect 18965 12547 19031 12550
rect 19149 12610 19215 12613
rect 19382 12610 19442 12686
rect 20897 12683 20963 12686
rect 21541 12683 21607 12686
rect 19149 12608 19442 12610
rect 19149 12552 19154 12608
rect 19210 12552 19442 12608
rect 19149 12550 19442 12552
rect 20161 12610 20227 12613
rect 20713 12610 20779 12613
rect 20161 12608 20779 12610
rect 20161 12552 20166 12608
rect 20222 12552 20718 12608
rect 20774 12552 20779 12608
rect 20161 12550 20779 12552
rect 19149 12547 19215 12550
rect 20161 12547 20227 12550
rect 20713 12547 20779 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 21081 12474 21147 12477
rect 22461 12474 22527 12477
rect 23749 12474 23815 12477
rect 21081 12472 23815 12474
rect 21081 12416 21086 12472
rect 21142 12416 22466 12472
rect 22522 12416 23754 12472
rect 23810 12416 23815 12472
rect 21081 12414 23815 12416
rect 21081 12411 21147 12414
rect 22461 12411 22527 12414
rect 23749 12411 23815 12414
rect 18873 12338 18939 12341
rect 23105 12338 23171 12341
rect 18873 12336 23171 12338
rect 18873 12280 18878 12336
rect 18934 12280 23110 12336
rect 23166 12280 23171 12336
rect 18873 12278 23171 12280
rect 18873 12275 18939 12278
rect 23105 12275 23171 12278
rect 24761 12338 24827 12341
rect 27520 12338 28000 12368
rect 24761 12336 28000 12338
rect 24761 12280 24766 12336
rect 24822 12280 28000 12336
rect 24761 12278 28000 12280
rect 24761 12275 24827 12278
rect 27520 12248 28000 12278
rect 10961 12202 11027 12205
rect 18137 12202 18203 12205
rect 10961 12200 18203 12202
rect 10961 12144 10966 12200
rect 11022 12144 18142 12200
rect 18198 12144 18203 12200
rect 10961 12142 18203 12144
rect 10961 12139 11027 12142
rect 18137 12139 18203 12142
rect 19885 12202 19951 12205
rect 22185 12202 22251 12205
rect 24577 12202 24643 12205
rect 19885 12200 22251 12202
rect 19885 12144 19890 12200
rect 19946 12144 22190 12200
rect 22246 12144 22251 12200
rect 19885 12142 22251 12144
rect 19885 12139 19951 12142
rect 22185 12139 22251 12142
rect 23246 12200 24643 12202
rect 23246 12144 24582 12200
rect 24638 12144 24643 12200
rect 23246 12142 24643 12144
rect 15377 12066 15443 12069
rect 19057 12066 19123 12069
rect 15377 12064 19123 12066
rect 15377 12008 15382 12064
rect 15438 12008 19062 12064
rect 19118 12008 19123 12064
rect 15377 12006 19123 12008
rect 15377 12003 15443 12006
rect 19057 12003 19123 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 18045 11930 18111 11933
rect 23246 11930 23306 12142
rect 24577 12139 24643 12142
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 23841 11932 23907 11933
rect 23790 11930 23796 11932
rect 18045 11928 23306 11930
rect 18045 11872 18050 11928
rect 18106 11872 23306 11928
rect 18045 11870 23306 11872
rect 23750 11870 23796 11930
rect 23860 11928 23907 11932
rect 23902 11872 23907 11928
rect 18045 11867 18111 11870
rect 23790 11868 23796 11870
rect 23860 11868 23907 11872
rect 23841 11867 23907 11868
rect 12157 11794 12223 11797
rect 17769 11794 17835 11797
rect 12157 11792 17835 11794
rect 12157 11736 12162 11792
rect 12218 11736 17774 11792
rect 17830 11736 17835 11792
rect 12157 11734 17835 11736
rect 12157 11731 12223 11734
rect 17769 11731 17835 11734
rect 21357 11794 21423 11797
rect 27520 11794 28000 11824
rect 21357 11792 28000 11794
rect 21357 11736 21362 11792
rect 21418 11736 28000 11792
rect 21357 11734 28000 11736
rect 21357 11731 21423 11734
rect 27520 11704 28000 11734
rect 381 11658 447 11661
rect 11053 11658 11119 11661
rect 381 11656 11119 11658
rect 381 11600 386 11656
rect 442 11600 11058 11656
rect 11114 11600 11119 11656
rect 381 11598 11119 11600
rect 381 11595 447 11598
rect 11053 11595 11119 11598
rect 13905 11658 13971 11661
rect 14457 11658 14523 11661
rect 13905 11656 14523 11658
rect 13905 11600 13910 11656
rect 13966 11600 14462 11656
rect 14518 11600 14523 11656
rect 13905 11598 14523 11600
rect 13905 11595 13971 11598
rect 14457 11595 14523 11598
rect 19241 11658 19307 11661
rect 20897 11658 20963 11661
rect 19241 11656 20963 11658
rect 19241 11600 19246 11656
rect 19302 11600 20902 11656
rect 20958 11600 20963 11656
rect 19241 11598 20963 11600
rect 19241 11595 19307 11598
rect 20897 11595 20963 11598
rect 20069 11522 20135 11525
rect 24117 11522 24183 11525
rect 20069 11520 24183 11522
rect 20069 11464 20074 11520
rect 20130 11464 24122 11520
rect 24178 11464 24183 11520
rect 20069 11462 24183 11464
rect 20069 11459 20135 11462
rect 24117 11459 24183 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 12249 11386 12315 11389
rect 17585 11386 17651 11389
rect 18045 11386 18111 11389
rect 12249 11384 18111 11386
rect 12249 11328 12254 11384
rect 12310 11328 17590 11384
rect 17646 11328 18050 11384
rect 18106 11328 18111 11384
rect 12249 11326 18111 11328
rect 12249 11323 12315 11326
rect 17585 11323 17651 11326
rect 18045 11323 18111 11326
rect 13629 11114 13695 11117
rect 15009 11114 15075 11117
rect 13629 11112 15075 11114
rect 13629 11056 13634 11112
rect 13690 11056 15014 11112
rect 15070 11056 15075 11112
rect 13629 11054 15075 11056
rect 13629 11051 13695 11054
rect 15009 11051 15075 11054
rect 18413 11114 18479 11117
rect 27520 11114 28000 11144
rect 18413 11112 28000 11114
rect 18413 11056 18418 11112
rect 18474 11056 28000 11112
rect 18413 11054 28000 11056
rect 18413 11051 18479 11054
rect 27520 11024 28000 11054
rect 21817 10978 21883 10981
rect 23013 10978 23079 10981
rect 21817 10976 23079 10978
rect 21817 10920 21822 10976
rect 21878 10920 23018 10976
rect 23074 10920 23079 10976
rect 21817 10918 23079 10920
rect 21817 10915 21883 10918
rect 23013 10915 23079 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 15653 10842 15719 10845
rect 15653 10840 24042 10842
rect 15653 10784 15658 10840
rect 15714 10784 24042 10840
rect 15653 10782 24042 10784
rect 15653 10779 15719 10782
rect 19241 10706 19307 10709
rect 19885 10706 19951 10709
rect 22737 10706 22803 10709
rect 19241 10704 22803 10706
rect 19241 10648 19246 10704
rect 19302 10648 19890 10704
rect 19946 10648 22742 10704
rect 22798 10648 22803 10704
rect 19241 10646 22803 10648
rect 19241 10643 19307 10646
rect 19885 10643 19951 10646
rect 22737 10643 22803 10646
rect 16665 10570 16731 10573
rect 21265 10570 21331 10573
rect 16665 10568 21331 10570
rect 16665 10512 16670 10568
rect 16726 10512 21270 10568
rect 21326 10512 21331 10568
rect 16665 10510 21331 10512
rect 16665 10507 16731 10510
rect 21265 10507 21331 10510
rect 13721 10434 13787 10437
rect 17953 10434 18019 10437
rect 13721 10432 18019 10434
rect 13721 10376 13726 10432
rect 13782 10376 17958 10432
rect 18014 10376 18019 10432
rect 13721 10374 18019 10376
rect 13721 10371 13787 10374
rect 17953 10371 18019 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 10777 10298 10843 10301
rect 15009 10298 15075 10301
rect 10777 10296 15075 10298
rect 10777 10240 10782 10296
rect 10838 10240 15014 10296
rect 15070 10240 15075 10296
rect 10777 10238 15075 10240
rect 10777 10235 10843 10238
rect 15009 10235 15075 10238
rect 1393 10162 1459 10165
rect 4981 10162 5047 10165
rect 12065 10162 12131 10165
rect 1393 10160 4906 10162
rect 1393 10104 1398 10160
rect 1454 10104 4906 10160
rect 1393 10102 4906 10104
rect 1393 10099 1459 10102
rect 4846 10026 4906 10102
rect 4981 10160 12131 10162
rect 4981 10104 4986 10160
rect 5042 10104 12070 10160
rect 12126 10104 12131 10160
rect 4981 10102 12131 10104
rect 4981 10099 5047 10102
rect 12065 10099 12131 10102
rect 12249 10162 12315 10165
rect 20345 10162 20411 10165
rect 12249 10160 20411 10162
rect 12249 10104 12254 10160
rect 12310 10104 20350 10160
rect 20406 10104 20411 10160
rect 12249 10102 20411 10104
rect 12249 10099 12315 10102
rect 20345 10099 20411 10102
rect 9949 10026 10015 10029
rect 11881 10026 11947 10029
rect 18321 10026 18387 10029
rect 20805 10026 20871 10029
rect 4846 10024 11714 10026
rect 4846 9968 9954 10024
rect 10010 9968 11714 10024
rect 4846 9966 11714 9968
rect 9949 9963 10015 9966
rect 11654 9890 11714 9966
rect 11881 10024 16130 10026
rect 11881 9968 11886 10024
rect 11942 9968 16130 10024
rect 11881 9966 16130 9968
rect 11881 9963 11947 9966
rect 12249 9890 12315 9893
rect 11654 9888 12315 9890
rect 11654 9832 12254 9888
rect 12310 9832 12315 9888
rect 11654 9830 12315 9832
rect 12249 9827 12315 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 16070 9754 16130 9966
rect 18321 10024 20871 10026
rect 18321 9968 18326 10024
rect 18382 9968 20810 10024
rect 20866 9968 20871 10024
rect 18321 9966 20871 9968
rect 23982 10026 24042 10782
rect 24117 10570 24183 10573
rect 27520 10570 28000 10600
rect 24117 10568 28000 10570
rect 24117 10512 24122 10568
rect 24178 10512 28000 10568
rect 24117 10510 28000 10512
rect 24117 10507 24183 10510
rect 27520 10480 28000 10510
rect 27520 10026 28000 10056
rect 23982 9966 28000 10026
rect 18321 9963 18387 9966
rect 20805 9963 20871 9966
rect 27520 9936 28000 9966
rect 16297 9890 16363 9893
rect 24117 9890 24183 9893
rect 16297 9888 24183 9890
rect 16297 9832 16302 9888
rect 16358 9832 24122 9888
rect 24178 9832 24183 9888
rect 16297 9830 24183 9832
rect 16297 9827 16363 9830
rect 24117 9827 24183 9830
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 16389 9754 16455 9757
rect 18321 9754 18387 9757
rect 21173 9754 21239 9757
rect 16070 9694 16314 9754
rect 13445 9618 13511 9621
rect 13905 9618 13971 9621
rect 13445 9616 13971 9618
rect 13445 9560 13450 9616
rect 13506 9560 13910 9616
rect 13966 9560 13971 9616
rect 13445 9558 13971 9560
rect 16254 9618 16314 9694
rect 16389 9752 18387 9754
rect 16389 9696 16394 9752
rect 16450 9696 18326 9752
rect 18382 9696 18387 9752
rect 16389 9694 18387 9696
rect 16389 9691 16455 9694
rect 18321 9691 18387 9694
rect 18462 9752 21239 9754
rect 18462 9696 21178 9752
rect 21234 9696 21239 9752
rect 18462 9694 21239 9696
rect 16389 9618 16455 9621
rect 18462 9618 18522 9694
rect 21173 9691 21239 9694
rect 16254 9616 18522 9618
rect 16254 9560 16394 9616
rect 16450 9560 18522 9616
rect 16254 9558 18522 9560
rect 19885 9618 19951 9621
rect 23473 9618 23539 9621
rect 19885 9616 23539 9618
rect 19885 9560 19890 9616
rect 19946 9560 23478 9616
rect 23534 9560 23539 9616
rect 19885 9558 23539 9560
rect 13445 9555 13511 9558
rect 13905 9555 13971 9558
rect 16389 9555 16455 9558
rect 19885 9555 19951 9558
rect 23473 9555 23539 9558
rect 15561 9484 15627 9485
rect 15510 9482 15516 9484
rect 15470 9422 15516 9482
rect 15580 9480 15627 9484
rect 15622 9424 15627 9480
rect 15510 9420 15516 9422
rect 15580 9420 15627 9424
rect 15561 9419 15627 9420
rect 24761 9482 24827 9485
rect 27520 9482 28000 9512
rect 24761 9480 28000 9482
rect 24761 9424 24766 9480
rect 24822 9424 28000 9480
rect 24761 9422 28000 9424
rect 24761 9419 24827 9422
rect 27520 9392 28000 9422
rect 11145 9346 11211 9349
rect 15377 9346 15443 9349
rect 15653 9346 15719 9349
rect 11145 9344 15719 9346
rect 11145 9288 11150 9344
rect 11206 9288 15382 9344
rect 15438 9288 15658 9344
rect 15714 9288 15719 9344
rect 11145 9286 15719 9288
rect 11145 9283 11211 9286
rect 15377 9283 15443 9286
rect 15653 9283 15719 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 11605 9210 11671 9213
rect 17217 9210 17283 9213
rect 11605 9208 17283 9210
rect 11605 9152 11610 9208
rect 11666 9152 17222 9208
rect 17278 9152 17283 9208
rect 11605 9150 17283 9152
rect 11605 9147 11671 9150
rect 17217 9147 17283 9150
rect 12341 9074 12407 9077
rect 16021 9074 16087 9077
rect 12341 9072 16087 9074
rect 12341 9016 12346 9072
rect 12402 9016 16026 9072
rect 16082 9016 16087 9072
rect 12341 9014 16087 9016
rect 12341 9011 12407 9014
rect 16021 9011 16087 9014
rect 17493 8938 17559 8941
rect 19425 8938 19491 8941
rect 17493 8936 19491 8938
rect 17493 8880 17498 8936
rect 17554 8880 19430 8936
rect 19486 8880 19491 8936
rect 17493 8878 19491 8880
rect 17493 8875 17559 8878
rect 19425 8875 19491 8878
rect 23841 8938 23907 8941
rect 27520 8938 28000 8968
rect 23841 8936 28000 8938
rect 23841 8880 23846 8936
rect 23902 8880 28000 8936
rect 23841 8878 28000 8880
rect 23841 8875 23907 8878
rect 27520 8848 28000 8878
rect 15469 8802 15535 8805
rect 23013 8802 23079 8805
rect 15469 8800 23079 8802
rect 15469 8744 15474 8800
rect 15530 8744 23018 8800
rect 23074 8744 23079 8800
rect 15469 8742 23079 8744
rect 15469 8739 15535 8742
rect 23013 8739 23079 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 13997 8530 14063 8533
rect 22277 8530 22343 8533
rect 23841 8530 23907 8533
rect 13997 8528 17418 8530
rect 13997 8472 14002 8528
rect 14058 8472 17418 8528
rect 13997 8470 17418 8472
rect 13997 8467 14063 8470
rect 10685 8394 10751 8397
rect 12433 8394 12499 8397
rect 10685 8392 12499 8394
rect 10685 8336 10690 8392
rect 10746 8336 12438 8392
rect 12494 8336 12499 8392
rect 10685 8334 12499 8336
rect 10685 8331 10751 8334
rect 12433 8331 12499 8334
rect 14273 8394 14339 8397
rect 17125 8394 17191 8397
rect 14273 8392 17191 8394
rect 14273 8336 14278 8392
rect 14334 8336 17130 8392
rect 17186 8336 17191 8392
rect 14273 8334 17191 8336
rect 17358 8394 17418 8470
rect 22277 8528 23907 8530
rect 22277 8472 22282 8528
rect 22338 8472 23846 8528
rect 23902 8472 23907 8528
rect 22277 8470 23907 8472
rect 22277 8467 22343 8470
rect 23841 8467 23907 8470
rect 18689 8394 18755 8397
rect 20621 8394 20687 8397
rect 22277 8394 22343 8397
rect 17358 8392 22343 8394
rect 17358 8336 18694 8392
rect 18750 8336 20626 8392
rect 20682 8336 22282 8392
rect 22338 8336 22343 8392
rect 17358 8334 22343 8336
rect 14273 8331 14339 8334
rect 17125 8331 17191 8334
rect 18689 8331 18755 8334
rect 20621 8331 20687 8334
rect 22277 8331 22343 8334
rect 11421 8258 11487 8261
rect 11789 8258 11855 8261
rect 11421 8256 11855 8258
rect 11421 8200 11426 8256
rect 11482 8200 11794 8256
rect 11850 8200 11855 8256
rect 11421 8198 11855 8200
rect 11421 8195 11487 8198
rect 11789 8195 11855 8198
rect 12617 8258 12683 8261
rect 18137 8258 18203 8261
rect 12617 8256 18203 8258
rect 12617 8200 12622 8256
rect 12678 8200 18142 8256
rect 18198 8200 18203 8256
rect 12617 8198 18203 8200
rect 12617 8195 12683 8198
rect 18137 8195 18203 8198
rect 20069 8258 20135 8261
rect 23289 8258 23355 8261
rect 20069 8256 23355 8258
rect 20069 8200 20074 8256
rect 20130 8200 23294 8256
rect 23350 8200 23355 8256
rect 20069 8198 23355 8200
rect 20069 8195 20135 8198
rect 23289 8195 23355 8198
rect 24209 8258 24275 8261
rect 27520 8258 28000 8288
rect 24209 8256 28000 8258
rect 24209 8200 24214 8256
rect 24270 8200 28000 8256
rect 24209 8198 28000 8200
rect 24209 8195 24275 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 289 8122 355 8125
rect 11973 8122 12039 8125
rect 14365 8122 14431 8125
rect 289 8120 7666 8122
rect 289 8064 294 8120
rect 350 8064 7666 8120
rect 289 8062 7666 8064
rect 289 8059 355 8062
rect 7606 7986 7666 8062
rect 11973 8120 14431 8122
rect 11973 8064 11978 8120
rect 12034 8064 14370 8120
rect 14426 8064 14431 8120
rect 11973 8062 14431 8064
rect 11973 8059 12039 8062
rect 14365 8059 14431 8062
rect 21081 8122 21147 8125
rect 22185 8122 22251 8125
rect 21081 8120 22251 8122
rect 21081 8064 21086 8120
rect 21142 8064 22190 8120
rect 22246 8064 22251 8120
rect 21081 8062 22251 8064
rect 21081 8059 21147 8062
rect 22185 8059 22251 8062
rect 23473 8122 23539 8125
rect 23473 8120 25146 8122
rect 23473 8064 23478 8120
rect 23534 8064 25146 8120
rect 23473 8062 25146 8064
rect 23473 8059 23539 8062
rect 14733 7986 14799 7989
rect 15469 7986 15535 7989
rect 18873 7986 18939 7989
rect 19149 7986 19215 7989
rect 24761 7986 24827 7989
rect 7606 7984 18706 7986
rect 7606 7928 14738 7984
rect 14794 7928 15474 7984
rect 15530 7928 18706 7984
rect 7606 7926 18706 7928
rect 14733 7923 14799 7926
rect 15469 7923 15535 7926
rect 3693 7850 3759 7853
rect 11237 7850 11303 7853
rect 3693 7848 11303 7850
rect 3693 7792 3698 7848
rect 3754 7792 11242 7848
rect 11298 7792 11303 7848
rect 3693 7790 11303 7792
rect 3693 7787 3759 7790
rect 11237 7787 11303 7790
rect 13721 7850 13787 7853
rect 18646 7850 18706 7926
rect 18873 7984 24827 7986
rect 18873 7928 18878 7984
rect 18934 7928 19154 7984
rect 19210 7928 24766 7984
rect 24822 7928 24827 7984
rect 18873 7926 24827 7928
rect 18873 7923 18939 7926
rect 19149 7923 19215 7926
rect 24761 7923 24827 7926
rect 19609 7850 19675 7853
rect 13721 7848 18522 7850
rect 13721 7792 13726 7848
rect 13782 7792 18522 7848
rect 13721 7790 18522 7792
rect 18646 7848 19675 7850
rect 18646 7792 19614 7848
rect 19670 7792 19675 7848
rect 18646 7790 19675 7792
rect 13721 7787 13787 7790
rect 9765 7714 9831 7717
rect 12525 7714 12591 7717
rect 9765 7712 12591 7714
rect 9765 7656 9770 7712
rect 9826 7656 12530 7712
rect 12586 7656 12591 7712
rect 9765 7654 12591 7656
rect 18462 7714 18522 7790
rect 19609 7787 19675 7790
rect 19793 7850 19859 7853
rect 19793 7848 24962 7850
rect 19793 7792 19798 7848
rect 19854 7792 24962 7848
rect 19793 7790 24962 7792
rect 19793 7787 19859 7790
rect 21265 7714 21331 7717
rect 18462 7712 21331 7714
rect 18462 7656 21270 7712
rect 21326 7656 21331 7712
rect 18462 7654 21331 7656
rect 9765 7651 9831 7654
rect 12525 7651 12591 7654
rect 21265 7651 21331 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 16757 7578 16823 7581
rect 16757 7576 24042 7578
rect 16757 7520 16762 7576
rect 16818 7520 24042 7576
rect 16757 7518 24042 7520
rect 16757 7515 16823 7518
rect 17585 7442 17651 7445
rect 21081 7442 21147 7445
rect 17585 7440 21147 7442
rect 17585 7384 17590 7440
rect 17646 7384 21086 7440
rect 21142 7384 21147 7440
rect 17585 7382 21147 7384
rect 23982 7442 24042 7518
rect 24761 7442 24827 7445
rect 23982 7440 24827 7442
rect 23982 7384 24766 7440
rect 24822 7384 24827 7440
rect 23982 7382 24827 7384
rect 17585 7379 17651 7382
rect 21081 7379 21147 7382
rect 24761 7379 24827 7382
rect 2313 7306 2379 7309
rect 10317 7306 10383 7309
rect 2313 7304 10383 7306
rect 2313 7248 2318 7304
rect 2374 7248 10322 7304
rect 10378 7248 10383 7304
rect 2313 7246 10383 7248
rect 2313 7243 2379 7246
rect 10317 7243 10383 7246
rect 16941 7306 17007 7309
rect 19517 7306 19583 7309
rect 16941 7304 19583 7306
rect 16941 7248 16946 7304
rect 17002 7248 19522 7304
rect 19578 7248 19583 7304
rect 16941 7246 19583 7248
rect 16941 7243 17007 7246
rect 19517 7243 19583 7246
rect 24902 7170 24962 7790
rect 25086 7714 25146 8062
rect 27520 7714 28000 7744
rect 25086 7654 28000 7714
rect 27520 7624 28000 7654
rect 27520 7170 28000 7200
rect 24902 7110 28000 7170
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 27520 7080 28000 7110
rect 19610 7039 19930 7040
rect 11053 7034 11119 7037
rect 11789 7034 11855 7037
rect 17217 7034 17283 7037
rect 0 6974 3986 7034
rect 0 6944 480 6974
rect 3926 6898 3986 6974
rect 11053 7032 17283 7034
rect 11053 6976 11058 7032
rect 11114 6976 11794 7032
rect 11850 6976 17222 7032
rect 17278 6976 17283 7032
rect 11053 6974 17283 6976
rect 11053 6971 11119 6974
rect 11789 6971 11855 6974
rect 17217 6971 17283 6974
rect 9857 6898 9923 6901
rect 3926 6896 9923 6898
rect 3926 6840 9862 6896
rect 9918 6840 9923 6896
rect 3926 6838 9923 6840
rect 9857 6835 9923 6838
rect 11881 6898 11947 6901
rect 17493 6898 17559 6901
rect 11881 6896 17559 6898
rect 11881 6840 11886 6896
rect 11942 6840 17498 6896
rect 17554 6840 17559 6896
rect 11881 6838 17559 6840
rect 11881 6835 11947 6838
rect 17493 6835 17559 6838
rect 12433 6762 12499 6765
rect 17677 6762 17743 6765
rect 23841 6762 23907 6765
rect 12433 6760 17743 6762
rect 12433 6704 12438 6760
rect 12494 6704 17682 6760
rect 17738 6704 17743 6760
rect 12433 6702 17743 6704
rect 12433 6699 12499 6702
rect 17677 6699 17743 6702
rect 23798 6760 23907 6762
rect 23798 6704 23846 6760
rect 23902 6704 23907 6760
rect 23798 6699 23907 6704
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 13813 6490 13879 6493
rect 14089 6490 14155 6493
rect 13813 6488 14155 6490
rect 13813 6432 13818 6488
rect 13874 6432 14094 6488
rect 14150 6432 14155 6488
rect 13813 6430 14155 6432
rect 13813 6427 13879 6430
rect 14089 6427 14155 6430
rect 16573 6490 16639 6493
rect 20069 6490 20135 6493
rect 16573 6488 20135 6490
rect 16573 6432 16578 6488
rect 16634 6432 20074 6488
rect 20130 6432 20135 6488
rect 16573 6430 20135 6432
rect 16573 6427 16639 6430
rect 20069 6427 20135 6430
rect 23798 6357 23858 6699
rect 24761 6626 24827 6629
rect 27520 6626 28000 6656
rect 24761 6624 28000 6626
rect 24761 6568 24766 6624
rect 24822 6568 28000 6624
rect 24761 6566 28000 6568
rect 24761 6563 24827 6566
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 11697 6354 11763 6357
rect 16297 6354 16363 6357
rect 11697 6352 23674 6354
rect 11697 6296 11702 6352
rect 11758 6296 16302 6352
rect 16358 6296 23674 6352
rect 11697 6294 23674 6296
rect 11697 6291 11763 6294
rect 16297 6291 16363 6294
rect 13445 6218 13511 6221
rect 16757 6218 16823 6221
rect 13445 6216 16823 6218
rect 13445 6160 13450 6216
rect 13506 6160 16762 6216
rect 16818 6160 16823 6216
rect 13445 6158 16823 6160
rect 13445 6155 13511 6158
rect 16757 6155 16823 6158
rect 19241 6218 19307 6221
rect 20713 6218 20779 6221
rect 19241 6216 20779 6218
rect 19241 6160 19246 6216
rect 19302 6160 20718 6216
rect 20774 6160 20779 6216
rect 19241 6158 20779 6160
rect 19241 6155 19307 6158
rect 20713 6155 20779 6158
rect 12065 6082 12131 6085
rect 15745 6082 15811 6085
rect 12065 6080 15811 6082
rect 12065 6024 12070 6080
rect 12126 6024 15750 6080
rect 15806 6024 15811 6080
rect 12065 6022 15811 6024
rect 23614 6082 23674 6294
rect 23749 6352 23858 6357
rect 23749 6296 23754 6352
rect 23810 6296 23858 6352
rect 23749 6294 23858 6296
rect 23749 6291 23815 6294
rect 27520 6082 28000 6112
rect 23614 6022 28000 6082
rect 12065 6019 12131 6022
rect 15745 6019 15811 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 16849 5810 16915 5813
rect 20069 5810 20135 5813
rect 22461 5810 22527 5813
rect 16849 5808 19994 5810
rect 16849 5752 16854 5808
rect 16910 5752 19994 5808
rect 16849 5750 19994 5752
rect 16849 5747 16915 5750
rect 13721 5674 13787 5677
rect 19517 5674 19583 5677
rect 13721 5672 19583 5674
rect 13721 5616 13726 5672
rect 13782 5616 19522 5672
rect 19578 5616 19583 5672
rect 13721 5614 19583 5616
rect 19934 5674 19994 5750
rect 20069 5808 22527 5810
rect 20069 5752 20074 5808
rect 20130 5752 22466 5808
rect 22522 5752 22527 5808
rect 20069 5750 22527 5752
rect 20069 5747 20135 5750
rect 22461 5747 22527 5750
rect 23105 5674 23171 5677
rect 19934 5672 23171 5674
rect 19934 5616 23110 5672
rect 23166 5616 23171 5672
rect 19934 5614 23171 5616
rect 13721 5611 13787 5614
rect 19517 5611 19583 5614
rect 23105 5611 23171 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 18781 5402 18847 5405
rect 23013 5402 23079 5405
rect 27520 5402 28000 5432
rect 18781 5400 23079 5402
rect 18781 5344 18786 5400
rect 18842 5344 23018 5400
rect 23074 5344 23079 5400
rect 18781 5342 23079 5344
rect 18781 5339 18847 5342
rect 23013 5339 23079 5342
rect 24902 5342 28000 5402
rect 21081 5266 21147 5269
rect 24761 5266 24827 5269
rect 21081 5264 24827 5266
rect 21081 5208 21086 5264
rect 21142 5208 24766 5264
rect 24822 5208 24827 5264
rect 21081 5206 24827 5208
rect 21081 5203 21147 5206
rect 24761 5203 24827 5206
rect 17677 5130 17743 5133
rect 18689 5130 18755 5133
rect 24902 5130 24962 5342
rect 27520 5312 28000 5342
rect 17677 5128 24962 5130
rect 17677 5072 17682 5128
rect 17738 5072 18694 5128
rect 18750 5072 24962 5128
rect 17677 5070 24962 5072
rect 17677 5067 17743 5070
rect 18689 5067 18755 5070
rect 10685 4994 10751 4997
rect 14089 4994 14155 4997
rect 10685 4992 14155 4994
rect 10685 4936 10690 4992
rect 10746 4936 14094 4992
rect 14150 4936 14155 4992
rect 10685 4934 14155 4936
rect 10685 4931 10751 4934
rect 14089 4931 14155 4934
rect 14825 4994 14891 4997
rect 17309 4994 17375 4997
rect 14825 4992 17375 4994
rect 14825 4936 14830 4992
rect 14886 4936 17314 4992
rect 17370 4936 17375 4992
rect 14825 4934 17375 4936
rect 14825 4931 14891 4934
rect 17309 4931 17375 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 13261 4858 13327 4861
rect 15837 4858 15903 4861
rect 13261 4856 15903 4858
rect 13261 4800 13266 4856
rect 13322 4800 15842 4856
rect 15898 4800 15903 4856
rect 13261 4798 15903 4800
rect 13261 4795 13327 4798
rect 15837 4795 15903 4798
rect 23013 4858 23079 4861
rect 24853 4858 24919 4861
rect 23013 4856 24919 4858
rect 23013 4800 23018 4856
rect 23074 4800 24858 4856
rect 24914 4800 24919 4856
rect 23013 4798 24919 4800
rect 23013 4795 23079 4798
rect 24853 4795 24919 4798
rect 25313 4858 25379 4861
rect 27520 4858 28000 4888
rect 25313 4856 28000 4858
rect 25313 4800 25318 4856
rect 25374 4800 28000 4856
rect 25313 4798 28000 4800
rect 25313 4795 25379 4798
rect 27520 4768 28000 4798
rect 12801 4722 12867 4725
rect 21081 4722 21147 4725
rect 12801 4720 21147 4722
rect 12801 4664 12806 4720
rect 12862 4664 21086 4720
rect 21142 4664 21147 4720
rect 12801 4662 21147 4664
rect 12801 4659 12867 4662
rect 21081 4659 21147 4662
rect 2957 4586 3023 4589
rect 11789 4586 11855 4589
rect 19701 4586 19767 4589
rect 2957 4584 6194 4586
rect 2957 4528 2962 4584
rect 3018 4528 6194 4584
rect 2957 4526 6194 4528
rect 2957 4523 3023 4526
rect 6134 4450 6194 4526
rect 11789 4584 19767 4586
rect 11789 4528 11794 4584
rect 11850 4528 19706 4584
rect 19762 4528 19767 4584
rect 11789 4526 19767 4528
rect 11789 4523 11855 4526
rect 19701 4523 19767 4526
rect 14733 4450 14799 4453
rect 6134 4448 14799 4450
rect 6134 4392 14738 4448
rect 14794 4392 14799 4448
rect 6134 4390 14799 4392
rect 14733 4387 14799 4390
rect 15510 4388 15516 4452
rect 15580 4450 15586 4452
rect 24117 4450 24183 4453
rect 15580 4448 24183 4450
rect 15580 4392 24122 4448
rect 24178 4392 24183 4448
rect 15580 4390 24183 4392
rect 15580 4388 15586 4390
rect 24117 4387 24183 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 26049 4314 26115 4317
rect 27520 4314 28000 4344
rect 26049 4312 28000 4314
rect 26049 4256 26054 4312
rect 26110 4256 28000 4312
rect 26049 4254 28000 4256
rect 26049 4251 26115 4254
rect 27520 4224 28000 4254
rect 933 4178 999 4181
rect 22645 4178 22711 4181
rect 24117 4178 24183 4181
rect 933 4176 15026 4178
rect 933 4120 938 4176
rect 994 4120 15026 4176
rect 933 4118 15026 4120
rect 933 4115 999 4118
rect 7097 4042 7163 4045
rect 10041 4042 10107 4045
rect 7097 4040 10107 4042
rect 7097 3984 7102 4040
rect 7158 3984 10046 4040
rect 10102 3984 10107 4040
rect 7097 3982 10107 3984
rect 14966 4042 15026 4118
rect 22645 4176 24183 4178
rect 22645 4120 22650 4176
rect 22706 4120 24122 4176
rect 24178 4120 24183 4176
rect 22645 4118 24183 4120
rect 22645 4115 22711 4118
rect 24117 4115 24183 4118
rect 21817 4042 21883 4045
rect 14966 4040 21883 4042
rect 14966 3984 21822 4040
rect 21878 3984 21883 4040
rect 14966 3982 21883 3984
rect 7097 3979 7163 3982
rect 10041 3979 10107 3982
rect 21817 3979 21883 3982
rect 22001 4042 22067 4045
rect 25313 4042 25379 4045
rect 22001 4040 25379 4042
rect 22001 3984 22006 4040
rect 22062 3984 25318 4040
rect 25374 3984 25379 4040
rect 22001 3982 25379 3984
rect 22001 3979 22067 3982
rect 25313 3979 25379 3982
rect 11881 3906 11947 3909
rect 15561 3906 15627 3909
rect 11881 3904 15627 3906
rect 11881 3848 11886 3904
rect 11942 3848 15566 3904
rect 15622 3848 15627 3904
rect 11881 3846 15627 3848
rect 11881 3843 11947 3846
rect 15561 3843 15627 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 11421 3770 11487 3773
rect 15285 3770 15351 3773
rect 11421 3768 15351 3770
rect 11421 3712 11426 3768
rect 11482 3712 15290 3768
rect 15346 3712 15351 3768
rect 11421 3710 15351 3712
rect 11421 3707 11487 3710
rect 15285 3707 15351 3710
rect 15469 3770 15535 3773
rect 17953 3770 18019 3773
rect 15469 3768 18019 3770
rect 15469 3712 15474 3768
rect 15530 3712 17958 3768
rect 18014 3712 18019 3768
rect 15469 3710 18019 3712
rect 15469 3707 15535 3710
rect 17953 3707 18019 3710
rect 22553 3770 22619 3773
rect 27520 3770 28000 3800
rect 22553 3768 28000 3770
rect 22553 3712 22558 3768
rect 22614 3712 28000 3768
rect 22553 3710 28000 3712
rect 22553 3707 22619 3710
rect 27520 3680 28000 3710
rect 4337 3634 4403 3637
rect 11973 3634 12039 3637
rect 4337 3632 12039 3634
rect 4337 3576 4342 3632
rect 4398 3576 11978 3632
rect 12034 3576 12039 3632
rect 4337 3574 12039 3576
rect 4337 3571 4403 3574
rect 11973 3571 12039 3574
rect 14733 3634 14799 3637
rect 19609 3634 19675 3637
rect 14733 3632 19675 3634
rect 14733 3576 14738 3632
rect 14794 3576 19614 3632
rect 19670 3576 19675 3632
rect 14733 3574 19675 3576
rect 14733 3571 14799 3574
rect 19609 3571 19675 3574
rect 11421 3498 11487 3501
rect 18045 3498 18111 3501
rect 11421 3496 18111 3498
rect 11421 3440 11426 3496
rect 11482 3440 18050 3496
rect 18106 3440 18111 3496
rect 11421 3438 18111 3440
rect 11421 3435 11487 3438
rect 18045 3435 18111 3438
rect 18505 3498 18571 3501
rect 20437 3498 20503 3501
rect 18505 3496 20503 3498
rect 18505 3440 18510 3496
rect 18566 3440 20442 3496
rect 20498 3440 20503 3496
rect 18505 3438 20503 3440
rect 18505 3435 18571 3438
rect 20437 3435 20503 3438
rect 8385 3362 8451 3365
rect 13077 3362 13143 3365
rect 8385 3360 13143 3362
rect 8385 3304 8390 3360
rect 8446 3304 13082 3360
rect 13138 3304 13143 3360
rect 8385 3302 13143 3304
rect 8385 3299 8451 3302
rect 13077 3299 13143 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 11881 3226 11947 3229
rect 15561 3228 15627 3229
rect 11881 3224 14842 3226
rect 11881 3168 11886 3224
rect 11942 3168 14842 3224
rect 11881 3166 14842 3168
rect 11881 3163 11947 3166
rect 6361 3090 6427 3093
rect 13353 3090 13419 3093
rect 6361 3088 13419 3090
rect 6361 3032 6366 3088
rect 6422 3032 13358 3088
rect 13414 3032 13419 3088
rect 6361 3030 13419 3032
rect 14782 3090 14842 3166
rect 15510 3164 15516 3228
rect 15580 3226 15627 3228
rect 27520 3226 28000 3256
rect 15580 3224 15672 3226
rect 15622 3168 15672 3224
rect 15580 3166 15672 3168
rect 24902 3166 28000 3226
rect 15580 3164 15627 3166
rect 15561 3163 15627 3164
rect 15745 3090 15811 3093
rect 14782 3088 15811 3090
rect 14782 3032 15750 3088
rect 15806 3032 15811 3088
rect 14782 3030 15811 3032
rect 6361 3027 6427 3030
rect 13353 3027 13419 3030
rect 15745 3027 15811 3030
rect 18137 3090 18203 3093
rect 21541 3090 21607 3093
rect 18137 3088 21607 3090
rect 18137 3032 18142 3088
rect 18198 3032 21546 3088
rect 21602 3032 21607 3088
rect 18137 3030 21607 3032
rect 18137 3027 18203 3030
rect 21541 3027 21607 3030
rect 21909 3090 21975 3093
rect 24902 3090 24962 3166
rect 27520 3136 28000 3166
rect 21909 3088 24962 3090
rect 21909 3032 21914 3088
rect 21970 3032 24962 3088
rect 21909 3030 24962 3032
rect 21909 3027 21975 3030
rect 11421 2954 11487 2957
rect 20345 2954 20411 2957
rect 23790 2954 23796 2956
rect 11421 2952 17050 2954
rect 11421 2896 11426 2952
rect 11482 2896 17050 2952
rect 11421 2894 17050 2896
rect 11421 2891 11487 2894
rect 10961 2818 11027 2821
rect 16849 2818 16915 2821
rect 10961 2816 16915 2818
rect 10961 2760 10966 2816
rect 11022 2760 16854 2816
rect 16910 2760 16915 2816
rect 10961 2758 16915 2760
rect 16990 2818 17050 2894
rect 20345 2952 23796 2954
rect 20345 2896 20350 2952
rect 20406 2896 23796 2952
rect 20345 2894 23796 2896
rect 20345 2891 20411 2894
rect 23790 2892 23796 2894
rect 23860 2954 23866 2956
rect 24577 2954 24643 2957
rect 23860 2952 24643 2954
rect 23860 2896 24582 2952
rect 24638 2896 24643 2952
rect 23860 2894 24643 2896
rect 23860 2892 23866 2894
rect 24577 2891 24643 2894
rect 19333 2818 19399 2821
rect 16990 2816 19399 2818
rect 16990 2760 19338 2816
rect 19394 2760 19399 2816
rect 16990 2758 19399 2760
rect 10961 2755 11027 2758
rect 16849 2755 16915 2758
rect 19333 2755 19399 2758
rect 20069 2818 20135 2821
rect 23473 2818 23539 2821
rect 20069 2816 23539 2818
rect 20069 2760 20074 2816
rect 20130 2760 23478 2816
rect 23534 2760 23539 2816
rect 20069 2758 23539 2760
rect 20069 2755 20135 2758
rect 23473 2755 23539 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 10869 2682 10935 2685
rect 16665 2682 16731 2685
rect 10869 2680 16731 2682
rect 10869 2624 10874 2680
rect 10930 2624 16670 2680
rect 16726 2624 16731 2680
rect 10869 2622 16731 2624
rect 10869 2619 10935 2622
rect 16665 2619 16731 2622
rect 1577 2546 1643 2549
rect 20897 2546 20963 2549
rect 1577 2544 20963 2546
rect 1577 2488 1582 2544
rect 1638 2488 20902 2544
rect 20958 2488 20963 2544
rect 1577 2486 20963 2488
rect 1577 2483 1643 2486
rect 20897 2483 20963 2486
rect 24577 2546 24643 2549
rect 27520 2546 28000 2576
rect 24577 2544 28000 2546
rect 24577 2488 24582 2544
rect 24638 2488 28000 2544
rect 24577 2486 28000 2488
rect 24577 2483 24643 2486
rect 27520 2456 28000 2486
rect 12893 2410 12959 2413
rect 22093 2410 22159 2413
rect 12893 2408 22159 2410
rect 12893 2352 12898 2408
rect 12954 2352 22098 2408
rect 22154 2352 22159 2408
rect 12893 2350 22159 2352
rect 12893 2347 12959 2350
rect 22093 2347 22159 2350
rect 16665 2274 16731 2277
rect 23974 2274 23980 2276
rect 16665 2272 23980 2274
rect 16665 2216 16670 2272
rect 16726 2216 23980 2272
rect 16665 2214 23980 2216
rect 16665 2211 16731 2214
rect 23974 2212 23980 2214
rect 24044 2212 24050 2276
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 11605 2002 11671 2005
rect 20713 2002 20779 2005
rect 27520 2002 28000 2032
rect 11605 2000 20779 2002
rect 11605 1944 11610 2000
rect 11666 1944 20718 2000
rect 20774 1944 20779 2000
rect 11605 1942 20779 1944
rect 11605 1939 11671 1942
rect 20713 1939 20779 1942
rect 26926 1942 28000 2002
rect 5717 1866 5783 1869
rect 13629 1866 13695 1869
rect 5717 1864 13695 1866
rect 5717 1808 5722 1864
rect 5778 1808 13634 1864
rect 13690 1808 13695 1864
rect 5717 1806 13695 1808
rect 5717 1803 5783 1806
rect 13629 1803 13695 1806
rect 17401 1866 17467 1869
rect 26926 1866 26986 1942
rect 27520 1912 28000 1942
rect 17401 1864 26986 1866
rect 17401 1808 17406 1864
rect 17462 1808 26986 1864
rect 17401 1806 26986 1808
rect 17401 1803 17467 1806
rect 9213 1730 9279 1733
rect 18873 1730 18939 1733
rect 9213 1728 18939 1730
rect 9213 1672 9218 1728
rect 9274 1672 18878 1728
rect 18934 1672 18939 1728
rect 9213 1670 18939 1672
rect 9213 1667 9279 1670
rect 18873 1667 18939 1670
rect 8753 1594 8819 1597
rect 14549 1594 14615 1597
rect 8753 1592 14615 1594
rect 8753 1536 8758 1592
rect 8814 1536 14554 1592
rect 14610 1536 14615 1592
rect 8753 1534 14615 1536
rect 8753 1531 8819 1534
rect 14549 1531 14615 1534
rect 15745 1594 15811 1597
rect 21357 1594 21423 1597
rect 15745 1592 21423 1594
rect 15745 1536 15750 1592
rect 15806 1536 21362 1592
rect 21418 1536 21423 1592
rect 15745 1534 21423 1536
rect 15745 1531 15811 1534
rect 21357 1531 21423 1534
rect 10501 1458 10567 1461
rect 18689 1458 18755 1461
rect 10501 1456 18755 1458
rect 10501 1400 10506 1456
rect 10562 1400 18694 1456
rect 18750 1400 18755 1456
rect 10501 1398 18755 1400
rect 10501 1395 10567 1398
rect 18689 1395 18755 1398
rect 23749 1458 23815 1461
rect 27520 1458 28000 1488
rect 23749 1456 28000 1458
rect 23749 1400 23754 1456
rect 23810 1400 28000 1456
rect 23749 1398 28000 1400
rect 23749 1395 23815 1398
rect 27520 1368 28000 1398
rect 18965 914 19031 917
rect 27520 914 28000 944
rect 18965 912 28000 914
rect 18965 856 18970 912
rect 19026 856 28000 912
rect 18965 854 28000 856
rect 18965 851 19031 854
rect 27520 824 28000 854
rect 23657 370 23723 373
rect 27520 370 28000 400
rect 23657 368 28000 370
rect 23657 312 23662 368
rect 23718 312 28000 368
rect 23657 310 28000 312
rect 23657 307 23723 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 14228 22612 14292 22676
rect 23980 22340 24044 22404
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 14228 19348 14292 19412
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 23796 11928 23860 11932
rect 23796 11872 23846 11928
rect 23846 11872 23860 11928
rect 23796 11868 23860 11872
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 15516 9480 15580 9484
rect 15516 9424 15566 9480
rect 15566 9424 15580 9480
rect 15516 9420 15580 9424
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 15516 4388 15580 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 15516 3224 15580 3228
rect 15516 3168 15566 3224
rect 15566 3168 15580 3224
rect 15516 3164 15580 3168
rect 23796 2892 23860 2956
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 23980 2212 24044 2276
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14227 22676 14293 22677
rect 14227 22612 14228 22676
rect 14292 22612 14293 22676
rect 14227 22611 14293 22612
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 14230 19413 14290 22611
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14227 19412 14293 19413
rect 14227 19348 14228 19412
rect 14292 19348 14293 19412
rect 14227 19347 14293 19348
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 23979 22404 24045 22405
rect 23979 22340 23980 22404
rect 24044 22340 24045 22404
rect 23979 22339 24045 22340
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 23795 11932 23861 11933
rect 23795 11868 23796 11932
rect 23860 11868 23861 11932
rect 23795 11867 23861 11868
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 15515 9484 15581 9485
rect 15515 9420 15516 9484
rect 15580 9420 15581 9484
rect 15515 9419 15581 9420
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 15518 4453 15578 9419
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 15515 4452 15581 4453
rect 15515 4388 15516 4452
rect 15580 4388 15581 4452
rect 15515 4387 15581 4388
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 15518 3229 15578 4387
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 15515 3228 15581 3229
rect 15515 3164 15516 3228
rect 15580 3164 15581 3228
rect 15515 3163 15581 3164
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 23798 2957 23858 11867
rect 23795 2956 23861 2957
rect 23795 2892 23796 2956
rect 23860 2892 23861 2956
rect 23795 2891 23861 2892
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 23982 2277 24042 22339
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 23979 2276 24045 2277
rect 23979 2212 23980 2276
rect 24044 2212 24045 2276
rect 23979 2211 24045 2212
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_128
timestamp 1604681595
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_130
timestamp 1604681595
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 12696 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_152
timestamp 1604681595
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1604681595
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 15548 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_176
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_180
timestamp 1604681595
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18124 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_201
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_205
timestamp 1604681595
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1604681595
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_227
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21436 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_1_235
timestamp 1604681595
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_231
timestamp 1604681595
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_234
timestamp 1604681595
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_238
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_246
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_255
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_251
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_255
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_267
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_263
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_267
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 24932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_275
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _039_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_102
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12328 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_114
timestamp 1604681595
transform 1 0 11592 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1604681595
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1604681595
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1604681595
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_164
timestamp 1604681595
transform 1 0 16192 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16560 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_184
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_192
timestamp 1604681595
transform 1 0 18768 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21712 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_223
timestamp 1604681595
transform 1 0 21620 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23920 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1604681595
transform 1 0 23184 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_244
timestamp 1604681595
transform 1 0 23552 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_257
timestamp 1604681595
transform 1 0 24748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_261
timestamp 1604681595
transform 1 0 25116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_265
timestamp 1604681595
transform 1 0 25484 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_273
timestamp 1604681595
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1604681595
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1604681595
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_145
timestamp 1604681595
transform 1 0 14444 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15640 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1604681595
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1604681595
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_174
timestamp 1604681595
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1604681595
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1604681595
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18584 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1604681595
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1604681595
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_223
timestamp 1604681595
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1604681595
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_254
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1604681595
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_266
timestamp 1604681595
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_270
timestamp 1604681595
transform 1 0 25944 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 11776 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_113
timestamp 1604681595
transform 1 0 11500 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_119
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 12788 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_131
timestamp 1604681595
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_135
timestamp 1604681595
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17296 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_170
timestamp 1604681595
transform 1 0 16744 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_185
timestamp 1604681595
transform 1 0 18124 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18860 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_207
timestamp 1604681595
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1604681595
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1604681595
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_225
timestamp 1604681595
transform 1 0 21804 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_229
timestamp 1604681595
transform 1 0 22172 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 22448 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_248
timestamp 1604681595
transform 1 0 23920 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_252
timestamp 1604681595
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_265
timestamp 1604681595
transform 1 0 25484 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_273
timestamp 1604681595
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 13064 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1604681595
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_151
timestamp 1604681595
transform 1 0 14996 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_180
timestamp 1604681595
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19964 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18400 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_201
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1604681595
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1604681595
transform 1 0 21804 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_229
timestamp 1604681595
transform 1 0 22172 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_261
timestamp 1604681595
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_265
timestamp 1604681595
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1604681595
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_100
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_104
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1604681595
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604681595
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_122
timestamp 1604681595
transform 1 0 12328 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 12052 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 1604681595
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_129
timestamp 1604681595
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_133
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 13064 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_139
timestamp 1604681595
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13708 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15916 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_174
timestamp 1604681595
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_170
timestamp 1604681595
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_175
timestamp 1604681595
transform 1 0 17204 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_170
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1604681595
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1604681595
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18676 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_194
timestamp 1604681595
transform 1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_199
timestamp 1604681595
transform 1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_188
timestamp 1604681595
transform 1 0 18400 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_207
timestamp 1604681595
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_211
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 20976 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1604681595
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_228
timestamp 1604681595
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604681595
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_236
timestamp 1604681595
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 22448 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_240
timestamp 1604681595
transform 1 0 23184 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23368 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23552 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_250
timestamp 1604681595
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_257
timestamp 1604681595
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1604681595
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24288 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24472 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_267
timestamp 1604681595
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_263
timestamp 1604681595
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1604681595
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 25116 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1604681595
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_275
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9752 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_110
timestamp 1604681595
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_114
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_132
timestamp 1604681595
transform 1 0 13248 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_169
timestamp 1604681595
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_176
timestamp 1604681595
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_189
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_194
timestamp 1604681595
transform 1 0 18952 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21252 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_210
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23828 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_235
timestamp 1604681595
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_243
timestamp 1604681595
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 25392 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_256
timestamp 1604681595
transform 1 0 24656 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_267
timestamp 1604681595
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1604681595
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1604681595
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_168
timestamp 1604681595
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_173
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_177
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18768 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_205
timestamp 1604681595
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20516 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1604681595
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_224
timestamp 1604681595
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_228
timestamp 1604681595
transform 1 0 22080 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 22356 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_235
timestamp 1604681595
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_239
timestamp 1604681595
transform 1 0 23092 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_261
timestamp 1604681595
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1604681595
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 1604681595
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1604681595
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_138
timestamp 1604681595
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_167
timestamp 1604681595
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1604681595
transform 1 0 17664 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_194
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_206
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_210
timestamp 1604681595
transform 1 0 20424 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_224
timestamp 1604681595
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_228
timestamp 1604681595
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 22540 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23644 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_232
timestamp 1604681595
transform 1 0 22448 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_236
timestamp 1604681595
transform 1 0 22816 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_242
timestamp 1604681595
transform 1 0 23368 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_261
timestamp 1604681595
transform 1 0 25116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_273
timestamp 1604681595
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_94
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_136
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1604681595
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14536 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_162
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1604681595
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1604681595
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_204
timestamp 1604681595
transform 1 0 19872 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20700 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 20332 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_212
timestamp 1604681595
transform 1 0 20608 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_229
timestamp 1604681595
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_233
timestamp 1604681595
transform 1 0 22540 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_237
timestamp 1604681595
transform 1 0 22908 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_249
timestamp 1604681595
transform 1 0 24012 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24104 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24288 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_261
timestamp 1604681595
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_265
timestamp 1604681595
transform 1 0 25484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_101
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11776 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1604681595
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1604681595
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_132
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_136
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1604681595
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_180
timestamp 1604681595
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_184
timestamp 1604681595
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_188
timestamp 1604681595
transform 1 0 18400 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23736 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22540 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23552 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_231
timestamp 1604681595
transform 1 0 22356 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_235
timestamp 1604681595
transform 1 0 22724 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_243
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_262
timestamp 1604681595
transform 1 0 25208 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_97
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1604681595
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_14_118
timestamp 1604681595
transform 1 0 11960 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_130
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1604681595
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12696 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_150
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_154
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1604681595
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1604681595
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_173
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1604681595
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17112 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1604681595
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1604681595
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1604681595
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_205
timestamp 1604681595
transform 1 0 19964 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19596 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1604681595
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20332 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604681595
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604681595
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1604681595
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21804 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_238
timestamp 1604681595
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_232
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_234
timestamp 1604681595
transform 1 0 22632 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 22724 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_242
timestamp 1604681595
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 23552 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23828 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23736 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_256
timestamp 1604681595
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_260
timestamp 1604681595
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_267
timestamp 1604681595
transform 1 0 25668 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_262
timestamp 1604681595
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_266
timestamp 1604681595
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_275
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604681595
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1604681595
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_160
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_204
timestamp 1604681595
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_211
timestamp 1604681595
transform 1 0 20516 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1604681595
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23736 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_255
timestamp 1604681595
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1604681595
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_270
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_274
timestamp 1604681595
transform 1 0 26312 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_121
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13524 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_126
timestamp 1604681595
transform 1 0 12696 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_144
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_167
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_171
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_175
timestamp 1604681595
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_192
timestamp 1604681595
transform 1 0 18768 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20976 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1604681595
transform 1 0 21804 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_229
timestamp 1604681595
transform 1 0 22172 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 22724 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22356 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_233
timestamp 1604681595
transform 1 0 22540 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 24932 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 24748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_255
timestamp 1604681595
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_104
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604681595
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12512 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_130
timestamp 1604681595
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_134
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16008 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_154
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1604681595
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_197
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_201
timestamp 1604681595
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_205
timestamp 1604681595
transform 1 0 19964 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20424 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_219
timestamp 1604681595
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_223
timestamp 1604681595
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1604681595
transform 1 0 24012 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24288 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_261
timestamp 1604681595
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_265
timestamp 1604681595
transform 1 0 25484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1604681595
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_194
timestamp 1604681595
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22540 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22908 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1604681595
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_235
timestamp 1604681595
transform 1 0 22724 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_242
timestamp 1604681595
transform 1 0 23368 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_247
timestamp 1604681595
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_101
timestamp 1604681595
transform 1 0 10396 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 10120 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_107
timestamp 1604681595
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11132 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1604681595
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_165
timestamp 1604681595
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_169
timestamp 1604681595
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1604681595
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18308 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17020 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18860 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19872 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1604681595
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_209
timestamp 1604681595
transform 1 0 20332 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1604681595
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_225
timestamp 1604681595
transform 1 0 21804 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_224
timestamp 1604681595
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21620 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_229
timestamp 1604681595
transform 1 0 22172 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_238
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_234
timestamp 1604681595
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22264 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_243
timestamp 1604681595
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23276 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1604681595
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_265
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9476 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 12604 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_128
timestamp 1604681595
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1604681595
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15180 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1604681595
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_204
timestamp 1604681595
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24564 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_251
timestamp 1604681595
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1604681595
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_268
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_99
timestamp 1604681595
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_103
timestamp 1604681595
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_123
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_127
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_160
timestamp 1604681595
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_164
timestamp 1604681595
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1604681595
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_186
timestamp 1604681595
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_194
timestamp 1604681595
transform 1 0 18952 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_224
timestamp 1604681595
transform 1 0 21712 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_229
timestamp 1604681595
transform 1 0 22172 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_241
timestamp 1604681595
transform 1 0 23276 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1604681595
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_258
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_262
timestamp 1604681595
transform 1 0 25208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 1604681595
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604681595
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12604 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14168 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_134
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1604681595
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1604681595
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19872 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_199
timestamp 1604681595
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_203
timestamp 1604681595
transform 1 0 19780 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_224
timestamp 1604681595
transform 1 0 21712 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 24104 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1604681595
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_270
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_274
timestamp 1604681595
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1604681595
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1604681595
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1604681595
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_137
timestamp 1604681595
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_148
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1604681595
transform 1 0 15916 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_165
timestamp 1604681595
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16652 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1604681595
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21068 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22172 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21804 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_223
timestamp 1604681595
transform 1 0 21620 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 22356 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_247
timestamp 1604681595
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24564 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_264
timestamp 1604681595
transform 1 0 25392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_268
timestamp 1604681595
transform 1 0 25760 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604681595
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_108
timestamp 1604681595
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1604681595
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_116
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_156
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_168
timestamp 1604681595
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1604681595
transform 1 0 16928 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_176
timestamp 1604681595
transform 1 0 17296 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20056 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1604681595
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1604681595
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21896 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_224
timestamp 1604681595
transform 1 0 21712 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_228
timestamp 1604681595
transform 1 0 22080 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 25576 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_262
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10856 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1604681595
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_139
timestamp 1604681595
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1604681595
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_150
timestamp 1604681595
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_147
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15548 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_27_173
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_174
timestamp 1604681595
transform 1 0 17112 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1604681595
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16928 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17664 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17848 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18124 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_194
timestamp 1604681595
transform 1 0 18952 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_199
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_199
timestamp 1604681595
transform 1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19688 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1604681595
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20976 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1604681595
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1604681595
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_229
timestamp 1604681595
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1604681595
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22632 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 22540 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_244
timestamp 1604681595
transform 1 0 23552 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_240
timestamp 1604681595
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23736 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23920 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_257
timestamp 1604681595
transform 1 0 24748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_261
timestamp 1604681595
transform 1 0 25116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_261
timestamp 1604681595
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1604681595
transform 1 0 25484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_273
timestamp 1604681595
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11684 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp 1604681595
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1604681595
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_142
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_148
timestamp 1604681595
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_160
timestamp 1604681595
transform 1 0 15824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_165
timestamp 1604681595
transform 1 0 16284 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16560 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_184
timestamp 1604681595
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 18952 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_188
timestamp 1604681595
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604681595
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_224
timestamp 1604681595
transform 1 0 21712 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_229
timestamp 1604681595
transform 1 0 22172 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 22908 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 22448 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_234
timestamp 1604681595
transform 1 0 22632 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 25116 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1604681595
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_257
timestamp 1604681595
transform 1 0 24748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1604681595
transform 1 0 25484 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 1604681595
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12788 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_140
timestamp 1604681595
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14996 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_148
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_160
timestamp 1604681595
transform 1 0 15824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 18216 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_174
timestamp 1604681595
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_178
timestamp 1604681595
transform 1 0 17480 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1604681595
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1604681595
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20792 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1604681595
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_223
timestamp 1604681595
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_227
timestamp 1604681595
transform 1 0 21988 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_254
timestamp 1604681595
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1604681595
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_266
timestamp 1604681595
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_270
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11408 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_111
timestamp 1604681595
transform 1 0 11316 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1604681595
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1604681595
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1604681595
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 14536 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_159
timestamp 1604681595
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17112 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1604681595
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1604681595
transform 1 0 17296 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_180
timestamp 1604681595
transform 1 0 17664 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1604681595
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_187
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18400 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_204
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 21160 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_222
timestamp 1604681595
transform 1 0 21528 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_226
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_229
timestamp 1604681595
transform 1 0 22172 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 22264 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23920 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_246
timestamp 1604681595
transform 1 0 23736 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1604681595
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24472 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_267
timestamp 1604681595
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_100
timestamp 1604681595
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_104
timestamp 1604681595
transform 1 0 10672 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1604681595
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_143
timestamp 1604681595
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1604681595
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_187
timestamp 1604681595
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_191
timestamp 1604681595
transform 1 0 18676 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1604681595
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_224
timestamp 1604681595
transform 1 0 21712 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1604681595
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_268
timestamp 1604681595
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_272
timestamp 1604681595
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_276
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1604681595
transform 1 0 11592 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_120
timestamp 1604681595
transform 1 0 12144 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_124
timestamp 1604681595
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_144
timestamp 1604681595
transform 1 0 14352 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15548 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1604681595
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1604681595
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_198
timestamp 1604681595
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 21160 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_210
timestamp 1604681595
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1604681595
transform 1 0 21528 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_226
timestamp 1604681595
transform 1 0 21896 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_229
timestamp 1604681595
transform 1 0 22172 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 22264 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23920 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_246
timestamp 1604681595
transform 1 0 23736 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1604681595
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24472 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1604681595
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_101
timestamp 1604681595
transform 1 0 10396 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_97
timestamp 1604681595
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10488 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_122
timestamp 1604681595
transform 1 0 12328 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1604681595
transform 1 0 11960 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_135
timestamp 1604681595
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_134
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_130
timestamp 1604681595
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_126
timestamp 1604681595
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_139
timestamp 1604681595
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 14260 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_150
timestamp 1604681595
transform 1 0 14904 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_146
timestamp 1604681595
transform 1 0 14536 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1604681595
transform 1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14720 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_158
timestamp 1604681595
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15640 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15824 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1604681595
transform 1 0 17296 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_182
timestamp 1604681595
transform 1 0 17848 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18032 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_193
timestamp 1604681595
transform 1 0 18860 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1604681595
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1604681595
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19228 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1604681595
transform 1 0 20056 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_199
timestamp 1604681595
transform 1 0 19412 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_216
timestamp 1604681595
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_212
timestamp 1604681595
transform 1 0 20608 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21068 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_219
timestamp 1604681595
transform 1 0 21252 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_223
timestamp 1604681595
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21804 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21436 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_237
timestamp 1604681595
transform 1 0 22908 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_241
timestamp 1604681595
transform 1 0 23276 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_254
timestamp 1604681595
transform 1 0 24472 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_266
timestamp 1604681595
transform 1 0 25576 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 25208 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_268
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_108
timestamp 1604681595
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_112
timestamp 1604681595
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14168 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_132
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_138
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_151
timestamp 1604681595
transform 1 0 14996 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1604681595
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1604681595
transform 1 0 17020 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_200
timestamp 1604681595
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1604681595
transform 1 0 19872 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20424 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1604681595
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_223
timestamp 1604681595
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1604681595
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 25484 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24196 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_263
timestamp 1604681595
transform 1 0 25300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 26036 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_101
timestamp 1604681595
transform 1 0 10396 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10948 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_123
timestamp 1604681595
transform 1 0 12420 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_131
timestamp 1604681595
transform 1 0 13156 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15640 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_167
timestamp 1604681595
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_171
timestamp 1604681595
transform 1 0 16836 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1604681595
transform 1 0 17388 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18676 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19044 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_189
timestamp 1604681595
transform 1 0 18492 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_193
timestamp 1604681595
transform 1 0 18860 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_206
timestamp 1604681595
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21068 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_210
timestamp 1604681595
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23828 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22724 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_233
timestamp 1604681595
transform 1 0 22540 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_237
timestamp 1604681595
transform 1 0 22908 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_245
timestamp 1604681595
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25116 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1604681595
transform 1 0 24380 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_267
timestamp 1604681595
transform 1 0 25668 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14444 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_139
timestamp 1604681595
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_143
timestamp 1604681595
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_156
timestamp 1604681595
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_160
timestamp 1604681595
transform 1 0 15824 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_181
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18952 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18768 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_188
timestamp 1604681595
transform 1 0 18400 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21160 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_210
timestamp 1604681595
transform 1 0 20424 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_214
timestamp 1604681595
transform 1 0 20792 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_217
timestamp 1604681595
transform 1 0 21068 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_234
timestamp 1604681595
transform 1 0 22632 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 24932 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 25484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_251
timestamp 1604681595
transform 1 0 24196 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_255
timestamp 1604681595
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_263
timestamp 1604681595
transform 1 0 25300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_267
timestamp 1604681595
transform 1 0 25668 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_275
timestamp 1604681595
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 11960 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_121
timestamp 1604681595
transform 1 0 12236 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_125
timestamp 1604681595
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1604681595
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17572 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16928 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17296 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_170
timestamp 1604681595
transform 1 0 16744 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_174
timestamp 1604681595
transform 1 0 17112 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 19780 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 19596 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_195
timestamp 1604681595
transform 1 0 19044 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_199
timestamp 1604681595
transform 1 0 19412 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_206
timestamp 1604681595
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_210
timestamp 1604681595
transform 1 0 20424 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_224
timestamp 1604681595
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_228
timestamp 1604681595
transform 1 0 22080 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 22540 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 22356 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_237
timestamp 1604681595
transform 1 0 22908 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24932 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_265
timestamp 1604681595
transform 1 0 25484 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_273
timestamp 1604681595
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_132
timestamp 1604681595
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604681595
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_142
timestamp 1604681595
transform 1 0 14168 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_137
timestamp 1604681595
transform 1 0 13708 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_136
timestamp 1604681595
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604681595
transform 1 0 14352 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 13800 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 13984 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_40_150
timestamp 1604681595
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_146
timestamp 1604681595
transform 1 0 14536 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_162
timestamp 1604681595
transform 1 0 16008 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_158
timestamp 1604681595
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_160
timestamp 1604681595
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_156
timestamp 1604681595
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604681595
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_173
timestamp 1604681595
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_187
timestamp 1604681595
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_183
timestamp 1604681595
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18124 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16468 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_40_195
timestamp 1604681595
transform 1 0 19044 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1604681595
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18492 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604681595
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 18676 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_200
timestamp 1604681595
transform 1 0 19504 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_205
timestamp 1604681595
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_197
timestamp 1604681595
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 19320 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 19596 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 19780 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_206
timestamp 1604681595
transform 1 0 20056 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_217
timestamp 1604681595
transform 1 0 21068 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_209
timestamp 1604681595
transform 1 0 20332 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1604681595
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_235
timestamp 1604681595
transform 1 0 22724 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_247
timestamp 1604681595
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 25484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1604681595
transform 1 0 24196 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_263
timestamp 1604681595
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_267
timestamp 1604681595
transform 1 0 25668 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_259
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1604681595
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 14260 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_131
timestamp 1604681595
transform 1 0 13156 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1604681595
transform 1 0 13892 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_145
timestamp 1604681595
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 15916 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15364 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_153
timestamp 1604681595
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_157
timestamp 1604681595
transform 1 0 15548 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_165
timestamp 1604681595
transform 1 0 16284 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604681595
transform 1 0 16468 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1604681595
transform 1 0 16652 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_173
timestamp 1604681595
transform 1 0 17020 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 19320 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 19964 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_188
timestamp 1604681595
transform 1 0 18400 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_192
timestamp 1604681595
transform 1 0 18768 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_195
timestamp 1604681595
transform 1 0 19044 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_202
timestamp 1604681595
transform 1 0 19688 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_207
timestamp 1604681595
transform 1 0 20148 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 21528 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 20424 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 22080 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 20976 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_214
timestamp 1604681595
transform 1 0 20792 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_218
timestamp 1604681595
transform 1 0 21160 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_226
timestamp 1604681595
transform 1 0 21896 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_230
timestamp 1604681595
transform 1 0 22264 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_234
timestamp 1604681595
transform 1 0 22632 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_242
timestamp 1604681595
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_259
timestamp 1604681595
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_275
timestamp 1604681595
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_147
timestamp 1604681595
transform 1 0 14628 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_159
timestamp 1604681595
transform 1 0 15732 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 16468 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_171
timestamp 1604681595
transform 1 0 16836 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_183
timestamp 1604681595
transform 1 0 17940 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 18860 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1604681595
transform 1 0 19228 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 21896 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1604681595
transform 1 0 20332 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 6944 480 7064 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 20952 480 21072 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27520 23672 28000 23792 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26882 0 26938 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 938 27520 994 28000 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 7746 27520 7802 28000 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 9126 27520 9182 28000 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1582 27520 1638 28000 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2962 27520 3018 28000 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4986 27520 5042 28000 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 5722 27520 5778 28000 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 23478 27520 23534 28000 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 25502 27520 25558 28000 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 26146 27520 26202 28000 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 26882 27520 26938 28000 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 27526 27520 27582 28000 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 15290 27520 15346 28000 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 17314 27520 17370 28000 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 20718 27520 20774 28000 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 prog_clk
port 123 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 124 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 125 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 126 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 127 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_bottom_grid_pin_38_
port 128 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 129 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 130 nsew default input
rlabel metal3 s 27520 4224 28000 4344 6 right_bottom_grid_pin_41_
port 131 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
