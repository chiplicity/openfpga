magic
tech sky130A
magscale 1 2
timestamp 1605014388
<< locali >>
rect 4445 29087 4479 29257
rect 11621 27455 11655 27625
rect 6837 25347 6871 25449
rect 6009 24667 6043 24837
rect 6377 24803 6411 24905
rect 13277 24599 13311 24837
rect 3709 16643 3743 16745
rect 8585 14875 8619 15113
rect 3617 13243 3651 13345
rect 12081 3927 12115 4233
rect 8125 2975 8159 3077
<< viali >>
rect 11785 36193 11819 36227
rect 11529 36125 11563 36159
rect 12909 35989 12943 36023
rect 7389 35785 7423 35819
rect 8493 35785 8527 35819
rect 11621 35785 11655 35819
rect 7205 35581 7239 35615
rect 8309 35581 8343 35615
rect 8861 35581 8895 35615
rect 11897 35513 11931 35547
rect 7849 35445 7883 35479
rect 2329 35241 2363 35275
rect 4261 35241 4295 35275
rect 5365 35241 5399 35275
rect 7665 35241 7699 35275
rect 9934 35173 9968 35207
rect 2145 35105 2179 35139
rect 4077 35105 4111 35139
rect 5181 35105 5215 35139
rect 6377 35105 6411 35139
rect 7481 35105 7515 35139
rect 9689 35105 9723 35139
rect 6561 34969 6595 35003
rect 5733 34901 5767 34935
rect 8125 34901 8159 34935
rect 11069 34901 11103 34935
rect 1593 34697 1627 34731
rect 2053 34697 2087 34731
rect 3801 34697 3835 34731
rect 5733 34697 5767 34731
rect 7021 34697 7055 34731
rect 7757 34697 7791 34731
rect 9413 34697 9447 34731
rect 10333 34697 10367 34731
rect 13645 34697 13679 34731
rect 2697 34629 2731 34663
rect 4261 34629 4295 34663
rect 2421 34561 2455 34595
rect 10977 34561 11011 34595
rect 11161 34561 11195 34595
rect 11529 34561 11563 34595
rect 1409 34493 1443 34527
rect 2513 34493 2547 34527
rect 3157 34493 3191 34527
rect 3617 34493 3651 34527
rect 5549 34493 5583 34527
rect 6469 34493 6503 34527
rect 6837 34493 6871 34527
rect 7389 34493 7423 34527
rect 8033 34493 8067 34527
rect 9965 34493 9999 34527
rect 10885 34493 10919 34527
rect 13461 34493 13495 34527
rect 14013 34493 14047 34527
rect 5181 34425 5215 34459
rect 8300 34425 8334 34459
rect 4629 34357 4663 34391
rect 10517 34357 10551 34391
rect 1593 34153 1627 34187
rect 2697 34153 2731 34187
rect 4261 34153 4295 34187
rect 5457 34153 5491 34187
rect 6929 34153 6963 34187
rect 8033 34153 8067 34187
rect 9873 34153 9907 34187
rect 11897 34153 11931 34187
rect 1409 34017 1443 34051
rect 2513 34017 2547 34051
rect 4077 34017 4111 34051
rect 5273 34017 5307 34051
rect 6745 34017 6779 34051
rect 7849 34017 7883 34051
rect 10784 34017 10818 34051
rect 10517 33949 10551 33983
rect 7389 33813 7423 33847
rect 8401 33813 8435 33847
rect 10333 33813 10367 33847
rect 1593 33609 1627 33643
rect 1961 33609 1995 33643
rect 2973 33609 3007 33643
rect 11161 33609 11195 33643
rect 6837 33473 6871 33507
rect 9689 33473 9723 33507
rect 10609 33473 10643 33507
rect 10793 33473 10827 33507
rect 1409 33405 1443 33439
rect 2789 33405 2823 33439
rect 6285 33337 6319 33371
rect 7104 33337 7138 33371
rect 10057 33337 10091 33371
rect 10517 33337 10551 33371
rect 2421 33269 2455 33303
rect 3341 33269 3375 33303
rect 4169 33269 4203 33303
rect 5365 33269 5399 33303
rect 6653 33269 6687 33303
rect 8217 33269 8251 33303
rect 10149 33269 10183 33303
rect 11529 33269 11563 33303
rect 12449 33269 12483 33303
rect 2789 33065 2823 33099
rect 6837 33065 6871 33099
rect 7849 33065 7883 33099
rect 10241 33065 10275 33099
rect 1685 32997 1719 33031
rect 11805 32997 11839 33031
rect 12265 32997 12299 33031
rect 1409 32929 1443 32963
rect 6929 32929 6963 32963
rect 8401 32929 8435 32963
rect 9505 32929 9539 32963
rect 10701 32929 10735 32963
rect 12357 32929 12391 32963
rect 7113 32861 7147 32895
rect 7573 32861 7607 32895
rect 8493 32861 8527 32895
rect 8585 32861 8619 32895
rect 10793 32861 10827 32895
rect 10977 32861 11011 32895
rect 12541 32861 12575 32895
rect 6469 32725 6503 32759
rect 8033 32725 8067 32759
rect 9137 32725 9171 32759
rect 10333 32725 10367 32759
rect 11897 32725 11931 32759
rect 13001 32725 13035 32759
rect 6193 32521 6227 32555
rect 8861 32521 8895 32555
rect 9965 32521 9999 32555
rect 10517 32521 10551 32555
rect 13553 32521 13587 32555
rect 6469 32453 6503 32487
rect 8677 32453 8711 32487
rect 7481 32385 7515 32419
rect 9413 32385 9447 32419
rect 10977 32385 11011 32419
rect 11069 32385 11103 32419
rect 13093 32385 13127 32419
rect 3525 32317 3559 32351
rect 3985 32317 4019 32351
rect 7297 32317 7331 32351
rect 9229 32317 9263 32351
rect 12817 32317 12851 32351
rect 3893 32249 3927 32283
rect 4252 32249 4286 32283
rect 7205 32249 7239 32283
rect 11897 32249 11931 32283
rect 12909 32249 12943 32283
rect 1685 32181 1719 32215
rect 5365 32181 5399 32215
rect 6837 32181 6871 32215
rect 7849 32181 7883 32215
rect 8217 32181 8251 32215
rect 9321 32181 9355 32215
rect 10333 32181 10367 32215
rect 10885 32181 10919 32215
rect 12173 32181 12207 32215
rect 12449 32181 12483 32215
rect 7481 31977 7515 32011
rect 9689 31977 9723 32011
rect 10793 31977 10827 32011
rect 11161 31977 11195 32011
rect 1685 31909 1719 31943
rect 5264 31909 5298 31943
rect 7849 31909 7883 31943
rect 8953 31909 8987 31943
rect 9505 31909 9539 31943
rect 11682 31909 11716 31943
rect 1409 31841 1443 31875
rect 4997 31841 5031 31875
rect 6929 31841 6963 31875
rect 7941 31841 7975 31875
rect 10057 31841 10091 31875
rect 11437 31841 11471 31875
rect 7389 31773 7423 31807
rect 8125 31773 8159 31807
rect 10149 31773 10183 31807
rect 10241 31773 10275 31807
rect 6377 31705 6411 31739
rect 8585 31637 8619 31671
rect 12817 31637 12851 31671
rect 5089 31433 5123 31467
rect 6653 31433 6687 31467
rect 7021 31433 7055 31467
rect 7481 31433 7515 31467
rect 8585 31433 8619 31467
rect 10241 31433 10275 31467
rect 11437 31433 11471 31467
rect 11989 31433 12023 31467
rect 12633 31433 12667 31467
rect 1685 31365 1719 31399
rect 8125 31297 8159 31331
rect 9413 31297 9447 31331
rect 10885 31297 10919 31331
rect 10977 31297 11011 31331
rect 5917 31229 5951 31263
rect 7941 31229 7975 31263
rect 6285 31161 6319 31195
rect 8033 31161 8067 31195
rect 5457 31093 5491 31127
rect 7573 31093 7607 31127
rect 9229 31093 9263 31127
rect 9873 31093 9907 31127
rect 10425 31093 10459 31127
rect 10793 31093 10827 31127
rect 6377 30889 6411 30923
rect 6837 30889 6871 30923
rect 8033 30889 8067 30923
rect 8493 30889 8527 30923
rect 10057 30889 10091 30923
rect 11069 30889 11103 30923
rect 7665 30821 7699 30855
rect 10793 30821 10827 30855
rect 11805 30821 11839 30855
rect 3893 30753 3927 30787
rect 4537 30753 4571 30787
rect 6929 30753 6963 30787
rect 8401 30753 8435 30787
rect 10149 30753 10183 30787
rect 11713 30753 11747 30787
rect 4629 30685 4663 30719
rect 4813 30685 4847 30719
rect 7021 30685 7055 30719
rect 8585 30685 8619 30719
rect 10241 30685 10275 30719
rect 11897 30685 11931 30719
rect 6469 30617 6503 30651
rect 9689 30617 9723 30651
rect 11345 30617 11379 30651
rect 4169 30549 4203 30583
rect 6009 30549 6043 30583
rect 6193 30345 6227 30379
rect 10057 30345 10091 30379
rect 10793 30345 10827 30379
rect 11345 30345 11379 30379
rect 11805 30345 11839 30379
rect 12081 30345 12115 30379
rect 2237 30277 2271 30311
rect 6285 30277 6319 30311
rect 9045 30277 9079 30311
rect 1593 30209 1627 30243
rect 3065 30209 3099 30243
rect 3525 30209 3559 30243
rect 1409 30141 1443 30175
rect 6469 30141 6503 30175
rect 7665 30141 7699 30175
rect 3433 30073 3467 30107
rect 3792 30073 3826 30107
rect 7910 30073 7944 30107
rect 10425 30073 10459 30107
rect 4905 30005 4939 30039
rect 5457 30005 5491 30039
rect 7113 30005 7147 30039
rect 7573 30005 7607 30039
rect 9781 30005 9815 30039
rect 3893 29801 3927 29835
rect 5641 29801 5675 29835
rect 7113 29801 7147 29835
rect 7573 29801 7607 29835
rect 8585 29801 8619 29835
rect 11069 29801 11103 29835
rect 2789 29733 2823 29767
rect 6745 29733 6779 29767
rect 9934 29733 9968 29767
rect 4445 29665 4479 29699
rect 6009 29665 6043 29699
rect 6101 29665 6135 29699
rect 8309 29665 8343 29699
rect 9689 29665 9723 29699
rect 2881 29597 2915 29631
rect 3065 29597 3099 29631
rect 4537 29597 4571 29631
rect 4721 29597 4755 29631
rect 6193 29597 6227 29631
rect 7665 29597 7699 29631
rect 7849 29597 7883 29631
rect 1685 29461 1719 29495
rect 2421 29461 2455 29495
rect 3525 29461 3559 29495
rect 4077 29461 4111 29495
rect 5181 29461 5215 29495
rect 7205 29461 7239 29495
rect 3249 29257 3283 29291
rect 4353 29257 4387 29291
rect 4445 29257 4479 29291
rect 4813 29257 4847 29291
rect 7849 29257 7883 29291
rect 9505 29257 9539 29291
rect 2513 29189 2547 29223
rect 3157 29121 3191 29155
rect 3801 29121 3835 29155
rect 6285 29189 6319 29223
rect 5365 29121 5399 29155
rect 7297 29121 7331 29155
rect 7481 29121 7515 29155
rect 10241 29121 10275 29155
rect 1409 29053 1443 29087
rect 3617 29053 3651 29087
rect 4445 29053 4479 29087
rect 5181 29053 5215 29087
rect 5273 29053 5307 29087
rect 8217 29053 8251 29087
rect 9229 29053 9263 29087
rect 10057 29053 10091 29087
rect 10149 29053 10183 29087
rect 1685 28985 1719 29019
rect 4721 28985 4755 29019
rect 5917 28985 5951 29019
rect 6653 28985 6687 29019
rect 7205 28985 7239 29019
rect 8861 28985 8895 29019
rect 3709 28917 3743 28951
rect 6837 28917 6871 28951
rect 9689 28917 9723 28951
rect 10793 28917 10827 28951
rect 2789 28713 2823 28747
rect 4353 28713 4387 28747
rect 4721 28713 4755 28747
rect 6193 28713 6227 28747
rect 6929 28713 6963 28747
rect 7665 28713 7699 28747
rect 9873 28713 9907 28747
rect 2513 28645 2547 28679
rect 6101 28645 6135 28679
rect 7297 28645 7331 28679
rect 11498 28645 11532 28679
rect 1409 28577 1443 28611
rect 8493 28577 8527 28611
rect 10609 28577 10643 28611
rect 11253 28577 11287 28611
rect 6285 28509 6319 28543
rect 1593 28441 1627 28475
rect 3893 28441 3927 28475
rect 9229 28441 9263 28475
rect 10425 28441 10459 28475
rect 3341 28373 3375 28407
rect 5181 28373 5215 28407
rect 5549 28373 5583 28407
rect 5733 28373 5767 28407
rect 8309 28373 8343 28407
rect 8861 28373 8895 28407
rect 12633 28373 12667 28407
rect 5457 28169 5491 28203
rect 5825 28169 5859 28203
rect 6101 28169 6135 28203
rect 9965 28169 9999 28203
rect 11253 28169 11287 28203
rect 11621 28169 11655 28203
rect 2053 28033 2087 28067
rect 2421 28033 2455 28067
rect 6653 28033 6687 28067
rect 7573 28033 7607 28067
rect 8401 28033 8435 28067
rect 1409 27965 1443 27999
rect 8585 27965 8619 27999
rect 8841 27965 8875 27999
rect 1593 27829 1627 27863
rect 7021 27829 7055 27863
rect 7389 27829 7423 27863
rect 7481 27829 7515 27863
rect 8125 27829 8159 27863
rect 10609 27829 10643 27863
rect 4077 27625 4111 27659
rect 8493 27625 8527 27659
rect 9689 27625 9723 27659
rect 11621 27625 11655 27659
rect 1685 27557 1719 27591
rect 6101 27557 6135 27591
rect 6469 27557 6503 27591
rect 10793 27557 10827 27591
rect 1409 27489 1443 27523
rect 4445 27489 4479 27523
rect 6745 27489 6779 27523
rect 7380 27489 7414 27523
rect 10057 27489 10091 27523
rect 11437 27489 11471 27523
rect 11980 27557 12014 27591
rect 4537 27421 4571 27455
rect 4721 27421 4755 27455
rect 7113 27421 7147 27455
rect 10149 27421 10183 27455
rect 10241 27421 10275 27455
rect 11621 27421 11655 27455
rect 11713 27421 11747 27455
rect 6561 27353 6595 27387
rect 9045 27285 9079 27319
rect 9413 27285 9447 27319
rect 11253 27285 11287 27319
rect 13093 27285 13127 27319
rect 1593 27081 1627 27115
rect 3525 27081 3559 27115
rect 3985 27081 4019 27115
rect 5641 27081 5675 27115
rect 8769 27081 8803 27115
rect 10425 27081 10459 27115
rect 12081 27081 12115 27115
rect 8953 27013 8987 27047
rect 11805 27013 11839 27047
rect 3157 26945 3191 26979
rect 4537 26945 4571 26979
rect 7389 26945 7423 26979
rect 9505 26945 9539 26979
rect 11161 26945 11195 26979
rect 6653 26877 6687 26911
rect 9413 26877 9447 26911
rect 10977 26877 11011 26911
rect 3893 26809 3927 26843
rect 4445 26809 4479 26843
rect 5733 26809 5767 26843
rect 6285 26809 6319 26843
rect 7205 26809 7239 26843
rect 7297 26809 7331 26843
rect 10885 26809 10919 26843
rect 4353 26741 4387 26775
rect 5089 26741 5123 26775
rect 6837 26741 6871 26775
rect 7941 26741 7975 26775
rect 8401 26741 8435 26775
rect 9321 26741 9355 26775
rect 9965 26741 9999 26775
rect 10517 26741 10551 26775
rect 4629 26537 4663 26571
rect 6653 26537 6687 26571
rect 7297 26537 7331 26571
rect 7573 26537 7607 26571
rect 8033 26537 8067 26571
rect 9137 26537 9171 26571
rect 9965 26537 9999 26571
rect 11897 26537 11931 26571
rect 5540 26469 5574 26503
rect 8401 26401 8435 26435
rect 10885 26401 10919 26435
rect 5273 26333 5307 26367
rect 8493 26333 8527 26367
rect 8677 26333 8711 26367
rect 9505 26333 9539 26367
rect 10977 26333 11011 26367
rect 11069 26333 11103 26367
rect 5181 26265 5215 26299
rect 10241 26265 10275 26299
rect 11529 26265 11563 26299
rect 4353 26197 4387 26231
rect 10517 26197 10551 26231
rect 3985 25993 4019 26027
rect 5457 25993 5491 26027
rect 8033 25993 8067 26027
rect 8769 25993 8803 26027
rect 11621 25993 11655 26027
rect 10333 25925 10367 25959
rect 11989 25925 12023 25959
rect 1593 25857 1627 25891
rect 7481 25857 7515 25891
rect 9413 25857 9447 25891
rect 11069 25857 11103 25891
rect 11253 25857 11287 25891
rect 1409 25789 1443 25823
rect 3617 25789 3651 25823
rect 4077 25789 4111 25823
rect 4333 25789 4367 25823
rect 6653 25789 6687 25823
rect 7205 25789 7239 25823
rect 8493 25789 8527 25823
rect 10517 25789 10551 25823
rect 10977 25789 11011 25823
rect 6285 25721 6319 25755
rect 7297 25721 7331 25755
rect 9137 25721 9171 25755
rect 2237 25653 2271 25687
rect 6837 25653 6871 25687
rect 9229 25653 9263 25687
rect 9781 25653 9815 25687
rect 10149 25653 10183 25687
rect 10609 25653 10643 25687
rect 12541 25653 12575 25687
rect 5457 25449 5491 25483
rect 6469 25449 6503 25483
rect 6837 25449 6871 25483
rect 8309 25449 8343 25483
rect 9229 25449 9263 25483
rect 10793 25449 10827 25483
rect 6101 25381 6135 25415
rect 11805 25381 11839 25415
rect 4077 25313 4111 25347
rect 4333 25313 4367 25347
rect 6745 25313 6779 25347
rect 6837 25313 6871 25347
rect 7185 25313 7219 25347
rect 10333 25313 10367 25347
rect 12725 25313 12759 25347
rect 12817 25313 12851 25347
rect 6929 25245 6963 25279
rect 10885 25245 10919 25279
rect 10977 25245 11011 25279
rect 12909 25245 12943 25279
rect 11529 25177 11563 25211
rect 12265 25177 12299 25211
rect 6561 25109 6595 25143
rect 9873 25109 9907 25143
rect 10425 25109 10459 25143
rect 12357 25109 12391 25143
rect 3801 24905 3835 24939
rect 5181 24905 5215 24939
rect 6193 24905 6227 24939
rect 6377 24905 6411 24939
rect 6653 24905 6687 24939
rect 9137 24905 9171 24939
rect 10149 24905 10183 24939
rect 13829 24905 13863 24939
rect 6009 24837 6043 24871
rect 5641 24769 5675 24803
rect 5825 24769 5859 24803
rect 5089 24701 5123 24735
rect 6837 24837 6871 24871
rect 12265 24837 12299 24871
rect 13277 24837 13311 24871
rect 6377 24769 6411 24803
rect 7297 24769 7331 24803
rect 7481 24769 7515 24803
rect 8309 24769 8343 24803
rect 8585 24769 8619 24803
rect 9689 24769 9723 24803
rect 11345 24769 11379 24803
rect 13093 24769 13127 24803
rect 7849 24701 7883 24735
rect 8953 24701 8987 24735
rect 11069 24701 11103 24735
rect 4721 24633 4755 24667
rect 5549 24633 5583 24667
rect 6009 24633 6043 24667
rect 7205 24633 7239 24667
rect 9597 24633 9631 24667
rect 11161 24633 11195 24667
rect 11897 24633 11931 24667
rect 12909 24633 12943 24667
rect 14197 24769 14231 24803
rect 13461 24633 13495 24667
rect 4169 24565 4203 24599
rect 9505 24565 9539 24599
rect 10517 24565 10551 24599
rect 10701 24565 10735 24599
rect 12449 24565 12483 24599
rect 12817 24565 12851 24599
rect 13277 24565 13311 24599
rect 5273 24361 5307 24395
rect 7573 24361 7607 24395
rect 9965 24361 9999 24395
rect 10517 24361 10551 24395
rect 11437 24361 11471 24395
rect 5908 24293 5942 24327
rect 11866 24293 11900 24327
rect 10425 24225 10459 24259
rect 5641 24157 5675 24191
rect 10609 24157 10643 24191
rect 11621 24157 11655 24191
rect 7021 24089 7055 24123
rect 9137 24021 9171 24055
rect 10057 24021 10091 24055
rect 11069 24021 11103 24055
rect 13001 24021 13035 24055
rect 5733 23817 5767 23851
rect 8677 23817 8711 23851
rect 10793 23817 10827 23851
rect 11069 23817 11103 23851
rect 11621 23817 11655 23851
rect 13001 23681 13035 23715
rect 8769 23613 8803 23647
rect 9025 23613 9059 23647
rect 12173 23613 12207 23647
rect 12909 23613 12943 23647
rect 13461 23613 13495 23647
rect 6101 23477 6135 23511
rect 10149 23477 10183 23511
rect 12449 23477 12483 23511
rect 12817 23477 12851 23511
rect 13829 23477 13863 23511
rect 5181 23273 5215 23307
rect 9321 23273 9355 23307
rect 10977 23273 11011 23307
rect 11621 23273 11655 23307
rect 10149 23205 10183 23239
rect 10885 23137 10919 23171
rect 12081 23137 12115 23171
rect 12337 23137 12371 23171
rect 5273 23069 5307 23103
rect 5457 23069 5491 23103
rect 11161 23069 11195 23103
rect 10517 23001 10551 23035
rect 2605 22933 2639 22967
rect 4813 22933 4847 22967
rect 5825 22933 5859 22967
rect 7665 22933 7699 22967
rect 8861 22933 8895 22967
rect 13461 22933 13495 22967
rect 4905 22729 4939 22763
rect 6285 22729 6319 22763
rect 7573 22729 7607 22763
rect 9137 22729 9171 22763
rect 9321 22729 9355 22763
rect 10609 22729 10643 22763
rect 10885 22729 10919 22763
rect 11345 22729 11379 22763
rect 12173 22729 12207 22763
rect 7481 22661 7515 22695
rect 2513 22593 2547 22627
rect 5733 22593 5767 22627
rect 6561 22593 6595 22627
rect 8033 22593 8067 22627
rect 8125 22593 8159 22627
rect 9873 22593 9907 22627
rect 4537 22525 4571 22559
rect 5549 22525 5583 22559
rect 9781 22525 9815 22559
rect 2421 22457 2455 22491
rect 2780 22457 2814 22491
rect 3893 22389 3927 22423
rect 5181 22389 5215 22423
rect 5641 22389 5675 22423
rect 7113 22389 7147 22423
rect 7941 22389 7975 22423
rect 9689 22389 9723 22423
rect 12633 22389 12667 22423
rect 8493 22185 8527 22219
rect 9689 22185 9723 22219
rect 10149 22185 10183 22219
rect 4322 22117 4356 22151
rect 2329 22049 2363 22083
rect 2789 22049 2823 22083
rect 2881 22049 2915 22083
rect 7113 22049 7147 22083
rect 7380 22049 7414 22083
rect 10057 22049 10091 22083
rect 12348 22049 12382 22083
rect 2973 21981 3007 22015
rect 4077 21981 4111 22015
rect 10241 21981 10275 22015
rect 12081 21981 12115 22015
rect 2421 21845 2455 21879
rect 3801 21845 3835 21879
rect 5457 21845 5491 21879
rect 6101 21845 6135 21879
rect 9413 21845 9447 21879
rect 13461 21845 13495 21879
rect 5365 21641 5399 21675
rect 6285 21641 6319 21675
rect 7849 21641 7883 21675
rect 9781 21641 9815 21675
rect 10425 21641 10459 21675
rect 12173 21641 12207 21675
rect 12633 21641 12667 21675
rect 13645 21641 13679 21675
rect 3985 21573 4019 21607
rect 3065 21505 3099 21539
rect 4445 21505 4479 21539
rect 4537 21505 4571 21539
rect 4997 21505 5031 21539
rect 6653 21505 6687 21539
rect 7389 21505 7423 21539
rect 8493 21505 8527 21539
rect 2329 21437 2363 21471
rect 3525 21437 3559 21471
rect 3893 21437 3927 21471
rect 8309 21437 8343 21471
rect 13461 21437 13495 21471
rect 14013 21437 14047 21471
rect 1961 21369 1995 21403
rect 2789 21369 2823 21403
rect 5549 21369 5583 21403
rect 2421 21301 2455 21335
rect 2881 21301 2915 21335
rect 4353 21301 4387 21335
rect 7757 21301 7791 21335
rect 8217 21301 8251 21335
rect 10057 21301 10091 21335
rect 2973 21097 3007 21131
rect 3249 21097 3283 21131
rect 4077 21097 4111 21131
rect 4445 21097 4479 21131
rect 4537 21097 4571 21131
rect 7205 21097 7239 21131
rect 7941 21097 7975 21131
rect 8309 21097 8343 21131
rect 2421 21029 2455 21063
rect 6070 21029 6104 21063
rect 2145 20961 2179 20995
rect 5825 20961 5859 20995
rect 10508 20961 10542 20995
rect 4629 20893 4663 20927
rect 9413 20893 9447 20927
rect 10241 20893 10275 20927
rect 3893 20825 3927 20859
rect 11621 20757 11655 20791
rect 2145 20553 2179 20587
rect 3341 20553 3375 20587
rect 4537 20553 4571 20587
rect 6193 20553 6227 20587
rect 11253 20553 11287 20587
rect 3709 20485 3743 20519
rect 3985 20417 4019 20451
rect 5089 20417 5123 20451
rect 6837 20417 6871 20451
rect 9321 20417 9355 20451
rect 4445 20281 4479 20315
rect 4905 20281 4939 20315
rect 6653 20281 6687 20315
rect 7082 20281 7116 20315
rect 9229 20281 9263 20315
rect 9588 20281 9622 20315
rect 4997 20213 5031 20247
rect 5917 20213 5951 20247
rect 8217 20213 8251 20247
rect 10701 20213 10735 20247
rect 11621 20213 11655 20247
rect 4905 20009 4939 20043
rect 5917 20009 5951 20043
rect 6929 20009 6963 20043
rect 9137 20009 9171 20043
rect 10333 20009 10367 20043
rect 11897 20009 11931 20043
rect 10784 19941 10818 19975
rect 6285 19873 6319 19907
rect 6377 19873 6411 19907
rect 10517 19873 10551 19907
rect 6561 19805 6595 19839
rect 13001 19805 13035 19839
rect 2605 19669 2639 19703
rect 4537 19669 4571 19703
rect 8677 19669 8711 19703
rect 9505 19669 9539 19703
rect 9873 19669 9907 19703
rect 12541 19669 12575 19703
rect 5641 19465 5675 19499
rect 10333 19397 10367 19431
rect 2605 19329 2639 19363
rect 10057 19329 10091 19363
rect 10977 19329 11011 19363
rect 12909 19329 12943 19363
rect 13001 19329 13035 19363
rect 9781 19261 9815 19295
rect 11345 19261 11379 19295
rect 2513 19193 2547 19227
rect 2850 19193 2884 19227
rect 7481 19193 7515 19227
rect 7573 19193 7607 19227
rect 10793 19193 10827 19227
rect 12173 19193 12207 19227
rect 3985 19125 4019 19159
rect 6009 19125 6043 19159
rect 6377 19125 6411 19159
rect 8861 19125 8895 19159
rect 9413 19125 9447 19159
rect 9873 19125 9907 19159
rect 10701 19125 10735 19159
rect 11805 19125 11839 19159
rect 12449 19125 12483 19159
rect 12817 19125 12851 19159
rect 2605 18921 2639 18955
rect 6285 18921 6319 18955
rect 7113 18921 7147 18955
rect 7941 18921 7975 18955
rect 8493 18921 8527 18955
rect 9689 18921 9723 18955
rect 11161 18921 11195 18955
rect 1685 18853 1719 18887
rect 9505 18853 9539 18887
rect 10057 18853 10091 18887
rect 1409 18785 1443 18819
rect 6193 18785 6227 18819
rect 8401 18785 8435 18819
rect 11785 18785 11819 18819
rect 6377 18717 6411 18751
rect 8585 18717 8619 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 11529 18717 11563 18751
rect 8033 18649 8067 18683
rect 5273 18581 5307 18615
rect 5825 18581 5859 18615
rect 7573 18581 7607 18615
rect 9137 18581 9171 18615
rect 10701 18581 10735 18615
rect 12909 18581 12943 18615
rect 3893 18377 3927 18411
rect 5089 18377 5123 18411
rect 6193 18377 6227 18411
rect 8585 18377 8619 18411
rect 9781 18377 9815 18411
rect 13829 18377 13863 18411
rect 1685 18309 1719 18343
rect 7113 18309 7147 18343
rect 8677 18309 8711 18343
rect 12173 18309 12207 18343
rect 4721 18241 4755 18275
rect 5825 18241 5859 18275
rect 7573 18241 7607 18275
rect 7665 18241 7699 18275
rect 9229 18241 9263 18275
rect 10885 18241 10919 18275
rect 13093 18241 13127 18275
rect 2513 18173 2547 18207
rect 5641 18173 5675 18207
rect 9045 18173 9079 18207
rect 9137 18173 9171 18207
rect 10793 18173 10827 18207
rect 11897 18173 11931 18207
rect 12817 18173 12851 18207
rect 2421 18105 2455 18139
rect 2758 18105 2792 18139
rect 5549 18105 5583 18139
rect 10701 18105 10735 18139
rect 13461 18105 13495 18139
rect 5181 18037 5215 18071
rect 6653 18037 6687 18071
rect 7481 18037 7515 18071
rect 8217 18037 8251 18071
rect 10149 18037 10183 18071
rect 10333 18037 10367 18071
rect 11437 18037 11471 18071
rect 12449 18037 12483 18071
rect 12909 18037 12943 18071
rect 8217 17833 8251 17867
rect 9689 17833 9723 17867
rect 10149 17833 10183 17867
rect 10793 17833 10827 17867
rect 11529 17833 11563 17867
rect 11989 17833 12023 17867
rect 4414 17765 4448 17799
rect 9505 17765 9539 17799
rect 12081 17765 12115 17799
rect 2329 17697 2363 17731
rect 2789 17697 2823 17731
rect 7104 17697 7138 17731
rect 10057 17697 10091 17731
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4169 17629 4203 17663
rect 6837 17629 6871 17663
rect 10241 17629 10275 17663
rect 12265 17629 12299 17663
rect 11621 17561 11655 17595
rect 2421 17493 2455 17527
rect 3525 17493 3559 17527
rect 5549 17493 5583 17527
rect 6101 17493 6135 17527
rect 6745 17493 6779 17527
rect 8769 17493 8803 17527
rect 11069 17493 11103 17527
rect 12725 17493 12759 17527
rect 13001 17493 13035 17527
rect 3433 17289 3467 17323
rect 4905 17289 4939 17323
rect 8125 17289 8159 17323
rect 9413 17289 9447 17323
rect 9781 17289 9815 17323
rect 10701 17289 10735 17323
rect 11897 17289 11931 17323
rect 12265 17289 12299 17323
rect 12449 17289 12483 17323
rect 2513 17221 2547 17255
rect 3341 17221 3375 17255
rect 4997 17221 5031 17255
rect 10793 17221 10827 17255
rect 1593 17153 1627 17187
rect 3893 17153 3927 17187
rect 4077 17153 4111 17187
rect 5549 17153 5583 17187
rect 7389 17153 7423 17187
rect 8033 17153 8067 17187
rect 8769 17153 8803 17187
rect 11345 17153 11379 17187
rect 13001 17153 13035 17187
rect 1409 17085 1443 17119
rect 5365 17085 5399 17119
rect 11253 17085 11287 17119
rect 12817 17085 12851 17119
rect 2973 17017 3007 17051
rect 3801 17017 3835 17051
rect 6837 17017 6871 17051
rect 10057 17017 10091 17051
rect 4445 16949 4479 16983
rect 5457 16949 5491 16983
rect 6561 16949 6595 16983
rect 8493 16949 8527 16983
rect 8585 16949 8619 16983
rect 11161 16949 11195 16983
rect 12909 16949 12943 16983
rect 13461 16949 13495 16983
rect 1593 16745 1627 16779
rect 2329 16745 2363 16779
rect 2421 16745 2455 16779
rect 3709 16745 3743 16779
rect 3801 16745 3835 16779
rect 4169 16745 4203 16779
rect 4537 16745 4571 16779
rect 4629 16745 4663 16779
rect 5549 16745 5583 16779
rect 7849 16745 7883 16779
rect 8769 16745 8803 16779
rect 10425 16745 10459 16779
rect 11897 16745 11931 16779
rect 13369 16745 13403 16779
rect 3525 16677 3559 16711
rect 6000 16677 6034 16711
rect 10885 16677 10919 16711
rect 2789 16609 2823 16643
rect 3709 16609 3743 16643
rect 5733 16609 5767 16643
rect 8217 16609 8251 16643
rect 10333 16609 10367 16643
rect 10793 16609 10827 16643
rect 11437 16609 11471 16643
rect 12245 16609 12279 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 4721 16541 4755 16575
rect 5181 16541 5215 16575
rect 9965 16541 9999 16575
rect 10977 16541 11011 16575
rect 11989 16541 12023 16575
rect 7113 16405 7147 16439
rect 2881 16201 2915 16235
rect 4537 16201 4571 16235
rect 4997 16201 5031 16235
rect 7021 16201 7055 16235
rect 9137 16201 9171 16235
rect 10793 16201 10827 16235
rect 12081 16201 12115 16235
rect 4261 16133 4295 16167
rect 9965 16133 9999 16167
rect 2513 16065 2547 16099
rect 5641 16065 5675 16099
rect 5825 16065 5859 16099
rect 7665 16065 7699 16099
rect 11437 16065 11471 16099
rect 7757 15997 7791 16031
rect 8024 15997 8058 16031
rect 10333 15997 10367 16031
rect 11161 15997 11195 16031
rect 5549 15929 5583 15963
rect 6561 15929 6595 15963
rect 10609 15929 10643 15963
rect 11253 15929 11287 15963
rect 3249 15861 3283 15895
rect 5181 15861 5215 15895
rect 6193 15861 6227 15895
rect 12633 15861 12667 15895
rect 5273 15657 5307 15691
rect 7757 15657 7791 15691
rect 8033 15657 8067 15691
rect 9045 15657 9079 15691
rect 10057 15657 10091 15691
rect 10517 15657 10551 15691
rect 11161 15657 11195 15691
rect 13001 15657 13035 15691
rect 6009 15521 6043 15555
rect 8401 15521 8435 15555
rect 8493 15521 8527 15555
rect 10425 15521 10459 15555
rect 11877 15521 11911 15555
rect 6101 15453 6135 15487
rect 6285 15453 6319 15487
rect 8585 15453 8619 15487
rect 10701 15453 10735 15487
rect 11621 15453 11655 15487
rect 9965 15385 9999 15419
rect 5641 15317 5675 15351
rect 6009 15113 6043 15147
rect 6377 15113 6411 15147
rect 8125 15113 8159 15147
rect 8585 15113 8619 15147
rect 8677 15113 8711 15147
rect 8861 15113 8895 15147
rect 10425 15113 10459 15147
rect 1593 14977 1627 15011
rect 1409 14909 1443 14943
rect 5733 14909 5767 14943
rect 9965 15045 9999 15079
rect 9413 14977 9447 15011
rect 11069 14977 11103 15011
rect 9321 14909 9355 14943
rect 8585 14841 8619 14875
rect 9229 14841 9263 14875
rect 10793 14841 10827 14875
rect 11989 14841 12023 14875
rect 2513 14773 2547 14807
rect 7757 14773 7791 14807
rect 10241 14773 10275 14807
rect 10885 14773 10919 14807
rect 11621 14773 11655 14807
rect 2421 14569 2455 14603
rect 3433 14569 3467 14603
rect 4077 14569 4111 14603
rect 4445 14569 4479 14603
rect 6101 14569 6135 14603
rect 8309 14569 8343 14603
rect 8953 14569 8987 14603
rect 9689 14569 9723 14603
rect 11161 14569 11195 14603
rect 6009 14501 6043 14535
rect 13553 14501 13587 14535
rect 2789 14433 2823 14467
rect 7573 14433 7607 14467
rect 13277 14433 13311 14467
rect 2881 14365 2915 14399
rect 3065 14365 3099 14399
rect 3893 14365 3927 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 6193 14365 6227 14399
rect 7665 14365 7699 14399
rect 7849 14365 7883 14399
rect 7021 14297 7055 14331
rect 10793 14297 10827 14331
rect 1685 14229 1719 14263
rect 2237 14229 2271 14263
rect 5641 14229 5675 14263
rect 7205 14229 7239 14263
rect 10425 14229 10459 14263
rect 1685 14025 1719 14059
rect 2145 14025 2179 14059
rect 3249 14025 3283 14059
rect 3617 14025 3651 14059
rect 5089 14025 5123 14059
rect 5733 14025 5767 14059
rect 6101 14025 6135 14059
rect 6653 14025 6687 14059
rect 2697 13889 2731 13923
rect 3709 13889 3743 13923
rect 6929 13889 6963 13923
rect 2053 13821 2087 13855
rect 2605 13821 2639 13855
rect 7185 13821 7219 13855
rect 8861 13821 8895 13855
rect 13277 13821 13311 13855
rect 3954 13753 3988 13787
rect 2513 13685 2547 13719
rect 8309 13685 8343 13719
rect 2237 13481 2271 13515
rect 4077 13481 4111 13515
rect 5641 13481 5675 13515
rect 6653 13481 6687 13515
rect 8217 13481 8251 13515
rect 4537 13413 4571 13447
rect 11980 13413 12014 13447
rect 2789 13345 2823 13379
rect 2881 13345 2915 13379
rect 3617 13345 3651 13379
rect 4445 13345 4479 13379
rect 7205 13345 7239 13379
rect 10333 13345 10367 13379
rect 3065 13277 3099 13311
rect 4629 13277 4663 13311
rect 7297 13277 7331 13311
rect 7481 13277 7515 13311
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 11713 13277 11747 13311
rect 1869 13209 1903 13243
rect 2421 13209 2455 13243
rect 3617 13209 3651 13243
rect 6837 13209 6871 13243
rect 7849 13209 7883 13243
rect 3709 13141 3743 13175
rect 5181 13141 5215 13175
rect 9965 13141 9999 13175
rect 10977 13141 11011 13175
rect 13093 13141 13127 13175
rect 2145 12937 2179 12971
rect 4261 12937 4295 12971
rect 7389 12937 7423 12971
rect 10517 12937 10551 12971
rect 11529 12937 11563 12971
rect 7113 12869 7147 12903
rect 10425 12869 10459 12903
rect 12633 12869 12667 12903
rect 2237 12801 2271 12835
rect 5549 12801 5583 12835
rect 7941 12801 7975 12835
rect 10977 12801 11011 12835
rect 11161 12801 11195 12835
rect 5457 12733 5491 12767
rect 6009 12733 6043 12767
rect 8033 12733 8067 12767
rect 8300 12733 8334 12767
rect 1777 12665 1811 12699
rect 2482 12665 2516 12699
rect 5365 12665 5399 12699
rect 6377 12665 6411 12699
rect 3617 12597 3651 12631
rect 4629 12597 4663 12631
rect 4997 12597 5031 12631
rect 9413 12597 9447 12631
rect 10057 12597 10091 12631
rect 10885 12597 10919 12631
rect 11989 12597 12023 12631
rect 6561 12393 6595 12427
rect 7113 12393 7147 12427
rect 7481 12393 7515 12427
rect 8401 12393 8435 12427
rect 9965 12393 9999 12427
rect 10057 12393 10091 12427
rect 1685 12325 1719 12359
rect 5426 12325 5460 12359
rect 11866 12325 11900 12359
rect 1409 12257 1443 12291
rect 5089 12257 5123 12291
rect 7941 12257 7975 12291
rect 10425 12257 10459 12291
rect 2881 12189 2915 12223
rect 4261 12189 4295 12223
rect 5181 12189 5215 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 10517 12189 10551 12223
rect 10701 12189 10735 12223
rect 11621 12189 11655 12223
rect 4905 12121 4939 12155
rect 8033 12121 8067 12155
rect 2421 12053 2455 12087
rect 3249 12053 3283 12087
rect 4813 12053 4847 12087
rect 11161 12053 11195 12087
rect 11529 12053 11563 12087
rect 13001 12053 13035 12087
rect 2513 11849 2547 11883
rect 5733 11849 5767 11883
rect 7021 11849 7055 11883
rect 10057 11849 10091 11883
rect 10977 11849 11011 11883
rect 12449 11849 12483 11883
rect 2237 11781 2271 11815
rect 4721 11781 4755 11815
rect 10701 11781 10735 11815
rect 12173 11781 12207 11815
rect 1593 11713 1627 11747
rect 3709 11713 3743 11747
rect 5181 11713 5215 11747
rect 5273 11713 5307 11747
rect 6653 11713 6687 11747
rect 7665 11713 7699 11747
rect 8677 11713 8711 11747
rect 11621 11713 11655 11747
rect 13093 11713 13127 11747
rect 1409 11645 1443 11679
rect 3617 11645 3651 11679
rect 4629 11645 4663 11679
rect 7389 11645 7423 11679
rect 8933 11645 8967 11679
rect 11345 11645 11379 11679
rect 3065 11577 3099 11611
rect 4261 11577 4295 11611
rect 5089 11577 5123 11611
rect 3157 11509 3191 11543
rect 3525 11509 3559 11543
rect 7481 11509 7515 11543
rect 8125 11509 8159 11543
rect 8493 11509 8527 11543
rect 11161 11509 11195 11543
rect 12817 11509 12851 11543
rect 12909 11509 12943 11543
rect 13461 11509 13495 11543
rect 1685 11305 1719 11339
rect 2053 11305 2087 11339
rect 3249 11305 3283 11339
rect 4997 11305 5031 11339
rect 5273 11305 5307 11339
rect 5457 11305 5491 11339
rect 5917 11305 5951 11339
rect 7481 11305 7515 11339
rect 8769 11305 8803 11339
rect 11069 11305 11103 11339
rect 12173 11305 12207 11339
rect 13185 11305 13219 11339
rect 9045 11237 9079 11271
rect 9505 11237 9539 11271
rect 11621 11237 11655 11271
rect 12633 11237 12667 11271
rect 5825 11169 5859 11203
rect 7849 11169 7883 11203
rect 9689 11169 9723 11203
rect 9956 11169 9990 11203
rect 12541 11169 12575 11203
rect 4629 11101 4663 11135
rect 6009 11101 6043 11135
rect 6745 11101 6779 11135
rect 7941 11101 7975 11135
rect 8033 11101 8067 11135
rect 12817 11101 12851 11135
rect 7113 11033 7147 11067
rect 5641 10761 5675 10795
rect 6469 10761 6503 10795
rect 8033 10761 8067 10795
rect 9781 10761 9815 10795
rect 10609 10761 10643 10795
rect 11805 10761 11839 10795
rect 12265 10761 12299 10795
rect 2973 10693 3007 10727
rect 4445 10693 4479 10727
rect 6101 10693 6135 10727
rect 1593 10625 1627 10659
rect 2881 10625 2915 10659
rect 3617 10625 3651 10659
rect 5089 10625 5123 10659
rect 8585 10625 8619 10659
rect 9045 10625 9079 10659
rect 10149 10625 10183 10659
rect 11253 10625 11287 10659
rect 12449 10625 12483 10659
rect 12909 10625 12943 10659
rect 1409 10557 1443 10591
rect 2513 10557 2547 10591
rect 3985 10557 4019 10591
rect 7941 10557 7975 10591
rect 8401 10557 8435 10591
rect 3341 10489 3375 10523
rect 4997 10489 5031 10523
rect 11069 10489 11103 10523
rect 3433 10421 3467 10455
rect 4537 10421 4571 10455
rect 4905 10421 4939 10455
rect 6837 10421 6871 10455
rect 7573 10421 7607 10455
rect 8493 10421 8527 10455
rect 10425 10421 10459 10455
rect 10977 10421 11011 10455
rect 3341 10217 3375 10251
rect 4445 10217 4479 10251
rect 4813 10217 4847 10251
rect 5549 10217 5583 10251
rect 6009 10217 6043 10251
rect 6469 10217 6503 10251
rect 8033 10217 8067 10251
rect 9045 10217 9079 10251
rect 9873 10217 9907 10251
rect 11529 10217 11563 10251
rect 6561 10149 6595 10183
rect 11989 10149 12023 10183
rect 2697 10081 2731 10115
rect 7757 10081 7791 10115
rect 8401 10081 8435 10115
rect 11897 10081 11931 10115
rect 2789 10013 2823 10047
rect 2881 10013 2915 10047
rect 4905 10013 4939 10047
rect 4997 10013 5031 10047
rect 6745 10013 6779 10047
rect 8493 10013 8527 10047
rect 8585 10013 8619 10047
rect 12081 10013 12115 10047
rect 6101 9945 6135 9979
rect 7389 9945 7423 9979
rect 1593 9877 1627 9911
rect 2053 9877 2087 9911
rect 2329 9877 2363 9911
rect 10609 9877 10643 9911
rect 1685 9673 1719 9707
rect 2053 9673 2087 9707
rect 6193 9673 6227 9707
rect 8677 9673 8711 9707
rect 11253 9673 11287 9707
rect 4261 9605 4295 9639
rect 5365 9605 5399 9639
rect 6469 9605 6503 9639
rect 7113 9605 7147 9639
rect 11621 9605 11655 9639
rect 2881 9537 2915 9571
rect 7849 9537 7883 9571
rect 8861 9537 8895 9571
rect 4905 9469 4939 9503
rect 5549 9469 5583 9503
rect 6653 9469 6687 9503
rect 7757 9469 7791 9503
rect 9321 9469 9355 9503
rect 10057 9469 10091 9503
rect 10333 9469 10367 9503
rect 3126 9401 3160 9435
rect 7665 9401 7699 9435
rect 8401 9401 8435 9435
rect 2329 9333 2363 9367
rect 2789 9333 2823 9367
rect 5181 9333 5215 9367
rect 7297 9333 7331 9367
rect 9873 9333 9907 9367
rect 11897 9333 11931 9367
rect 2881 9129 2915 9163
rect 3433 9129 3467 9163
rect 4353 9129 4387 9163
rect 5273 9129 5307 9163
rect 6745 9129 6779 9163
rect 7849 9129 7883 9163
rect 7297 9061 7331 9095
rect 1501 8993 1535 9027
rect 1768 8993 1802 9027
rect 5365 8993 5399 9027
rect 5632 8993 5666 9027
rect 8217 8993 8251 9027
rect 4813 8925 4847 8959
rect 8309 8925 8343 8959
rect 8493 8925 8527 8959
rect 7757 8857 7791 8891
rect 9505 8789 9539 8823
rect 2697 8585 2731 8619
rect 5641 8585 5675 8619
rect 6193 8585 6227 8619
rect 6653 8585 6687 8619
rect 8769 8585 8803 8619
rect 9229 8585 9263 8619
rect 1593 8449 1627 8483
rect 3249 8449 3283 8483
rect 4261 8449 4295 8483
rect 9873 8449 9907 8483
rect 10057 8449 10091 8483
rect 1409 8381 1443 8415
rect 2605 8381 2639 8415
rect 3065 8381 3099 8415
rect 6837 8381 6871 8415
rect 7093 8381 7127 8415
rect 2237 8313 2271 8347
rect 4169 8313 4203 8347
rect 4528 8313 4562 8347
rect 9781 8313 9815 8347
rect 3157 8245 3191 8279
rect 3709 8245 3743 8279
rect 8217 8245 8251 8279
rect 9413 8245 9447 8279
rect 10517 8245 10551 8279
rect 2421 8041 2455 8075
rect 4077 8041 4111 8075
rect 5181 8041 5215 8075
rect 5457 8041 5491 8075
rect 6561 8041 6595 8075
rect 7021 8041 7055 8075
rect 8493 8041 8527 8075
rect 10793 8041 10827 8075
rect 13093 8041 13127 8075
rect 2053 7973 2087 8007
rect 2789 7973 2823 8007
rect 1685 7905 1719 7939
rect 2881 7905 2915 7939
rect 4445 7905 4479 7939
rect 4537 7905 4571 7939
rect 7369 7905 7403 7939
rect 10057 7905 10091 7939
rect 11980 7905 12014 7939
rect 2973 7837 3007 7871
rect 4721 7837 4755 7871
rect 6193 7837 6227 7871
rect 7113 7837 7147 7871
rect 10149 7837 10183 7871
rect 10333 7837 10367 7871
rect 11713 7837 11747 7871
rect 9413 7769 9447 7803
rect 9137 7701 9171 7735
rect 9689 7701 9723 7735
rect 11529 7701 11563 7735
rect 1869 7497 1903 7531
rect 4077 7497 4111 7531
rect 5181 7497 5215 7531
rect 6653 7497 6687 7531
rect 7481 7497 7515 7531
rect 11253 7497 11287 7531
rect 11897 7497 11931 7531
rect 12173 7497 12207 7531
rect 12449 7497 12483 7531
rect 1777 7429 1811 7463
rect 9321 7429 9355 7463
rect 2329 7361 2363 7395
rect 2421 7361 2455 7395
rect 7941 7361 7975 7395
rect 8953 7361 8987 7395
rect 13001 7361 13035 7395
rect 2237 7293 2271 7327
rect 3341 7293 3375 7327
rect 3801 7293 3835 7327
rect 4905 7293 4939 7327
rect 6837 7293 6871 7327
rect 8217 7293 8251 7327
rect 8769 7293 8803 7327
rect 9873 7293 9907 7327
rect 10140 7225 10174 7259
rect 12909 7225 12943 7259
rect 13461 7225 13495 7259
rect 2973 7157 3007 7191
rect 4445 7157 4479 7191
rect 4721 7157 4755 7191
rect 7021 7157 7055 7191
rect 8033 7157 8067 7191
rect 8309 7157 8343 7191
rect 8677 7157 8711 7191
rect 9689 7157 9723 7191
rect 12817 7157 12851 7191
rect 13829 7157 13863 7191
rect 1961 6953 1995 6987
rect 2697 6953 2731 6987
rect 7205 6953 7239 6987
rect 7573 6953 7607 6987
rect 9137 6953 9171 6987
rect 9873 6953 9907 6987
rect 10241 6953 10275 6987
rect 12817 6953 12851 6987
rect 2053 6817 2087 6851
rect 5181 6817 5215 6851
rect 6285 6817 6319 6851
rect 7941 6817 7975 6851
rect 8401 6817 8435 6851
rect 10333 6817 10367 6851
rect 10977 6817 11011 6851
rect 11693 6817 11727 6851
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 10425 6749 10459 6783
rect 11437 6749 11471 6783
rect 9505 6681 9539 6715
rect 2237 6613 2271 6647
rect 5365 6613 5399 6647
rect 6469 6613 6503 6647
rect 8033 6613 8067 6647
rect 11253 6613 11287 6647
rect 1777 6409 1811 6443
rect 5181 6409 5215 6443
rect 6561 6409 6595 6443
rect 7573 6409 7607 6443
rect 9045 6409 9079 6443
rect 10057 6409 10091 6443
rect 10517 6409 10551 6443
rect 10793 6409 10827 6443
rect 11805 6409 11839 6443
rect 2053 6341 2087 6375
rect 3617 6341 3651 6375
rect 5825 6341 5859 6375
rect 6193 6341 6227 6375
rect 8585 6273 8619 6307
rect 9505 6273 9539 6307
rect 9597 6273 9631 6307
rect 11437 6273 11471 6307
rect 1869 6205 1903 6239
rect 2973 6205 3007 6239
rect 4445 6205 4479 6239
rect 4537 6205 4571 6239
rect 5641 6205 5675 6239
rect 7021 6205 7055 6239
rect 2513 6069 2547 6103
rect 3157 6069 3191 6103
rect 4721 6069 4755 6103
rect 7205 6069 7239 6103
rect 8125 6069 8159 6103
rect 8953 6069 8987 6103
rect 9413 6069 9447 6103
rect 11161 6069 11195 6103
rect 11253 6069 11287 6103
rect 12173 6069 12207 6103
rect 12449 6069 12483 6103
rect 6101 5865 6135 5899
rect 7573 5865 7607 5899
rect 7941 5865 7975 5899
rect 9505 5865 9539 5899
rect 10701 5865 10735 5899
rect 9137 5797 9171 5831
rect 2329 5729 2363 5763
rect 4077 5729 4111 5763
rect 6009 5729 6043 5763
rect 8401 5729 8435 5763
rect 10241 5729 10275 5763
rect 11897 5729 11931 5763
rect 6193 5661 6227 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 10793 5661 10827 5695
rect 10885 5661 10919 5695
rect 13001 5661 13035 5695
rect 4261 5593 4295 5627
rect 5641 5593 5675 5627
rect 11437 5593 11471 5627
rect 12541 5593 12575 5627
rect 2513 5525 2547 5559
rect 5549 5525 5583 5559
rect 6929 5525 6963 5559
rect 8033 5525 8067 5559
rect 10333 5525 10367 5559
rect 12081 5525 12115 5559
rect 12817 5525 12851 5559
rect 2881 5321 2915 5355
rect 4813 5321 4847 5355
rect 6101 5321 6135 5355
rect 11253 5321 11287 5355
rect 11989 5321 12023 5355
rect 12449 5321 12483 5355
rect 11621 5253 11655 5287
rect 2329 5185 2363 5219
rect 13093 5185 13127 5219
rect 2053 5117 2087 5151
rect 2145 5117 2179 5151
rect 3433 5117 3467 5151
rect 6837 5117 6871 5151
rect 9321 5117 9355 5151
rect 3341 5049 3375 5083
rect 3700 5049 3734 5083
rect 5733 5049 5767 5083
rect 6653 5049 6687 5083
rect 7082 5049 7116 5083
rect 8861 5049 8895 5083
rect 9229 5049 9263 5083
rect 9588 5049 9622 5083
rect 12909 5049 12943 5083
rect 8217 4981 8251 5015
rect 10701 4981 10735 5015
rect 12817 4981 12851 5015
rect 13461 4981 13495 5015
rect 2421 4777 2455 4811
rect 3525 4777 3559 4811
rect 4353 4777 4387 4811
rect 4813 4777 4847 4811
rect 7021 4777 7055 4811
rect 7849 4777 7883 4811
rect 9321 4777 9355 4811
rect 10701 4777 10735 4811
rect 11805 4777 11839 4811
rect 12265 4709 12299 4743
rect 2789 4641 2823 4675
rect 4997 4641 5031 4675
rect 5253 4641 5287 4675
rect 10609 4641 10643 4675
rect 11253 4641 11287 4675
rect 12173 4641 12207 4675
rect 12817 4641 12851 4675
rect 13369 4641 13403 4675
rect 2329 4573 2363 4607
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 10885 4573 10919 4607
rect 12449 4573 12483 4607
rect 6377 4505 6411 4539
rect 7481 4505 7515 4539
rect 8861 4505 8895 4539
rect 10241 4505 10275 4539
rect 13185 4505 13219 4539
rect 1685 4437 1719 4471
rect 7297 4437 7331 4471
rect 8493 4437 8527 4471
rect 9965 4437 9999 4471
rect 11713 4437 11747 4471
rect 13553 4437 13587 4471
rect 2513 4233 2547 4267
rect 4445 4233 4479 4267
rect 10425 4233 10459 4267
rect 10793 4233 10827 4267
rect 12081 4233 12115 4267
rect 12173 4233 12207 4267
rect 12449 4233 12483 4267
rect 13461 4233 13495 4267
rect 1593 4097 1627 4131
rect 6837 4097 6871 4131
rect 9137 4097 9171 4131
rect 9873 4097 9907 4131
rect 1409 4029 1443 4063
rect 3065 4029 3099 4063
rect 3332 4029 3366 4063
rect 5549 4029 5583 4063
rect 6193 4029 6227 4063
rect 7104 4029 7138 4063
rect 8769 4029 8803 4063
rect 9689 4029 9723 4063
rect 10885 4029 10919 4063
rect 11437 4029 11471 4063
rect 2973 3961 3007 3995
rect 5089 3961 5123 3995
rect 5457 3961 5491 3995
rect 6653 3961 6687 3995
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 5733 3893 5767 3927
rect 8217 3893 8251 3927
rect 9321 3893 9355 3927
rect 9781 3893 9815 3927
rect 11069 3893 11103 3927
rect 11897 3893 11931 3927
rect 12081 3893 12115 3927
rect 12817 3893 12851 3927
rect 1961 3689 1995 3723
rect 2421 3689 2455 3723
rect 3433 3689 3467 3723
rect 4537 3689 4571 3723
rect 5457 3689 5491 3723
rect 6561 3689 6595 3723
rect 7021 3689 7055 3723
rect 7941 3689 7975 3723
rect 9321 3689 9355 3723
rect 9873 3689 9907 3723
rect 10425 3689 10459 3723
rect 13001 3689 13035 3723
rect 4905 3621 4939 3655
rect 6009 3621 6043 3655
rect 6469 3621 6503 3655
rect 7665 3621 7699 3655
rect 8861 3621 8895 3655
rect 11529 3621 11563 3655
rect 11888 3621 11922 3655
rect 2329 3553 2363 3587
rect 2789 3553 2823 3587
rect 5365 3553 5399 3587
rect 6929 3553 6963 3587
rect 8125 3553 8159 3587
rect 1409 3485 1443 3519
rect 2881 3485 2915 3519
rect 3065 3485 3099 3519
rect 5549 3485 5583 3519
rect 7113 3485 7147 3519
rect 10517 3485 10551 3519
rect 10701 3485 10735 3519
rect 11069 3485 11103 3519
rect 11621 3485 11655 3519
rect 4997 3417 5031 3451
rect 10057 3417 10091 3451
rect 8309 3349 8343 3383
rect 1685 3145 1719 3179
rect 4905 3145 4939 3179
rect 6653 3145 6687 3179
rect 7021 3145 7055 3179
rect 7205 3145 7239 3179
rect 8309 3145 8343 3179
rect 8677 3145 8711 3179
rect 10149 3145 10183 3179
rect 10701 3145 10735 3179
rect 11161 3145 11195 3179
rect 11805 3145 11839 3179
rect 12449 3145 12483 3179
rect 4445 3077 4479 3111
rect 8125 3077 8159 3111
rect 11437 3077 11471 3111
rect 4813 3009 4847 3043
rect 5457 3009 5491 3043
rect 7849 3009 7883 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 2145 2941 2179 2975
rect 5273 2941 5307 2975
rect 7573 2941 7607 2975
rect 8125 2941 8159 2975
rect 8769 2941 8803 2975
rect 9025 2941 9059 2975
rect 11253 2941 11287 2975
rect 13829 2941 13863 2975
rect 1961 2873 1995 2907
rect 2390 2873 2424 2907
rect 5365 2873 5399 2907
rect 5917 2873 5951 2907
rect 7665 2873 7699 2907
rect 12265 2873 12299 2907
rect 12817 2873 12851 2907
rect 3525 2805 3559 2839
rect 13461 2805 13495 2839
rect 1685 2601 1719 2635
rect 2421 2601 2455 2635
rect 2789 2601 2823 2635
rect 4905 2601 4939 2635
rect 5365 2601 5399 2635
rect 6377 2601 6411 2635
rect 7941 2601 7975 2635
rect 8125 2601 8159 2635
rect 8585 2601 8619 2635
rect 11437 2601 11471 2635
rect 12633 2601 12667 2635
rect 13001 2601 13035 2635
rect 14013 2601 14047 2635
rect 4353 2533 4387 2567
rect 4813 2533 4847 2567
rect 6653 2533 6687 2567
rect 7665 2533 7699 2567
rect 9229 2533 9263 2567
rect 9597 2533 9631 2567
rect 10302 2533 10336 2567
rect 12081 2533 12115 2567
rect 1777 2465 1811 2499
rect 2881 2465 2915 2499
rect 5273 2465 5307 2499
rect 6929 2465 6963 2499
rect 8493 2465 8527 2499
rect 10057 2465 10091 2499
rect 12449 2465 12483 2499
rect 13093 2465 13127 2499
rect 3525 2397 3559 2431
rect 5457 2397 5491 2431
rect 5917 2397 5951 2431
rect 8769 2397 8803 2431
rect 13277 2397 13311 2431
rect 13645 2397 13679 2431
rect 1961 2329 1995 2363
rect 3065 2261 3099 2295
rect 7113 2261 7147 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 11606 36184 11612 36236
rect 11664 36224 11670 36236
rect 11773 36227 11831 36233
rect 11773 36224 11785 36227
rect 11664 36196 11785 36224
rect 11664 36184 11670 36196
rect 11773 36193 11785 36196
rect 11819 36193 11831 36227
rect 11773 36187 11831 36193
rect 11422 36116 11428 36168
rect 11480 36156 11486 36168
rect 11517 36159 11575 36165
rect 11517 36156 11529 36159
rect 11480 36128 11529 36156
rect 11480 36116 11486 36128
rect 11517 36125 11529 36128
rect 11563 36125 11575 36159
rect 11517 36119 11575 36125
rect 12434 35980 12440 36032
rect 12492 36020 12498 36032
rect 12897 36023 12955 36029
rect 12897 36020 12909 36023
rect 12492 35992 12909 36020
rect 12492 35980 12498 35992
rect 12897 35989 12909 35992
rect 12943 35989 12955 36023
rect 12897 35983 12955 35989
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 198 35776 204 35828
rect 256 35816 262 35828
rect 1302 35816 1308 35828
rect 256 35788 1308 35816
rect 256 35776 262 35788
rect 1302 35776 1308 35788
rect 1360 35776 1366 35828
rect 6914 35776 6920 35828
rect 6972 35816 6978 35828
rect 7377 35819 7435 35825
rect 7377 35816 7389 35819
rect 6972 35788 7389 35816
rect 6972 35776 6978 35788
rect 7377 35785 7389 35788
rect 7423 35785 7435 35819
rect 8478 35816 8484 35828
rect 8439 35788 8484 35816
rect 7377 35779 7435 35785
rect 8478 35776 8484 35788
rect 8536 35776 8542 35828
rect 11606 35816 11612 35828
rect 11567 35788 11612 35816
rect 11606 35776 11612 35788
rect 11664 35816 11670 35828
rect 11974 35816 11980 35828
rect 11664 35788 11980 35816
rect 11664 35776 11670 35788
rect 11974 35776 11980 35788
rect 12032 35776 12038 35828
rect 7193 35615 7251 35621
rect 7193 35581 7205 35615
rect 7239 35612 7251 35615
rect 8297 35615 8355 35621
rect 7239 35584 7880 35612
rect 7239 35581 7251 35584
rect 7193 35575 7251 35581
rect 7852 35485 7880 35584
rect 8297 35581 8309 35615
rect 8343 35612 8355 35615
rect 8849 35615 8907 35621
rect 8849 35612 8861 35615
rect 8343 35584 8861 35612
rect 8343 35581 8355 35584
rect 8297 35575 8355 35581
rect 8849 35581 8861 35584
rect 8895 35612 8907 35615
rect 10042 35612 10048 35624
rect 8895 35584 10048 35612
rect 8895 35581 8907 35584
rect 8849 35575 8907 35581
rect 10042 35572 10048 35584
rect 10100 35572 10106 35624
rect 11422 35504 11428 35556
rect 11480 35544 11486 35556
rect 11885 35547 11943 35553
rect 11885 35544 11897 35547
rect 11480 35516 11897 35544
rect 11480 35504 11486 35516
rect 11885 35513 11897 35516
rect 11931 35513 11943 35547
rect 11885 35507 11943 35513
rect 7837 35479 7895 35485
rect 7837 35445 7849 35479
rect 7883 35476 7895 35479
rect 8018 35476 8024 35488
rect 7883 35448 8024 35476
rect 7883 35445 7895 35448
rect 7837 35439 7895 35445
rect 8018 35436 8024 35448
rect 8076 35436 8082 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 1762 35232 1768 35284
rect 1820 35272 1826 35284
rect 2317 35275 2375 35281
rect 2317 35272 2329 35275
rect 1820 35244 2329 35272
rect 1820 35232 1826 35244
rect 2317 35241 2329 35244
rect 2363 35241 2375 35275
rect 2317 35235 2375 35241
rect 3970 35232 3976 35284
rect 4028 35272 4034 35284
rect 4249 35275 4307 35281
rect 4249 35272 4261 35275
rect 4028 35244 4261 35272
rect 4028 35232 4034 35244
rect 4249 35241 4261 35244
rect 4295 35241 4307 35275
rect 4249 35235 4307 35241
rect 5353 35275 5411 35281
rect 5353 35241 5365 35275
rect 5399 35272 5411 35275
rect 5442 35272 5448 35284
rect 5399 35244 5448 35272
rect 5399 35241 5411 35244
rect 5353 35235 5411 35241
rect 5442 35232 5448 35244
rect 5500 35232 5506 35284
rect 7374 35232 7380 35284
rect 7432 35272 7438 35284
rect 7653 35275 7711 35281
rect 7653 35272 7665 35275
rect 7432 35244 7665 35272
rect 7432 35232 7438 35244
rect 7653 35241 7665 35244
rect 7699 35241 7711 35275
rect 7653 35235 7711 35241
rect 9858 35164 9864 35216
rect 9916 35213 9922 35216
rect 9916 35207 9980 35213
rect 9916 35173 9934 35207
rect 9968 35173 9980 35207
rect 9916 35167 9980 35173
rect 9916 35164 9922 35167
rect 2133 35139 2191 35145
rect 2133 35105 2145 35139
rect 2179 35136 2191 35139
rect 2406 35136 2412 35148
rect 2179 35108 2412 35136
rect 2179 35105 2191 35108
rect 2133 35099 2191 35105
rect 2406 35096 2412 35108
rect 2464 35096 2470 35148
rect 4062 35136 4068 35148
rect 4023 35108 4068 35136
rect 4062 35096 4068 35108
rect 4120 35096 4126 35148
rect 5166 35136 5172 35148
rect 5127 35108 5172 35136
rect 5166 35096 5172 35108
rect 5224 35096 5230 35148
rect 6365 35139 6423 35145
rect 6365 35105 6377 35139
rect 6411 35136 6423 35139
rect 6730 35136 6736 35148
rect 6411 35108 6736 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 6730 35096 6736 35108
rect 6788 35096 6794 35148
rect 7466 35136 7472 35148
rect 7427 35108 7472 35136
rect 7466 35096 7472 35108
rect 7524 35096 7530 35148
rect 9677 35139 9735 35145
rect 9677 35105 9689 35139
rect 9723 35136 9735 35139
rect 11422 35136 11428 35148
rect 9723 35108 11428 35136
rect 9723 35105 9735 35108
rect 9677 35099 9735 35105
rect 11422 35096 11428 35108
rect 11480 35096 11486 35148
rect 4154 34960 4160 35012
rect 4212 35000 4218 35012
rect 6549 35003 6607 35009
rect 6549 35000 6561 35003
rect 4212 34972 6561 35000
rect 4212 34960 4218 34972
rect 6549 34969 6561 34972
rect 6595 34969 6607 35003
rect 6549 34963 6607 34969
rect 5718 34932 5724 34944
rect 5679 34904 5724 34932
rect 5718 34892 5724 34904
rect 5776 34892 5782 34944
rect 8110 34932 8116 34944
rect 8071 34904 8116 34932
rect 8110 34892 8116 34904
rect 8168 34892 8174 34944
rect 11057 34935 11115 34941
rect 11057 34901 11069 34935
rect 11103 34932 11115 34935
rect 11146 34932 11152 34944
rect 11103 34904 11152 34932
rect 11103 34901 11115 34904
rect 11057 34895 11115 34901
rect 11146 34892 11152 34904
rect 11204 34892 11210 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 566 34688 572 34740
rect 624 34728 630 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 624 34700 1593 34728
rect 624 34688 630 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 2038 34728 2044 34740
rect 1999 34700 2044 34728
rect 1581 34691 1639 34697
rect 2038 34688 2044 34700
rect 2096 34688 2102 34740
rect 2590 34688 2596 34740
rect 2648 34728 2654 34740
rect 3789 34731 3847 34737
rect 3789 34728 3801 34731
rect 2648 34700 3801 34728
rect 2648 34688 2654 34700
rect 3789 34697 3801 34700
rect 3835 34697 3847 34731
rect 3789 34691 3847 34697
rect 5721 34731 5779 34737
rect 5721 34697 5733 34731
rect 5767 34728 5779 34731
rect 6178 34728 6184 34740
rect 5767 34700 6184 34728
rect 5767 34697 5779 34700
rect 5721 34691 5779 34697
rect 6178 34688 6184 34700
rect 6236 34688 6242 34740
rect 6638 34688 6644 34740
rect 6696 34728 6702 34740
rect 7009 34731 7067 34737
rect 7009 34728 7021 34731
rect 6696 34700 7021 34728
rect 6696 34688 6702 34700
rect 7009 34697 7021 34700
rect 7055 34697 7067 34731
rect 7009 34691 7067 34697
rect 7466 34688 7472 34740
rect 7524 34728 7530 34740
rect 7745 34731 7803 34737
rect 7745 34728 7757 34731
rect 7524 34700 7757 34728
rect 7524 34688 7530 34700
rect 7745 34697 7757 34700
rect 7791 34697 7803 34731
rect 7745 34691 7803 34697
rect 8294 34688 8300 34740
rect 8352 34728 8358 34740
rect 9401 34731 9459 34737
rect 9401 34728 9413 34731
rect 8352 34700 9413 34728
rect 8352 34688 8358 34700
rect 9401 34697 9413 34700
rect 9447 34728 9459 34731
rect 9858 34728 9864 34740
rect 9447 34700 9864 34728
rect 9447 34697 9459 34700
rect 9401 34691 9459 34697
rect 9858 34688 9864 34700
rect 9916 34688 9922 34740
rect 10318 34728 10324 34740
rect 10279 34700 10324 34728
rect 10318 34688 10324 34700
rect 10376 34728 10382 34740
rect 13630 34728 13636 34740
rect 10376 34700 11008 34728
rect 13591 34700 13636 34728
rect 10376 34688 10382 34700
rect 1394 34620 1400 34672
rect 1452 34660 1458 34672
rect 2685 34663 2743 34669
rect 2685 34660 2697 34663
rect 1452 34632 2697 34660
rect 1452 34620 1458 34632
rect 2685 34629 2697 34632
rect 2731 34629 2743 34663
rect 2685 34623 2743 34629
rect 4249 34663 4307 34669
rect 4249 34629 4261 34663
rect 4295 34660 4307 34663
rect 4890 34660 4896 34672
rect 4295 34632 4896 34660
rect 4295 34629 4307 34632
rect 4249 34623 4307 34629
rect 2406 34592 2412 34604
rect 2319 34564 2412 34592
rect 2406 34552 2412 34564
rect 2464 34592 2470 34604
rect 2590 34592 2596 34604
rect 2464 34564 2596 34592
rect 2464 34552 2470 34564
rect 2590 34552 2596 34564
rect 2648 34552 2654 34604
rect 3326 34552 3332 34604
rect 3384 34592 3390 34604
rect 4154 34592 4160 34604
rect 3384 34564 4160 34592
rect 3384 34552 3390 34564
rect 4154 34552 4160 34564
rect 4212 34552 4218 34604
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 2038 34524 2044 34536
rect 1443 34496 2044 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2501 34527 2559 34533
rect 2501 34493 2513 34527
rect 2547 34524 2559 34527
rect 3145 34527 3203 34533
rect 3145 34524 3157 34527
rect 2547 34496 3157 34524
rect 2547 34493 2559 34496
rect 2501 34487 2559 34493
rect 3145 34493 3157 34496
rect 3191 34524 3203 34527
rect 3234 34524 3240 34536
rect 3191 34496 3240 34524
rect 3191 34493 3203 34496
rect 3145 34487 3203 34493
rect 3234 34484 3240 34496
rect 3292 34484 3298 34536
rect 3605 34527 3663 34533
rect 3605 34493 3617 34527
rect 3651 34524 3663 34527
rect 4264 34524 4292 34623
rect 4890 34620 4896 34632
rect 4948 34620 4954 34672
rect 10980 34601 11008 34700
rect 13630 34688 13636 34700
rect 13688 34688 13694 34740
rect 10965 34595 11023 34601
rect 10965 34561 10977 34595
rect 11011 34561 11023 34595
rect 11146 34592 11152 34604
rect 11107 34564 11152 34592
rect 10965 34555 11023 34561
rect 11146 34552 11152 34564
rect 11204 34592 11210 34604
rect 11517 34595 11575 34601
rect 11517 34592 11529 34595
rect 11204 34564 11529 34592
rect 11204 34552 11210 34564
rect 11517 34561 11529 34564
rect 11563 34561 11575 34595
rect 11517 34555 11575 34561
rect 3651 34496 4292 34524
rect 5537 34527 5595 34533
rect 3651 34493 3663 34496
rect 3605 34487 3663 34493
rect 5537 34493 5549 34527
rect 5583 34524 5595 34527
rect 5718 34524 5724 34536
rect 5583 34496 5724 34524
rect 5583 34493 5595 34496
rect 5537 34487 5595 34493
rect 5718 34484 5724 34496
rect 5776 34484 5782 34536
rect 6457 34527 6515 34533
rect 6457 34493 6469 34527
rect 6503 34524 6515 34527
rect 6730 34524 6736 34536
rect 6503 34496 6736 34524
rect 6503 34493 6515 34496
rect 6457 34487 6515 34493
rect 6730 34484 6736 34496
rect 6788 34484 6794 34536
rect 6825 34527 6883 34533
rect 6825 34493 6837 34527
rect 6871 34524 6883 34527
rect 7190 34524 7196 34536
rect 6871 34496 7196 34524
rect 6871 34493 6883 34496
rect 6825 34487 6883 34493
rect 7190 34484 7196 34496
rect 7248 34524 7254 34536
rect 7377 34527 7435 34533
rect 7377 34524 7389 34527
rect 7248 34496 7389 34524
rect 7248 34484 7254 34496
rect 7377 34493 7389 34496
rect 7423 34493 7435 34527
rect 7377 34487 7435 34493
rect 7926 34484 7932 34536
rect 7984 34524 7990 34536
rect 8021 34527 8079 34533
rect 8021 34524 8033 34527
rect 7984 34496 8033 34524
rect 7984 34484 7990 34496
rect 8021 34493 8033 34496
rect 8067 34493 8079 34527
rect 9950 34524 9956 34536
rect 9911 34496 9956 34524
rect 8021 34487 8079 34493
rect 9950 34484 9956 34496
rect 10008 34524 10014 34536
rect 10873 34527 10931 34533
rect 10873 34524 10885 34527
rect 10008 34496 10885 34524
rect 10008 34484 10014 34496
rect 10873 34493 10885 34496
rect 10919 34493 10931 34527
rect 13446 34524 13452 34536
rect 13407 34496 13452 34524
rect 10873 34487 10931 34493
rect 13446 34484 13452 34496
rect 13504 34524 13510 34536
rect 14001 34527 14059 34533
rect 14001 34524 14013 34527
rect 13504 34496 14013 34524
rect 13504 34484 13510 34496
rect 14001 34493 14013 34496
rect 14047 34493 14059 34527
rect 14001 34487 14059 34493
rect 4338 34416 4344 34468
rect 4396 34456 4402 34468
rect 5166 34456 5172 34468
rect 4396 34428 5172 34456
rect 4396 34416 4402 34428
rect 5166 34416 5172 34428
rect 5224 34416 5230 34468
rect 8110 34416 8116 34468
rect 8168 34456 8174 34468
rect 8288 34459 8346 34465
rect 8288 34456 8300 34459
rect 8168 34428 8300 34456
rect 8168 34416 8174 34428
rect 8288 34425 8300 34428
rect 8334 34456 8346 34459
rect 8570 34456 8576 34468
rect 8334 34428 8576 34456
rect 8334 34425 8346 34428
rect 8288 34419 8346 34425
rect 8570 34416 8576 34428
rect 8628 34416 8634 34468
rect 4062 34348 4068 34400
rect 4120 34388 4126 34400
rect 4617 34391 4675 34397
rect 4617 34388 4629 34391
rect 4120 34360 4629 34388
rect 4120 34348 4126 34360
rect 4617 34357 4629 34360
rect 4663 34388 4675 34391
rect 5258 34388 5264 34400
rect 4663 34360 5264 34388
rect 4663 34357 4675 34360
rect 4617 34351 4675 34357
rect 5258 34348 5264 34360
rect 5316 34348 5322 34400
rect 10502 34388 10508 34400
rect 10463 34360 10508 34388
rect 10502 34348 10508 34360
rect 10560 34348 10566 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1394 34144 1400 34196
rect 1452 34184 1458 34196
rect 1581 34187 1639 34193
rect 1581 34184 1593 34187
rect 1452 34156 1593 34184
rect 1452 34144 1458 34156
rect 1581 34153 1593 34156
rect 1627 34153 1639 34187
rect 1581 34147 1639 34153
rect 2130 34144 2136 34196
rect 2188 34184 2194 34196
rect 2685 34187 2743 34193
rect 2685 34184 2697 34187
rect 2188 34156 2697 34184
rect 2188 34144 2194 34156
rect 2685 34153 2697 34156
rect 2731 34153 2743 34187
rect 2685 34147 2743 34153
rect 4154 34144 4160 34196
rect 4212 34184 4218 34196
rect 4249 34187 4307 34193
rect 4249 34184 4261 34187
rect 4212 34156 4261 34184
rect 4212 34144 4218 34156
rect 4249 34153 4261 34156
rect 4295 34153 4307 34187
rect 4249 34147 4307 34153
rect 4982 34144 4988 34196
rect 5040 34184 5046 34196
rect 5445 34187 5503 34193
rect 5445 34184 5457 34187
rect 5040 34156 5457 34184
rect 5040 34144 5046 34156
rect 5445 34153 5457 34156
rect 5491 34153 5503 34187
rect 6914 34184 6920 34196
rect 6875 34156 6920 34184
rect 5445 34147 5503 34153
rect 6914 34144 6920 34156
rect 6972 34144 6978 34196
rect 7742 34144 7748 34196
rect 7800 34184 7806 34196
rect 8021 34187 8079 34193
rect 8021 34184 8033 34187
rect 7800 34156 8033 34184
rect 7800 34144 7806 34156
rect 8021 34153 8033 34156
rect 8067 34153 8079 34187
rect 9858 34184 9864 34196
rect 9819 34156 9864 34184
rect 8021 34147 8079 34153
rect 9858 34144 9864 34156
rect 9916 34144 9922 34196
rect 11885 34187 11943 34193
rect 11885 34153 11897 34187
rect 11931 34184 11943 34187
rect 11974 34184 11980 34196
rect 11931 34156 11980 34184
rect 11931 34153 11943 34156
rect 11885 34147 11943 34153
rect 11974 34144 11980 34156
rect 12032 34144 12038 34196
rect 1397 34051 1455 34057
rect 1397 34017 1409 34051
rect 1443 34048 1455 34051
rect 1946 34048 1952 34060
rect 1443 34020 1952 34048
rect 1443 34017 1455 34020
rect 1397 34011 1455 34017
rect 1946 34008 1952 34020
rect 2004 34008 2010 34060
rect 2501 34051 2559 34057
rect 2501 34017 2513 34051
rect 2547 34048 2559 34051
rect 3326 34048 3332 34060
rect 2547 34020 3332 34048
rect 2547 34017 2559 34020
rect 2501 34011 2559 34017
rect 3326 34008 3332 34020
rect 3384 34008 3390 34060
rect 4062 34048 4068 34060
rect 4023 34020 4068 34048
rect 4062 34008 4068 34020
rect 4120 34008 4126 34060
rect 5261 34051 5319 34057
rect 5261 34017 5273 34051
rect 5307 34048 5319 34051
rect 5442 34048 5448 34060
rect 5307 34020 5448 34048
rect 5307 34017 5319 34020
rect 5261 34011 5319 34017
rect 5442 34008 5448 34020
rect 5500 34008 5506 34060
rect 6638 34008 6644 34060
rect 6696 34048 6702 34060
rect 6733 34051 6791 34057
rect 6733 34048 6745 34051
rect 6696 34020 6745 34048
rect 6696 34008 6702 34020
rect 6733 34017 6745 34020
rect 6779 34017 6791 34051
rect 6733 34011 6791 34017
rect 7558 34008 7564 34060
rect 7616 34048 7622 34060
rect 7837 34051 7895 34057
rect 7837 34048 7849 34051
rect 7616 34020 7849 34048
rect 7616 34008 7622 34020
rect 7837 34017 7849 34020
rect 7883 34017 7895 34051
rect 7837 34011 7895 34017
rect 10772 34051 10830 34057
rect 10772 34017 10784 34051
rect 10818 34048 10830 34051
rect 11146 34048 11152 34060
rect 10818 34020 11152 34048
rect 10818 34017 10830 34020
rect 10772 34011 10830 34017
rect 11146 34008 11152 34020
rect 11204 34008 11210 34060
rect 10505 33983 10563 33989
rect 10505 33949 10517 33983
rect 10551 33949 10563 33983
rect 10505 33943 10563 33949
rect 6822 33804 6828 33856
rect 6880 33844 6886 33856
rect 7377 33847 7435 33853
rect 7377 33844 7389 33847
rect 6880 33816 7389 33844
rect 6880 33804 6886 33816
rect 7377 33813 7389 33816
rect 7423 33844 7435 33847
rect 7926 33844 7932 33856
rect 7423 33816 7932 33844
rect 7423 33813 7435 33816
rect 7377 33807 7435 33813
rect 7926 33804 7932 33816
rect 7984 33844 7990 33856
rect 8294 33844 8300 33856
rect 7984 33816 8300 33844
rect 7984 33804 7990 33816
rect 8294 33804 8300 33816
rect 8352 33844 8358 33856
rect 8389 33847 8447 33853
rect 8389 33844 8401 33847
rect 8352 33816 8401 33844
rect 8352 33804 8358 33816
rect 8389 33813 8401 33816
rect 8435 33813 8447 33847
rect 8389 33807 8447 33813
rect 10321 33847 10379 33853
rect 10321 33813 10333 33847
rect 10367 33844 10379 33847
rect 10520 33844 10548 33943
rect 11422 33844 11428 33856
rect 10367 33816 11428 33844
rect 10367 33813 10379 33816
rect 10321 33807 10379 33813
rect 11422 33804 11428 33816
rect 11480 33804 11486 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 934 33600 940 33652
rect 992 33640 998 33652
rect 1581 33643 1639 33649
rect 1581 33640 1593 33643
rect 992 33612 1593 33640
rect 992 33600 998 33612
rect 1581 33609 1593 33612
rect 1627 33609 1639 33643
rect 1946 33640 1952 33652
rect 1907 33612 1952 33640
rect 1581 33603 1639 33609
rect 1946 33600 1952 33612
rect 2004 33600 2010 33652
rect 2958 33640 2964 33652
rect 2919 33612 2964 33640
rect 2958 33600 2964 33612
rect 3016 33600 3022 33652
rect 11146 33640 11152 33652
rect 11107 33612 11152 33640
rect 11146 33600 11152 33612
rect 11204 33600 11210 33652
rect 6822 33504 6828 33516
rect 6783 33476 6828 33504
rect 6822 33464 6828 33476
rect 6880 33464 6886 33516
rect 9677 33507 9735 33513
rect 9677 33473 9689 33507
rect 9723 33504 9735 33507
rect 10502 33504 10508 33516
rect 9723 33476 10508 33504
rect 9723 33473 9735 33476
rect 9677 33467 9735 33473
rect 10502 33464 10508 33476
rect 10560 33504 10566 33516
rect 10597 33507 10655 33513
rect 10597 33504 10609 33507
rect 10560 33476 10609 33504
rect 10560 33464 10566 33476
rect 10597 33473 10609 33476
rect 10643 33473 10655 33507
rect 10778 33504 10784 33516
rect 10691 33476 10784 33504
rect 10597 33467 10655 33473
rect 10778 33464 10784 33476
rect 10836 33504 10842 33516
rect 11974 33504 11980 33516
rect 10836 33476 11980 33504
rect 10836 33464 10842 33476
rect 11974 33464 11980 33476
rect 12032 33464 12038 33516
rect 1397 33439 1455 33445
rect 1397 33405 1409 33439
rect 1443 33436 1455 33439
rect 2774 33436 2780 33448
rect 1443 33408 2452 33436
rect 2735 33408 2780 33436
rect 1443 33405 1455 33408
rect 1397 33399 1455 33405
rect 2424 33312 2452 33408
rect 2774 33396 2780 33408
rect 2832 33396 2838 33448
rect 6273 33371 6331 33377
rect 6273 33337 6285 33371
rect 6319 33368 6331 33371
rect 7092 33371 7150 33377
rect 7092 33368 7104 33371
rect 6319 33340 7104 33368
rect 6319 33337 6331 33340
rect 6273 33331 6331 33337
rect 7092 33337 7104 33340
rect 7138 33368 7150 33371
rect 7374 33368 7380 33380
rect 7138 33340 7380 33368
rect 7138 33337 7150 33340
rect 7092 33331 7150 33337
rect 7374 33328 7380 33340
rect 7432 33328 7438 33380
rect 9858 33328 9864 33380
rect 9916 33368 9922 33380
rect 10045 33371 10103 33377
rect 10045 33368 10057 33371
rect 9916 33340 10057 33368
rect 9916 33328 9922 33340
rect 10045 33337 10057 33340
rect 10091 33368 10103 33371
rect 10505 33371 10563 33377
rect 10505 33368 10517 33371
rect 10091 33340 10517 33368
rect 10091 33337 10103 33340
rect 10045 33331 10103 33337
rect 10505 33337 10517 33340
rect 10551 33337 10563 33371
rect 10505 33331 10563 33337
rect 2406 33300 2412 33312
rect 2367 33272 2412 33300
rect 2406 33260 2412 33272
rect 2464 33260 2470 33312
rect 3326 33300 3332 33312
rect 3287 33272 3332 33300
rect 3326 33260 3332 33272
rect 3384 33260 3390 33312
rect 4062 33260 4068 33312
rect 4120 33300 4126 33312
rect 4157 33303 4215 33309
rect 4157 33300 4169 33303
rect 4120 33272 4169 33300
rect 4120 33260 4126 33272
rect 4157 33269 4169 33272
rect 4203 33300 4215 33303
rect 4706 33300 4712 33312
rect 4203 33272 4712 33300
rect 4203 33269 4215 33272
rect 4157 33263 4215 33269
rect 4706 33260 4712 33272
rect 4764 33260 4770 33312
rect 5353 33303 5411 33309
rect 5353 33269 5365 33303
rect 5399 33300 5411 33303
rect 5442 33300 5448 33312
rect 5399 33272 5448 33300
rect 5399 33269 5411 33272
rect 5353 33263 5411 33269
rect 5442 33260 5448 33272
rect 5500 33260 5506 33312
rect 6638 33300 6644 33312
rect 6551 33272 6644 33300
rect 6638 33260 6644 33272
rect 6696 33300 6702 33312
rect 7282 33300 7288 33312
rect 6696 33272 7288 33300
rect 6696 33260 6702 33272
rect 7282 33260 7288 33272
rect 7340 33260 7346 33312
rect 8202 33300 8208 33312
rect 8163 33272 8208 33300
rect 8202 33260 8208 33272
rect 8260 33260 8266 33312
rect 10134 33300 10140 33312
rect 10095 33272 10140 33300
rect 10134 33260 10140 33272
rect 10192 33260 10198 33312
rect 11422 33260 11428 33312
rect 11480 33300 11486 33312
rect 11517 33303 11575 33309
rect 11517 33300 11529 33303
rect 11480 33272 11529 33300
rect 11480 33260 11486 33272
rect 11517 33269 11529 33272
rect 11563 33269 11575 33303
rect 11517 33263 11575 33269
rect 12250 33260 12256 33312
rect 12308 33300 12314 33312
rect 12437 33303 12495 33309
rect 12437 33300 12449 33303
rect 12308 33272 12449 33300
rect 12308 33260 12314 33272
rect 12437 33269 12449 33272
rect 12483 33269 12495 33303
rect 12437 33263 12495 33269
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 2774 33096 2780 33108
rect 2735 33068 2780 33096
rect 2774 33056 2780 33068
rect 2832 33056 2838 33108
rect 6822 33096 6828 33108
rect 6783 33068 6828 33096
rect 6822 33056 6828 33068
rect 6880 33056 6886 33108
rect 7558 33056 7564 33108
rect 7616 33096 7622 33108
rect 7837 33099 7895 33105
rect 7837 33096 7849 33099
rect 7616 33068 7849 33096
rect 7616 33056 7622 33068
rect 7837 33065 7849 33068
rect 7883 33065 7895 33099
rect 7837 33059 7895 33065
rect 10229 33099 10287 33105
rect 10229 33065 10241 33099
rect 10275 33096 10287 33099
rect 10778 33096 10784 33108
rect 10275 33068 10784 33096
rect 10275 33065 10287 33068
rect 10229 33059 10287 33065
rect 10778 33056 10784 33068
rect 10836 33056 10842 33108
rect 1486 32988 1492 33040
rect 1544 33028 1550 33040
rect 1673 33031 1731 33037
rect 1673 33028 1685 33031
rect 1544 33000 1685 33028
rect 1544 32988 1550 33000
rect 1673 32997 1685 33000
rect 1719 32997 1731 33031
rect 1673 32991 1731 32997
rect 11793 33031 11851 33037
rect 11793 32997 11805 33031
rect 11839 33028 11851 33031
rect 12250 33028 12256 33040
rect 11839 33000 12256 33028
rect 11839 32997 11851 33000
rect 11793 32991 11851 32997
rect 12250 32988 12256 33000
rect 12308 32988 12314 33040
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32960 1455 32963
rect 1762 32960 1768 32972
rect 1443 32932 1768 32960
rect 1443 32929 1455 32932
rect 1397 32923 1455 32929
rect 1762 32920 1768 32932
rect 1820 32920 1826 32972
rect 5810 32920 5816 32972
rect 5868 32960 5874 32972
rect 6917 32963 6975 32969
rect 6917 32960 6929 32963
rect 5868 32932 6929 32960
rect 5868 32920 5874 32932
rect 6917 32929 6929 32932
rect 6963 32929 6975 32963
rect 8386 32960 8392 32972
rect 8347 32932 8392 32960
rect 6917 32923 6975 32929
rect 8386 32920 8392 32932
rect 8444 32920 8450 32972
rect 9493 32963 9551 32969
rect 9493 32929 9505 32963
rect 9539 32960 9551 32963
rect 10502 32960 10508 32972
rect 9539 32932 10508 32960
rect 9539 32929 9551 32932
rect 9493 32923 9551 32929
rect 10502 32920 10508 32932
rect 10560 32960 10566 32972
rect 10689 32963 10747 32969
rect 10689 32960 10701 32963
rect 10560 32932 10701 32960
rect 10560 32920 10566 32932
rect 10689 32929 10701 32932
rect 10735 32929 10747 32963
rect 10689 32923 10747 32929
rect 12345 32963 12403 32969
rect 12345 32929 12357 32963
rect 12391 32960 12403 32963
rect 13538 32960 13544 32972
rect 12391 32932 13544 32960
rect 12391 32929 12403 32932
rect 12345 32923 12403 32929
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 7101 32895 7159 32901
rect 7101 32861 7113 32895
rect 7147 32892 7159 32895
rect 7374 32892 7380 32904
rect 7147 32864 7380 32892
rect 7147 32861 7159 32864
rect 7101 32855 7159 32861
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 7561 32895 7619 32901
rect 7561 32861 7573 32895
rect 7607 32892 7619 32895
rect 8478 32892 8484 32904
rect 7607 32864 8484 32892
rect 7607 32861 7619 32864
rect 7561 32855 7619 32861
rect 8478 32852 8484 32864
rect 8536 32852 8542 32904
rect 8570 32852 8576 32904
rect 8628 32892 8634 32904
rect 8628 32864 8673 32892
rect 8628 32852 8634 32864
rect 10134 32852 10140 32904
rect 10192 32892 10198 32904
rect 10781 32895 10839 32901
rect 10781 32892 10793 32895
rect 10192 32864 10793 32892
rect 10192 32852 10198 32864
rect 10781 32861 10793 32864
rect 10827 32861 10839 32895
rect 10781 32855 10839 32861
rect 10965 32895 11023 32901
rect 10965 32861 10977 32895
rect 11011 32892 11023 32895
rect 11146 32892 11152 32904
rect 11011 32864 11152 32892
rect 11011 32861 11023 32864
rect 10965 32855 11023 32861
rect 11146 32852 11152 32864
rect 11204 32892 11210 32904
rect 12250 32892 12256 32904
rect 11204 32864 12256 32892
rect 11204 32852 11210 32864
rect 12250 32852 12256 32864
rect 12308 32852 12314 32904
rect 12529 32895 12587 32901
rect 12529 32861 12541 32895
rect 12575 32892 12587 32895
rect 12575 32864 13032 32892
rect 12575 32861 12587 32864
rect 12529 32855 12587 32861
rect 12066 32784 12072 32836
rect 12124 32824 12130 32836
rect 12544 32824 12572 32855
rect 12124 32796 12572 32824
rect 12124 32784 12130 32796
rect 6457 32759 6515 32765
rect 6457 32725 6469 32759
rect 6503 32756 6515 32759
rect 7006 32756 7012 32768
rect 6503 32728 7012 32756
rect 6503 32725 6515 32728
rect 6457 32719 6515 32725
rect 7006 32716 7012 32728
rect 7064 32716 7070 32768
rect 7926 32716 7932 32768
rect 7984 32756 7990 32768
rect 8021 32759 8079 32765
rect 8021 32756 8033 32759
rect 7984 32728 8033 32756
rect 7984 32716 7990 32728
rect 8021 32725 8033 32728
rect 8067 32725 8079 32759
rect 8021 32719 8079 32725
rect 9125 32759 9183 32765
rect 9125 32725 9137 32759
rect 9171 32756 9183 32759
rect 9398 32756 9404 32768
rect 9171 32728 9404 32756
rect 9171 32725 9183 32728
rect 9125 32719 9183 32725
rect 9398 32716 9404 32728
rect 9456 32716 9462 32768
rect 10318 32756 10324 32768
rect 10279 32728 10324 32756
rect 10318 32716 10324 32728
rect 10376 32716 10382 32768
rect 11885 32759 11943 32765
rect 11885 32725 11897 32759
rect 11931 32756 11943 32759
rect 11974 32756 11980 32768
rect 11931 32728 11980 32756
rect 11931 32725 11943 32728
rect 11885 32719 11943 32725
rect 11974 32716 11980 32728
rect 12032 32716 12038 32768
rect 13004 32765 13032 32864
rect 12989 32759 13047 32765
rect 12989 32725 13001 32759
rect 13035 32756 13047 32759
rect 13078 32756 13084 32768
rect 13035 32728 13084 32756
rect 13035 32725 13047 32728
rect 12989 32719 13047 32725
rect 13078 32716 13084 32728
rect 13136 32716 13142 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 6181 32555 6239 32561
rect 6181 32521 6193 32555
rect 6227 32552 6239 32555
rect 6822 32552 6828 32564
rect 6227 32524 6828 32552
rect 6227 32521 6239 32524
rect 6181 32515 6239 32521
rect 6822 32512 6828 32524
rect 6880 32512 6886 32564
rect 8478 32512 8484 32564
rect 8536 32552 8542 32564
rect 8849 32555 8907 32561
rect 8849 32552 8861 32555
rect 8536 32524 8861 32552
rect 8536 32512 8542 32524
rect 8849 32521 8861 32524
rect 8895 32521 8907 32555
rect 8849 32515 8907 32521
rect 9674 32512 9680 32564
rect 9732 32552 9738 32564
rect 9953 32555 10011 32561
rect 9953 32552 9965 32555
rect 9732 32524 9965 32552
rect 9732 32512 9738 32524
rect 9953 32521 9965 32524
rect 9999 32521 10011 32555
rect 10502 32552 10508 32564
rect 10463 32524 10508 32552
rect 9953 32515 10011 32521
rect 5810 32444 5816 32496
rect 5868 32484 5874 32496
rect 6457 32487 6515 32493
rect 6457 32484 6469 32487
rect 5868 32456 6469 32484
rect 5868 32444 5874 32456
rect 6457 32453 6469 32456
rect 6503 32453 6515 32487
rect 8662 32484 8668 32496
rect 8623 32456 8668 32484
rect 6457 32447 6515 32453
rect 8662 32444 8668 32456
rect 8720 32444 8726 32496
rect 7374 32376 7380 32428
rect 7432 32416 7438 32428
rect 7469 32419 7527 32425
rect 7469 32416 7481 32419
rect 7432 32388 7481 32416
rect 7432 32376 7438 32388
rect 7469 32385 7481 32388
rect 7515 32416 7527 32419
rect 7834 32416 7840 32428
rect 7515 32388 7840 32416
rect 7515 32385 7527 32388
rect 7469 32379 7527 32385
rect 7834 32376 7840 32388
rect 7892 32376 7898 32428
rect 3513 32351 3571 32357
rect 3513 32317 3525 32351
rect 3559 32348 3571 32351
rect 3970 32348 3976 32360
rect 3559 32320 3976 32348
rect 3559 32317 3571 32320
rect 3513 32311 3571 32317
rect 3970 32308 3976 32320
rect 4028 32308 4034 32360
rect 6914 32308 6920 32360
rect 6972 32348 6978 32360
rect 7285 32351 7343 32357
rect 7285 32348 7297 32351
rect 6972 32320 7297 32348
rect 6972 32308 6978 32320
rect 7285 32317 7297 32320
rect 7331 32317 7343 32351
rect 8680 32348 8708 32444
rect 9398 32416 9404 32428
rect 9359 32388 9404 32416
rect 9398 32376 9404 32388
rect 9456 32376 9462 32428
rect 9490 32376 9496 32428
rect 9548 32376 9554 32428
rect 9968 32416 9996 32515
rect 10502 32512 10508 32524
rect 10560 32512 10566 32564
rect 13538 32552 13544 32564
rect 13499 32524 13544 32552
rect 13538 32512 13544 32524
rect 13596 32512 13602 32564
rect 10778 32444 10784 32496
rect 10836 32484 10842 32496
rect 10836 32456 11100 32484
rect 10836 32444 10842 32456
rect 11072 32425 11100 32456
rect 10965 32419 11023 32425
rect 10965 32416 10977 32419
rect 9968 32388 10977 32416
rect 10965 32385 10977 32388
rect 11011 32385 11023 32419
rect 10965 32379 11023 32385
rect 11057 32419 11115 32425
rect 11057 32385 11069 32419
rect 11103 32385 11115 32419
rect 13078 32416 13084 32428
rect 13039 32388 13084 32416
rect 11057 32379 11115 32385
rect 13078 32376 13084 32388
rect 13136 32376 13142 32428
rect 9217 32351 9275 32357
rect 9217 32348 9229 32351
rect 8680 32320 9229 32348
rect 7285 32311 7343 32317
rect 9217 32317 9229 32320
rect 9263 32348 9275 32351
rect 9306 32348 9312 32360
rect 9263 32320 9312 32348
rect 9263 32317 9275 32320
rect 9217 32311 9275 32317
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 3881 32283 3939 32289
rect 3881 32249 3893 32283
rect 3927 32280 3939 32283
rect 4240 32283 4298 32289
rect 4240 32280 4252 32283
rect 3927 32252 4252 32280
rect 3927 32249 3939 32252
rect 3881 32243 3939 32249
rect 4240 32249 4252 32252
rect 4286 32280 4298 32283
rect 4890 32280 4896 32292
rect 4286 32252 4896 32280
rect 4286 32249 4298 32252
rect 4240 32243 4298 32249
rect 4890 32240 4896 32252
rect 4948 32240 4954 32292
rect 7193 32283 7251 32289
rect 7193 32249 7205 32283
rect 7239 32280 7251 32283
rect 7374 32280 7380 32292
rect 7239 32252 7380 32280
rect 7239 32249 7251 32252
rect 7193 32243 7251 32249
rect 7374 32240 7380 32252
rect 7432 32280 7438 32292
rect 8478 32280 8484 32292
rect 7432 32252 8484 32280
rect 7432 32240 7438 32252
rect 8478 32240 8484 32252
rect 8536 32280 8542 32292
rect 8754 32280 8760 32292
rect 8536 32252 8760 32280
rect 8536 32240 8542 32252
rect 8754 32240 8760 32252
rect 8812 32240 8818 32292
rect 1673 32215 1731 32221
rect 1673 32181 1685 32215
rect 1719 32212 1731 32215
rect 1762 32212 1768 32224
rect 1719 32184 1768 32212
rect 1719 32181 1731 32184
rect 1673 32175 1731 32181
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 5350 32212 5356 32224
rect 5311 32184 5356 32212
rect 5350 32172 5356 32184
rect 5408 32172 5414 32224
rect 6822 32212 6828 32224
rect 6783 32184 6828 32212
rect 6822 32172 6828 32184
rect 6880 32172 6886 32224
rect 7834 32212 7840 32224
rect 7795 32184 7840 32212
rect 7834 32172 7840 32184
rect 7892 32212 7898 32224
rect 8205 32215 8263 32221
rect 8205 32212 8217 32215
rect 7892 32184 8217 32212
rect 7892 32172 7898 32184
rect 8205 32181 8217 32184
rect 8251 32181 8263 32215
rect 8205 32175 8263 32181
rect 8938 32172 8944 32224
rect 8996 32212 9002 32224
rect 9309 32215 9367 32221
rect 9309 32212 9321 32215
rect 8996 32184 9321 32212
rect 8996 32172 9002 32184
rect 9309 32181 9321 32184
rect 9355 32212 9367 32215
rect 9508 32212 9536 32376
rect 12805 32351 12863 32357
rect 12805 32348 12817 32351
rect 11808 32320 12817 32348
rect 9355 32184 9536 32212
rect 9355 32181 9367 32184
rect 9309 32175 9367 32181
rect 10042 32172 10048 32224
rect 10100 32212 10106 32224
rect 10321 32215 10379 32221
rect 10321 32212 10333 32215
rect 10100 32184 10333 32212
rect 10100 32172 10106 32184
rect 10321 32181 10333 32184
rect 10367 32212 10379 32215
rect 10873 32215 10931 32221
rect 10873 32212 10885 32215
rect 10367 32184 10885 32212
rect 10367 32181 10379 32184
rect 10321 32175 10379 32181
rect 10873 32181 10885 32184
rect 10919 32181 10931 32215
rect 10873 32175 10931 32181
rect 11330 32172 11336 32224
rect 11388 32212 11394 32224
rect 11808 32212 11836 32320
rect 12805 32317 12817 32320
rect 12851 32317 12863 32351
rect 12805 32311 12863 32317
rect 11885 32283 11943 32289
rect 11885 32249 11897 32283
rect 11931 32280 11943 32283
rect 12066 32280 12072 32292
rect 11931 32252 12072 32280
rect 11931 32249 11943 32252
rect 11885 32243 11943 32249
rect 12066 32240 12072 32252
rect 12124 32280 12130 32292
rect 12526 32280 12532 32292
rect 12124 32252 12532 32280
rect 12124 32240 12130 32252
rect 12526 32240 12532 32252
rect 12584 32280 12590 32292
rect 12897 32283 12955 32289
rect 12897 32280 12909 32283
rect 12584 32252 12909 32280
rect 12584 32240 12590 32252
rect 12897 32249 12909 32252
rect 12943 32249 12955 32283
rect 12897 32243 12955 32249
rect 12161 32215 12219 32221
rect 12161 32212 12173 32215
rect 11388 32184 12173 32212
rect 11388 32172 11394 32184
rect 12161 32181 12173 32184
rect 12207 32181 12219 32215
rect 12434 32212 12440 32224
rect 12395 32184 12440 32212
rect 12161 32175 12219 32181
rect 12434 32172 12440 32184
rect 12492 32172 12498 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 5902 31968 5908 32020
rect 5960 32008 5966 32020
rect 7469 32011 7527 32017
rect 7469 32008 7481 32011
rect 5960 31980 7481 32008
rect 5960 31968 5966 31980
rect 7469 31977 7481 31980
rect 7515 31977 7527 32011
rect 7469 31971 7527 31977
rect 8386 31968 8392 32020
rect 8444 32008 8450 32020
rect 9677 32011 9735 32017
rect 9677 32008 9689 32011
rect 8444 31980 9689 32008
rect 8444 31968 8450 31980
rect 9677 31977 9689 31980
rect 9723 31977 9735 32011
rect 10778 32008 10784 32020
rect 10739 31980 10784 32008
rect 9677 31971 9735 31977
rect 10778 31968 10784 31980
rect 10836 31968 10842 32020
rect 11146 32008 11152 32020
rect 11107 31980 11152 32008
rect 11146 31968 11152 31980
rect 11204 31968 11210 32020
rect 1670 31940 1676 31952
rect 1631 31912 1676 31940
rect 1670 31900 1676 31912
rect 1728 31900 1734 31952
rect 5074 31900 5080 31952
rect 5132 31940 5138 31952
rect 5252 31943 5310 31949
rect 5252 31940 5264 31943
rect 5132 31912 5264 31940
rect 5132 31900 5138 31912
rect 5252 31909 5264 31912
rect 5298 31940 5310 31943
rect 5350 31940 5356 31952
rect 5298 31912 5356 31940
rect 5298 31909 5310 31912
rect 5252 31903 5310 31909
rect 5350 31900 5356 31912
rect 5408 31900 5414 31952
rect 5442 31900 5448 31952
rect 5500 31900 5506 31952
rect 6822 31900 6828 31952
rect 6880 31940 6886 31952
rect 7837 31943 7895 31949
rect 7837 31940 7849 31943
rect 6880 31912 7849 31940
rect 6880 31900 6886 31912
rect 7837 31909 7849 31912
rect 7883 31909 7895 31943
rect 8938 31940 8944 31952
rect 8899 31912 8944 31940
rect 7837 31903 7895 31909
rect 8938 31900 8944 31912
rect 8996 31900 9002 31952
rect 9493 31943 9551 31949
rect 9493 31909 9505 31943
rect 9539 31940 9551 31943
rect 10134 31940 10140 31952
rect 9539 31912 10140 31940
rect 9539 31909 9551 31912
rect 9493 31903 9551 31909
rect 10134 31900 10140 31912
rect 10192 31900 10198 31952
rect 11164 31940 11192 31968
rect 11670 31943 11728 31949
rect 11670 31940 11682 31943
rect 11164 31912 11682 31940
rect 11670 31909 11682 31912
rect 11716 31909 11728 31943
rect 11670 31903 11728 31909
rect 1397 31875 1455 31881
rect 1397 31841 1409 31875
rect 1443 31841 1455 31875
rect 1397 31835 1455 31841
rect 1412 31804 1440 31835
rect 3970 31832 3976 31884
rect 4028 31872 4034 31884
rect 4985 31875 5043 31881
rect 4985 31872 4997 31875
rect 4028 31844 4997 31872
rect 4028 31832 4034 31844
rect 4985 31841 4997 31844
rect 5031 31872 5043 31875
rect 5460 31872 5488 31900
rect 6914 31872 6920 31884
rect 5031 31844 5488 31872
rect 6875 31844 6920 31872
rect 5031 31841 5043 31844
rect 4985 31835 5043 31841
rect 6914 31832 6920 31844
rect 6972 31832 6978 31884
rect 7006 31832 7012 31884
rect 7064 31872 7070 31884
rect 7929 31875 7987 31881
rect 7929 31872 7941 31875
rect 7064 31844 7941 31872
rect 7064 31832 7070 31844
rect 7929 31841 7941 31844
rect 7975 31841 7987 31875
rect 10042 31872 10048 31884
rect 10003 31844 10048 31872
rect 7929 31835 7987 31841
rect 10042 31832 10048 31844
rect 10100 31832 10106 31884
rect 10870 31872 10876 31884
rect 10152 31844 10876 31872
rect 10152 31816 10180 31844
rect 10870 31832 10876 31844
rect 10928 31832 10934 31884
rect 11422 31872 11428 31884
rect 11335 31844 11428 31872
rect 11422 31832 11428 31844
rect 11480 31872 11486 31884
rect 12250 31872 12256 31884
rect 11480 31844 12256 31872
rect 11480 31832 11486 31844
rect 12250 31832 12256 31844
rect 12308 31832 12314 31884
rect 1670 31804 1676 31816
rect 1412 31776 1676 31804
rect 1670 31764 1676 31776
rect 1728 31764 1734 31816
rect 7374 31804 7380 31816
rect 7335 31776 7380 31804
rect 7374 31764 7380 31776
rect 7432 31764 7438 31816
rect 8113 31807 8171 31813
rect 8113 31773 8125 31807
rect 8159 31804 8171 31807
rect 10134 31804 10140 31816
rect 8159 31776 8193 31804
rect 10047 31776 10140 31804
rect 8159 31773 8171 31776
rect 8113 31767 8171 31773
rect 6365 31739 6423 31745
rect 6365 31705 6377 31739
rect 6411 31736 6423 31739
rect 7834 31736 7840 31748
rect 6411 31708 7840 31736
rect 6411 31705 6423 31708
rect 6365 31699 6423 31705
rect 7834 31696 7840 31708
rect 7892 31696 7898 31748
rect 8128 31736 8156 31767
rect 10134 31764 10140 31776
rect 10192 31764 10198 31816
rect 10229 31807 10287 31813
rect 10229 31773 10241 31807
rect 10275 31804 10287 31807
rect 10275 31776 10309 31804
rect 10275 31773 10287 31776
rect 10229 31767 10287 31773
rect 8202 31736 8208 31748
rect 8128 31708 8208 31736
rect 8202 31696 8208 31708
rect 8260 31696 8266 31748
rect 9490 31696 9496 31748
rect 9548 31736 9554 31748
rect 10244 31736 10272 31767
rect 9548 31708 10272 31736
rect 9548 31696 9554 31708
rect 13998 31696 14004 31748
rect 14056 31736 14062 31748
rect 14918 31736 14924 31748
rect 14056 31708 14924 31736
rect 14056 31696 14062 31708
rect 14918 31696 14924 31708
rect 14976 31696 14982 31748
rect 8573 31671 8631 31677
rect 8573 31637 8585 31671
rect 8619 31668 8631 31671
rect 8662 31668 8668 31680
rect 8619 31640 8668 31668
rect 8619 31637 8631 31640
rect 8573 31631 8631 31637
rect 8662 31628 8668 31640
rect 8720 31628 8726 31680
rect 12802 31668 12808 31680
rect 12763 31640 12808 31668
rect 12802 31628 12808 31640
rect 12860 31628 12866 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 4246 31424 4252 31476
rect 4304 31464 4310 31476
rect 5074 31464 5080 31476
rect 4304 31436 5080 31464
rect 4304 31424 4310 31436
rect 5074 31424 5080 31436
rect 5132 31424 5138 31476
rect 6641 31467 6699 31473
rect 6641 31433 6653 31467
rect 6687 31464 6699 31467
rect 6822 31464 6828 31476
rect 6687 31436 6828 31464
rect 6687 31433 6699 31436
rect 6641 31427 6699 31433
rect 6822 31424 6828 31436
rect 6880 31424 6886 31476
rect 7006 31464 7012 31476
rect 6967 31436 7012 31464
rect 7006 31424 7012 31436
rect 7064 31424 7070 31476
rect 7466 31464 7472 31476
rect 7379 31436 7472 31464
rect 7466 31424 7472 31436
rect 7524 31464 7530 31476
rect 8202 31464 8208 31476
rect 7524 31436 8208 31464
rect 7524 31424 7530 31436
rect 8202 31424 8208 31436
rect 8260 31424 8266 31476
rect 8386 31424 8392 31476
rect 8444 31464 8450 31476
rect 8573 31467 8631 31473
rect 8573 31464 8585 31467
rect 8444 31436 8585 31464
rect 8444 31424 8450 31436
rect 8573 31433 8585 31436
rect 8619 31433 8631 31467
rect 10042 31464 10048 31476
rect 8573 31427 8631 31433
rect 9416 31436 10048 31464
rect 1670 31396 1676 31408
rect 1631 31368 1676 31396
rect 1670 31356 1676 31368
rect 1728 31356 1734 31408
rect 7650 31288 7656 31340
rect 7708 31328 7714 31340
rect 8110 31328 8116 31340
rect 7708 31300 8116 31328
rect 7708 31288 7714 31300
rect 8110 31288 8116 31300
rect 8168 31288 8174 31340
rect 9416 31337 9444 31436
rect 10042 31424 10048 31436
rect 10100 31464 10106 31476
rect 10229 31467 10287 31473
rect 10229 31464 10241 31467
rect 10100 31436 10241 31464
rect 10100 31424 10106 31436
rect 10229 31433 10241 31436
rect 10275 31433 10287 31467
rect 10229 31427 10287 31433
rect 11146 31424 11152 31476
rect 11204 31464 11210 31476
rect 11425 31467 11483 31473
rect 11425 31464 11437 31467
rect 11204 31436 11437 31464
rect 11204 31424 11210 31436
rect 11425 31433 11437 31436
rect 11471 31433 11483 31467
rect 11425 31427 11483 31433
rect 11977 31467 12035 31473
rect 11977 31433 11989 31467
rect 12023 31464 12035 31467
rect 12158 31464 12164 31476
rect 12023 31436 12164 31464
rect 12023 31433 12035 31436
rect 11977 31427 12035 31433
rect 12158 31424 12164 31436
rect 12216 31424 12222 31476
rect 12250 31424 12256 31476
rect 12308 31464 12314 31476
rect 12621 31467 12679 31473
rect 12621 31464 12633 31467
rect 12308 31436 12633 31464
rect 12308 31424 12314 31436
rect 12621 31433 12633 31436
rect 12667 31433 12679 31467
rect 12621 31427 12679 31433
rect 9401 31331 9459 31337
rect 9401 31297 9413 31331
rect 9447 31297 9459 31331
rect 9401 31291 9459 31297
rect 10318 31288 10324 31340
rect 10376 31328 10382 31340
rect 10870 31328 10876 31340
rect 10376 31300 10876 31328
rect 10376 31288 10382 31300
rect 10870 31288 10876 31300
rect 10928 31288 10934 31340
rect 10962 31288 10968 31340
rect 11020 31328 11026 31340
rect 11020 31300 11065 31328
rect 11020 31288 11026 31300
rect 5905 31263 5963 31269
rect 5905 31229 5917 31263
rect 5951 31260 5963 31263
rect 7926 31260 7932 31272
rect 5951 31232 7932 31260
rect 5951 31229 5963 31232
rect 5905 31223 5963 31229
rect 7926 31220 7932 31232
rect 7984 31220 7990 31272
rect 9766 31220 9772 31272
rect 9824 31260 9830 31272
rect 10042 31260 10048 31272
rect 9824 31232 10048 31260
rect 9824 31220 9830 31232
rect 10042 31220 10048 31232
rect 10100 31220 10106 31272
rect 6273 31195 6331 31201
rect 6273 31161 6285 31195
rect 6319 31192 6331 31195
rect 6638 31192 6644 31204
rect 6319 31164 6644 31192
rect 6319 31161 6331 31164
rect 6273 31155 6331 31161
rect 6638 31152 6644 31164
rect 6696 31192 6702 31204
rect 8021 31195 8079 31201
rect 8021 31192 8033 31195
rect 6696 31164 8033 31192
rect 6696 31152 6702 31164
rect 8021 31161 8033 31164
rect 8067 31161 8079 31195
rect 8021 31155 8079 31161
rect 5442 31124 5448 31136
rect 5403 31096 5448 31124
rect 5442 31084 5448 31096
rect 5500 31084 5506 31136
rect 7558 31124 7564 31136
rect 7519 31096 7564 31124
rect 7558 31084 7564 31096
rect 7616 31084 7622 31136
rect 8570 31084 8576 31136
rect 8628 31124 8634 31136
rect 9217 31127 9275 31133
rect 9217 31124 9229 31127
rect 8628 31096 9229 31124
rect 8628 31084 8634 31096
rect 9217 31093 9229 31096
rect 9263 31124 9275 31127
rect 9490 31124 9496 31136
rect 9263 31096 9496 31124
rect 9263 31093 9275 31096
rect 9217 31087 9275 31093
rect 9490 31084 9496 31096
rect 9548 31084 9554 31136
rect 9766 31084 9772 31136
rect 9824 31124 9830 31136
rect 9861 31127 9919 31133
rect 9861 31124 9873 31127
rect 9824 31096 9873 31124
rect 9824 31084 9830 31096
rect 9861 31093 9873 31096
rect 9907 31124 9919 31127
rect 10134 31124 10140 31136
rect 9907 31096 10140 31124
rect 9907 31093 9919 31096
rect 9861 31087 9919 31093
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 10410 31124 10416 31136
rect 10371 31096 10416 31124
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10778 31124 10784 31136
rect 10739 31096 10784 31124
rect 10778 31084 10784 31096
rect 10836 31084 10842 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 6365 30923 6423 30929
rect 6365 30889 6377 30923
rect 6411 30920 6423 30923
rect 6825 30923 6883 30929
rect 6825 30920 6837 30923
rect 6411 30892 6837 30920
rect 6411 30889 6423 30892
rect 6365 30883 6423 30889
rect 6825 30889 6837 30892
rect 6871 30920 6883 30923
rect 8021 30923 8079 30929
rect 8021 30920 8033 30923
rect 6871 30892 8033 30920
rect 6871 30889 6883 30892
rect 6825 30883 6883 30889
rect 8021 30889 8033 30892
rect 8067 30889 8079 30923
rect 8478 30920 8484 30932
rect 8439 30892 8484 30920
rect 8021 30883 8079 30889
rect 8478 30880 8484 30892
rect 8536 30880 8542 30932
rect 10045 30923 10103 30929
rect 10045 30889 10057 30923
rect 10091 30920 10103 30923
rect 10134 30920 10140 30932
rect 10091 30892 10140 30920
rect 10091 30889 10103 30892
rect 10045 30883 10103 30889
rect 10134 30880 10140 30892
rect 10192 30920 10198 30932
rect 10502 30920 10508 30932
rect 10192 30892 10508 30920
rect 10192 30880 10198 30892
rect 10502 30880 10508 30892
rect 10560 30880 10566 30932
rect 10870 30880 10876 30932
rect 10928 30920 10934 30932
rect 11057 30923 11115 30929
rect 11057 30920 11069 30923
rect 10928 30892 11069 30920
rect 10928 30880 10934 30892
rect 11057 30889 11069 30892
rect 11103 30889 11115 30923
rect 11057 30883 11115 30889
rect 7650 30852 7656 30864
rect 7611 30824 7656 30852
rect 7650 30812 7656 30824
rect 7708 30812 7714 30864
rect 10781 30855 10839 30861
rect 10781 30821 10793 30855
rect 10827 30852 10839 30855
rect 10962 30852 10968 30864
rect 10827 30824 10968 30852
rect 10827 30821 10839 30824
rect 10781 30815 10839 30821
rect 10962 30812 10968 30824
rect 11020 30812 11026 30864
rect 11790 30852 11796 30864
rect 11751 30824 11796 30852
rect 11790 30812 11796 30824
rect 11848 30812 11854 30864
rect 11882 30812 11888 30864
rect 11940 30852 11946 30864
rect 12434 30852 12440 30864
rect 11940 30824 12440 30852
rect 11940 30812 11946 30824
rect 12434 30812 12440 30824
rect 12492 30812 12498 30864
rect 3881 30787 3939 30793
rect 3881 30753 3893 30787
rect 3927 30784 3939 30787
rect 4522 30784 4528 30796
rect 3927 30756 4528 30784
rect 3927 30753 3939 30756
rect 3881 30747 3939 30753
rect 4522 30744 4528 30756
rect 4580 30744 4586 30796
rect 6917 30787 6975 30793
rect 6917 30753 6929 30787
rect 6963 30784 6975 30787
rect 7098 30784 7104 30796
rect 6963 30756 7104 30784
rect 6963 30753 6975 30756
rect 6917 30747 6975 30753
rect 7098 30744 7104 30756
rect 7156 30744 7162 30796
rect 8202 30744 8208 30796
rect 8260 30784 8266 30796
rect 8389 30787 8447 30793
rect 8389 30784 8401 30787
rect 8260 30756 8401 30784
rect 8260 30744 8266 30756
rect 8389 30753 8401 30756
rect 8435 30753 8447 30787
rect 8389 30747 8447 30753
rect 9858 30744 9864 30796
rect 9916 30784 9922 30796
rect 10137 30787 10195 30793
rect 10137 30784 10149 30787
rect 9916 30756 10149 30784
rect 9916 30744 9922 30756
rect 10137 30753 10149 30756
rect 10183 30753 10195 30787
rect 10137 30747 10195 30753
rect 11701 30787 11759 30793
rect 11701 30753 11713 30787
rect 11747 30784 11759 30787
rect 11974 30784 11980 30796
rect 11747 30756 11980 30784
rect 11747 30753 11759 30756
rect 11701 30747 11759 30753
rect 11974 30744 11980 30756
rect 12032 30744 12038 30796
rect 4614 30716 4620 30728
rect 4575 30688 4620 30716
rect 4614 30676 4620 30688
rect 4672 30676 4678 30728
rect 4801 30719 4859 30725
rect 4801 30685 4813 30719
rect 4847 30716 4859 30719
rect 4890 30716 4896 30728
rect 4847 30688 4896 30716
rect 4847 30685 4859 30688
rect 4801 30679 4859 30685
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 7006 30716 7012 30728
rect 6967 30688 7012 30716
rect 7006 30676 7012 30688
rect 7064 30676 7070 30728
rect 8570 30716 8576 30728
rect 8531 30688 8576 30716
rect 8570 30676 8576 30688
rect 8628 30676 8634 30728
rect 10226 30716 10232 30728
rect 10187 30688 10232 30716
rect 10226 30676 10232 30688
rect 10284 30676 10290 30728
rect 11146 30676 11152 30728
rect 11204 30716 11210 30728
rect 11885 30719 11943 30725
rect 11885 30716 11897 30719
rect 11204 30688 11897 30716
rect 11204 30676 11210 30688
rect 11885 30685 11897 30688
rect 11931 30685 11943 30719
rect 11885 30679 11943 30685
rect 6457 30651 6515 30657
rect 6457 30617 6469 30651
rect 6503 30648 6515 30651
rect 6638 30648 6644 30660
rect 6503 30620 6644 30648
rect 6503 30617 6515 30620
rect 6457 30611 6515 30617
rect 6638 30608 6644 30620
rect 6696 30608 6702 30660
rect 9674 30648 9680 30660
rect 9635 30620 9680 30648
rect 9674 30608 9680 30620
rect 9732 30608 9738 30660
rect 10778 30608 10784 30660
rect 10836 30648 10842 30660
rect 11333 30651 11391 30657
rect 11333 30648 11345 30651
rect 10836 30620 11345 30648
rect 10836 30608 10842 30620
rect 11333 30617 11345 30620
rect 11379 30617 11391 30651
rect 11333 30611 11391 30617
rect 4154 30580 4160 30592
rect 4115 30552 4160 30580
rect 4154 30540 4160 30552
rect 4212 30540 4218 30592
rect 5994 30580 6000 30592
rect 5955 30552 6000 30580
rect 5994 30540 6000 30552
rect 6052 30540 6058 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 6181 30379 6239 30385
rect 3528 30348 5488 30376
rect 2222 30308 2228 30320
rect 1412 30280 2228 30308
rect 1412 30181 1440 30280
rect 2222 30268 2228 30280
rect 2280 30268 2286 30320
rect 1578 30240 1584 30252
rect 1539 30212 1584 30240
rect 1578 30200 1584 30212
rect 1636 30200 1642 30252
rect 3528 30249 3556 30348
rect 5460 30320 5488 30348
rect 6181 30345 6193 30379
rect 6227 30376 6239 30379
rect 7006 30376 7012 30388
rect 6227 30348 7012 30376
rect 6227 30345 6239 30348
rect 6181 30339 6239 30345
rect 7006 30336 7012 30348
rect 7064 30376 7070 30388
rect 7064 30348 8616 30376
rect 7064 30336 7070 30348
rect 5442 30268 5448 30320
rect 5500 30308 5506 30320
rect 6273 30311 6331 30317
rect 6273 30308 6285 30311
rect 5500 30280 6285 30308
rect 5500 30268 5506 30280
rect 6196 30252 6224 30280
rect 6273 30277 6285 30280
rect 6319 30308 6331 30311
rect 8588 30308 8616 30348
rect 9490 30336 9496 30388
rect 9548 30376 9554 30388
rect 10045 30379 10103 30385
rect 10045 30376 10057 30379
rect 9548 30348 10057 30376
rect 9548 30336 9554 30348
rect 10045 30345 10057 30348
rect 10091 30376 10103 30379
rect 10226 30376 10232 30388
rect 10091 30348 10232 30376
rect 10091 30345 10103 30348
rect 10045 30339 10103 30345
rect 10226 30336 10232 30348
rect 10284 30336 10290 30388
rect 10778 30376 10784 30388
rect 10739 30348 10784 30376
rect 10778 30336 10784 30348
rect 10836 30336 10842 30388
rect 11146 30336 11152 30388
rect 11204 30376 11210 30388
rect 11333 30379 11391 30385
rect 11333 30376 11345 30379
rect 11204 30348 11345 30376
rect 11204 30336 11210 30348
rect 11333 30345 11345 30348
rect 11379 30345 11391 30379
rect 11790 30376 11796 30388
rect 11751 30348 11796 30376
rect 11333 30339 11391 30345
rect 11790 30336 11796 30348
rect 11848 30336 11854 30388
rect 11974 30336 11980 30388
rect 12032 30376 12038 30388
rect 12069 30379 12127 30385
rect 12069 30376 12081 30379
rect 12032 30348 12081 30376
rect 12032 30336 12038 30348
rect 12069 30345 12081 30348
rect 12115 30345 12127 30379
rect 12069 30339 12127 30345
rect 8662 30308 8668 30320
rect 6319 30280 7696 30308
rect 8575 30280 8668 30308
rect 6319 30277 6331 30280
rect 6273 30271 6331 30277
rect 3053 30243 3111 30249
rect 3053 30209 3065 30243
rect 3099 30240 3111 30243
rect 3513 30243 3571 30249
rect 3513 30240 3525 30243
rect 3099 30212 3525 30240
rect 3099 30209 3111 30212
rect 3053 30203 3111 30209
rect 3513 30209 3525 30212
rect 3559 30209 3571 30243
rect 3513 30203 3571 30209
rect 6178 30200 6184 30252
rect 6236 30200 6242 30252
rect 1397 30175 1455 30181
rect 1397 30141 1409 30175
rect 1443 30141 1455 30175
rect 1397 30135 1455 30141
rect 5994 30132 6000 30184
rect 6052 30172 6058 30184
rect 6457 30175 6515 30181
rect 6457 30172 6469 30175
rect 6052 30144 6469 30172
rect 6052 30132 6058 30144
rect 6457 30141 6469 30144
rect 6503 30172 6515 30175
rect 6638 30172 6644 30184
rect 6503 30144 6644 30172
rect 6503 30141 6515 30144
rect 6457 30135 6515 30141
rect 6638 30132 6644 30144
rect 6696 30132 6702 30184
rect 7668 30181 7696 30280
rect 8662 30268 8668 30280
rect 8720 30308 8726 30320
rect 9033 30311 9091 30317
rect 9033 30308 9045 30311
rect 8720 30280 9045 30308
rect 8720 30268 8726 30280
rect 9033 30277 9045 30280
rect 9079 30277 9091 30311
rect 9033 30271 9091 30277
rect 7653 30175 7711 30181
rect 7653 30141 7665 30175
rect 7699 30172 7711 30175
rect 8294 30172 8300 30184
rect 7699 30144 8300 30172
rect 7699 30141 7711 30144
rect 7653 30135 7711 30141
rect 8294 30132 8300 30144
rect 8352 30132 8358 30184
rect 3421 30107 3479 30113
rect 3421 30073 3433 30107
rect 3467 30104 3479 30107
rect 3780 30107 3838 30113
rect 3780 30104 3792 30107
rect 3467 30076 3792 30104
rect 3467 30073 3479 30076
rect 3421 30067 3479 30073
rect 3780 30073 3792 30076
rect 3826 30104 3838 30107
rect 4798 30104 4804 30116
rect 3826 30076 4804 30104
rect 3826 30073 3838 30076
rect 3780 30067 3838 30073
rect 4798 30064 4804 30076
rect 4856 30064 4862 30116
rect 7898 30107 7956 30113
rect 7898 30104 7910 30107
rect 7116 30076 7910 30104
rect 7116 30048 7144 30076
rect 7898 30073 7910 30076
rect 7944 30104 7956 30107
rect 8570 30104 8576 30116
rect 7944 30076 8576 30104
rect 7944 30073 7956 30076
rect 7898 30067 7956 30073
rect 8570 30064 8576 30076
rect 8628 30064 8634 30116
rect 9674 30064 9680 30116
rect 9732 30104 9738 30116
rect 9858 30104 9864 30116
rect 9732 30076 9864 30104
rect 9732 30064 9738 30076
rect 9858 30064 9864 30076
rect 9916 30104 9922 30116
rect 10413 30107 10471 30113
rect 10413 30104 10425 30107
rect 9916 30076 10425 30104
rect 9916 30064 9922 30076
rect 10413 30073 10425 30076
rect 10459 30073 10471 30107
rect 10413 30067 10471 30073
rect 4890 30036 4896 30048
rect 4851 30008 4896 30036
rect 4890 29996 4896 30008
rect 4948 30036 4954 30048
rect 5445 30039 5503 30045
rect 5445 30036 5457 30039
rect 4948 30008 5457 30036
rect 4948 29996 4954 30008
rect 5445 30005 5457 30008
rect 5491 30005 5503 30039
rect 7098 30036 7104 30048
rect 7059 30008 7104 30036
rect 5445 29999 5503 30005
rect 7098 29996 7104 30008
rect 7156 29996 7162 30048
rect 7558 30036 7564 30048
rect 7519 30008 7564 30036
rect 7558 29996 7564 30008
rect 7616 30036 7622 30048
rect 8202 30036 8208 30048
rect 7616 30008 8208 30036
rect 7616 29996 7622 30008
rect 8202 29996 8208 30008
rect 8260 29996 8266 30048
rect 9769 30039 9827 30045
rect 9769 30005 9781 30039
rect 9815 30036 9827 30039
rect 10134 30036 10140 30048
rect 9815 30008 10140 30036
rect 9815 30005 9827 30008
rect 9769 29999 9827 30005
rect 10134 29996 10140 30008
rect 10192 29996 10198 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 3881 29835 3939 29841
rect 3881 29801 3893 29835
rect 3927 29832 3939 29835
rect 4614 29832 4620 29844
rect 3927 29804 4620 29832
rect 3927 29801 3939 29804
rect 3881 29795 3939 29801
rect 4614 29792 4620 29804
rect 4672 29832 4678 29844
rect 5629 29835 5687 29841
rect 5629 29832 5641 29835
rect 4672 29804 5641 29832
rect 4672 29792 4678 29804
rect 5629 29801 5641 29804
rect 5675 29801 5687 29835
rect 7098 29832 7104 29844
rect 7059 29804 7104 29832
rect 5629 29795 5687 29801
rect 7098 29792 7104 29804
rect 7156 29792 7162 29844
rect 7282 29792 7288 29844
rect 7340 29832 7346 29844
rect 7561 29835 7619 29841
rect 7561 29832 7573 29835
rect 7340 29804 7573 29832
rect 7340 29792 7346 29804
rect 7561 29801 7573 29804
rect 7607 29832 7619 29835
rect 7650 29832 7656 29844
rect 7607 29804 7656 29832
rect 7607 29801 7619 29804
rect 7561 29795 7619 29801
rect 7650 29792 7656 29804
rect 7708 29792 7714 29844
rect 8294 29792 8300 29844
rect 8352 29832 8358 29844
rect 8573 29835 8631 29841
rect 8573 29832 8585 29835
rect 8352 29804 8585 29832
rect 8352 29792 8358 29804
rect 8573 29801 8585 29804
rect 8619 29801 8631 29835
rect 8573 29795 8631 29801
rect 10226 29792 10232 29844
rect 10284 29832 10290 29844
rect 11057 29835 11115 29841
rect 11057 29832 11069 29835
rect 10284 29804 11069 29832
rect 10284 29792 10290 29804
rect 11057 29801 11069 29804
rect 11103 29801 11115 29835
rect 11057 29795 11115 29801
rect 2774 29724 2780 29776
rect 2832 29764 2838 29776
rect 4062 29764 4068 29776
rect 2832 29736 4068 29764
rect 2832 29724 2838 29736
rect 4062 29724 4068 29736
rect 4120 29724 4126 29776
rect 6733 29767 6791 29773
rect 6733 29733 6745 29767
rect 6779 29764 6791 29767
rect 7006 29764 7012 29776
rect 6779 29736 7012 29764
rect 6779 29733 6791 29736
rect 6733 29727 6791 29733
rect 7006 29724 7012 29736
rect 7064 29724 7070 29776
rect 9858 29724 9864 29776
rect 9916 29773 9922 29776
rect 9916 29767 9980 29773
rect 9916 29733 9934 29767
rect 9968 29733 9980 29767
rect 9916 29727 9980 29733
rect 9916 29724 9922 29727
rect 2958 29656 2964 29708
rect 3016 29696 3022 29708
rect 4154 29696 4160 29708
rect 3016 29668 4160 29696
rect 3016 29656 3022 29668
rect 4154 29656 4160 29668
rect 4212 29696 4218 29708
rect 4433 29699 4491 29705
rect 4433 29696 4445 29699
rect 4212 29668 4445 29696
rect 4212 29656 4218 29668
rect 4433 29665 4445 29668
rect 4479 29665 4491 29699
rect 4433 29659 4491 29665
rect 5718 29656 5724 29708
rect 5776 29696 5782 29708
rect 5994 29696 6000 29708
rect 5776 29668 6000 29696
rect 5776 29656 5782 29668
rect 5994 29656 6000 29668
rect 6052 29656 6058 29708
rect 6089 29699 6147 29705
rect 6089 29665 6101 29699
rect 6135 29696 6147 29699
rect 6270 29696 6276 29708
rect 6135 29668 6276 29696
rect 6135 29665 6147 29668
rect 6089 29659 6147 29665
rect 6270 29656 6276 29668
rect 6328 29656 6334 29708
rect 8297 29699 8355 29705
rect 8297 29665 8309 29699
rect 8343 29696 8355 29699
rect 8478 29696 8484 29708
rect 8343 29668 8484 29696
rect 8343 29665 8355 29668
rect 8297 29659 8355 29665
rect 8478 29656 8484 29668
rect 8536 29696 8542 29708
rect 9490 29696 9496 29708
rect 8536 29668 9496 29696
rect 8536 29656 8542 29668
rect 9490 29656 9496 29668
rect 9548 29656 9554 29708
rect 9677 29699 9735 29705
rect 9677 29665 9689 29699
rect 9723 29696 9735 29699
rect 10778 29696 10784 29708
rect 9723 29668 10784 29696
rect 9723 29665 9735 29668
rect 9677 29659 9735 29665
rect 10778 29656 10784 29668
rect 10836 29656 10842 29708
rect 2866 29628 2872 29640
rect 2827 29600 2872 29628
rect 2866 29588 2872 29600
rect 2924 29588 2930 29640
rect 3050 29628 3056 29640
rect 2963 29600 3056 29628
rect 3050 29588 3056 29600
rect 3108 29628 3114 29640
rect 4246 29628 4252 29640
rect 3108 29600 4252 29628
rect 3108 29588 3114 29600
rect 4246 29588 4252 29600
rect 4304 29588 4310 29640
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29628 4583 29631
rect 4614 29628 4620 29640
rect 4571 29600 4620 29628
rect 4571 29597 4583 29600
rect 4525 29591 4583 29597
rect 4614 29588 4620 29600
rect 4672 29588 4678 29640
rect 4709 29631 4767 29637
rect 4709 29597 4721 29631
rect 4755 29628 4767 29631
rect 4798 29628 4804 29640
rect 4755 29600 4804 29628
rect 4755 29597 4767 29600
rect 4709 29591 4767 29597
rect 4798 29588 4804 29600
rect 4856 29628 4862 29640
rect 5350 29628 5356 29640
rect 4856 29600 5356 29628
rect 4856 29588 4862 29600
rect 5350 29588 5356 29600
rect 5408 29588 5414 29640
rect 6181 29631 6239 29637
rect 6181 29597 6193 29631
rect 6227 29597 6239 29631
rect 7650 29628 7656 29640
rect 7611 29600 7656 29628
rect 6181 29591 6239 29597
rect 5368 29560 5396 29588
rect 6196 29560 6224 29591
rect 7650 29588 7656 29600
rect 7708 29588 7714 29640
rect 7834 29628 7840 29640
rect 7795 29600 7840 29628
rect 7834 29588 7840 29600
rect 7892 29588 7898 29640
rect 5368 29532 6224 29560
rect 1394 29452 1400 29504
rect 1452 29492 1458 29504
rect 1673 29495 1731 29501
rect 1673 29492 1685 29495
rect 1452 29464 1685 29492
rect 1452 29452 1458 29464
rect 1673 29461 1685 29464
rect 1719 29492 1731 29495
rect 2409 29495 2467 29501
rect 2409 29492 2421 29495
rect 1719 29464 2421 29492
rect 1719 29461 1731 29464
rect 1673 29455 1731 29461
rect 2409 29461 2421 29464
rect 2455 29461 2467 29495
rect 3510 29492 3516 29504
rect 3423 29464 3516 29492
rect 2409 29455 2467 29461
rect 3510 29452 3516 29464
rect 3568 29492 3574 29504
rect 4065 29495 4123 29501
rect 4065 29492 4077 29495
rect 3568 29464 4077 29492
rect 3568 29452 3574 29464
rect 4065 29461 4077 29464
rect 4111 29461 4123 29495
rect 5166 29492 5172 29504
rect 5127 29464 5172 29492
rect 4065 29455 4123 29461
rect 5166 29452 5172 29464
rect 5224 29452 5230 29504
rect 7190 29492 7196 29504
rect 7151 29464 7196 29492
rect 7190 29452 7196 29464
rect 7248 29452 7254 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 2866 29248 2872 29300
rect 2924 29288 2930 29300
rect 3237 29291 3295 29297
rect 3237 29288 3249 29291
rect 2924 29260 3249 29288
rect 2924 29248 2930 29260
rect 3237 29257 3249 29260
rect 3283 29257 3295 29291
rect 3237 29251 3295 29257
rect 4154 29248 4160 29300
rect 4212 29288 4218 29300
rect 4341 29291 4399 29297
rect 4341 29288 4353 29291
rect 4212 29260 4353 29288
rect 4212 29248 4218 29260
rect 4341 29257 4353 29260
rect 4387 29288 4399 29291
rect 4433 29291 4491 29297
rect 4433 29288 4445 29291
rect 4387 29260 4445 29288
rect 4387 29257 4399 29260
rect 4341 29251 4399 29257
rect 4433 29257 4445 29260
rect 4479 29257 4491 29291
rect 4433 29251 4491 29257
rect 4522 29248 4528 29300
rect 4580 29288 4586 29300
rect 4801 29291 4859 29297
rect 4801 29288 4813 29291
rect 4580 29260 4813 29288
rect 4580 29248 4586 29260
rect 4801 29257 4813 29260
rect 4847 29257 4859 29291
rect 4801 29251 4859 29257
rect 7650 29248 7656 29300
rect 7708 29288 7714 29300
rect 7837 29291 7895 29297
rect 7837 29288 7849 29291
rect 7708 29260 7849 29288
rect 7708 29248 7714 29260
rect 7837 29257 7849 29260
rect 7883 29257 7895 29291
rect 7837 29251 7895 29257
rect 8662 29248 8668 29300
rect 8720 29288 8726 29300
rect 9493 29291 9551 29297
rect 9493 29288 9505 29291
rect 8720 29260 9505 29288
rect 8720 29248 8726 29260
rect 9493 29257 9505 29260
rect 9539 29288 9551 29291
rect 9539 29260 10364 29288
rect 9539 29257 9551 29260
rect 9493 29251 9551 29257
rect 2501 29223 2559 29229
rect 2501 29189 2513 29223
rect 2547 29220 2559 29223
rect 3050 29220 3056 29232
rect 2547 29192 3056 29220
rect 2547 29189 2559 29192
rect 2501 29183 2559 29189
rect 3050 29180 3056 29192
rect 3108 29180 3114 29232
rect 4246 29180 4252 29232
rect 4304 29220 4310 29232
rect 5258 29220 5264 29232
rect 4304 29192 5264 29220
rect 4304 29180 4310 29192
rect 5258 29180 5264 29192
rect 5316 29180 5322 29232
rect 6270 29220 6276 29232
rect 6231 29192 6276 29220
rect 6270 29180 6276 29192
rect 6328 29180 6334 29232
rect 9214 29180 9220 29232
rect 9272 29220 9278 29232
rect 9582 29220 9588 29232
rect 9272 29192 9588 29220
rect 9272 29180 9278 29192
rect 9582 29180 9588 29192
rect 9640 29180 9646 29232
rect 3145 29155 3203 29161
rect 3145 29121 3157 29155
rect 3191 29152 3203 29155
rect 3789 29155 3847 29161
rect 3789 29152 3801 29155
rect 3191 29124 3801 29152
rect 3191 29121 3203 29124
rect 3145 29115 3203 29121
rect 3789 29121 3801 29124
rect 3835 29152 3847 29155
rect 4890 29152 4896 29164
rect 3835 29124 4896 29152
rect 3835 29121 3847 29124
rect 3789 29115 3847 29121
rect 4890 29112 4896 29124
rect 4948 29112 4954 29164
rect 5350 29152 5356 29164
rect 5311 29124 5356 29152
rect 5350 29112 5356 29124
rect 5408 29112 5414 29164
rect 5534 29112 5540 29164
rect 5592 29152 5598 29164
rect 5592 29124 6684 29152
rect 5592 29112 5598 29124
rect 1394 29084 1400 29096
rect 1355 29056 1400 29084
rect 1394 29044 1400 29056
rect 1452 29044 1458 29096
rect 3602 29084 3608 29096
rect 3563 29056 3608 29084
rect 3602 29044 3608 29056
rect 3660 29044 3666 29096
rect 4433 29087 4491 29093
rect 4433 29053 4445 29087
rect 4479 29084 4491 29087
rect 4798 29084 4804 29096
rect 4479 29056 4804 29084
rect 4479 29053 4491 29056
rect 4433 29047 4491 29053
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 5166 29084 5172 29096
rect 5127 29056 5172 29084
rect 5166 29044 5172 29056
rect 5224 29044 5230 29096
rect 5261 29087 5319 29093
rect 5261 29053 5273 29087
rect 5307 29084 5319 29087
rect 6086 29084 6092 29096
rect 5307 29056 6092 29084
rect 5307 29053 5319 29056
rect 5261 29047 5319 29053
rect 1486 28976 1492 29028
rect 1544 29016 1550 29028
rect 1673 29019 1731 29025
rect 1673 29016 1685 29019
rect 1544 28988 1685 29016
rect 1544 28976 1550 28988
rect 1673 28985 1685 28988
rect 1719 28985 1731 29019
rect 1673 28979 1731 28985
rect 4709 29019 4767 29025
rect 4709 28985 4721 29019
rect 4755 29016 4767 29019
rect 5276 29016 5304 29047
rect 6086 29044 6092 29056
rect 6144 29044 6150 29096
rect 4755 28988 5304 29016
rect 5905 29019 5963 29025
rect 4755 28985 4767 28988
rect 4709 28979 4767 28985
rect 5905 28985 5917 29019
rect 5951 29016 5963 29019
rect 5994 29016 6000 29028
rect 5951 28988 6000 29016
rect 5951 28985 5963 28988
rect 5905 28979 5963 28985
rect 5994 28976 6000 28988
rect 6052 28976 6058 29028
rect 6656 29025 6684 29124
rect 7190 29112 7196 29164
rect 7248 29152 7254 29164
rect 7285 29155 7343 29161
rect 7285 29152 7297 29155
rect 7248 29124 7297 29152
rect 7248 29112 7254 29124
rect 7285 29121 7297 29124
rect 7331 29121 7343 29155
rect 7466 29152 7472 29164
rect 7427 29124 7472 29152
rect 7285 29115 7343 29121
rect 7300 29084 7328 29115
rect 7466 29112 7472 29124
rect 7524 29112 7530 29164
rect 9858 29112 9864 29164
rect 9916 29152 9922 29164
rect 10229 29155 10287 29161
rect 10229 29152 10241 29155
rect 9916 29124 10241 29152
rect 9916 29112 9922 29124
rect 10229 29121 10241 29124
rect 10275 29121 10287 29155
rect 10229 29115 10287 29121
rect 8205 29087 8263 29093
rect 8205 29084 8217 29087
rect 7300 29056 8217 29084
rect 8205 29053 8217 29056
rect 8251 29053 8263 29087
rect 8205 29047 8263 29053
rect 9217 29087 9275 29093
rect 9217 29053 9229 29087
rect 9263 29084 9275 29087
rect 9306 29084 9312 29096
rect 9263 29056 9312 29084
rect 9263 29053 9275 29056
rect 9217 29047 9275 29053
rect 9306 29044 9312 29056
rect 9364 29084 9370 29096
rect 9582 29084 9588 29096
rect 9364 29056 9588 29084
rect 9364 29044 9370 29056
rect 9582 29044 9588 29056
rect 9640 29084 9646 29096
rect 10045 29087 10103 29093
rect 10045 29084 10057 29087
rect 9640 29056 10057 29084
rect 9640 29044 9646 29056
rect 10045 29053 10057 29056
rect 10091 29053 10103 29087
rect 10045 29047 10103 29053
rect 10137 29087 10195 29093
rect 10137 29053 10149 29087
rect 10183 29084 10195 29087
rect 10336 29084 10364 29260
rect 10410 29084 10416 29096
rect 10183 29056 10416 29084
rect 10183 29053 10195 29056
rect 10137 29047 10195 29053
rect 10410 29044 10416 29056
rect 10468 29044 10474 29096
rect 6641 29019 6699 29025
rect 6641 28985 6653 29019
rect 6687 29016 6699 29019
rect 7193 29019 7251 29025
rect 7193 29016 7205 29019
rect 6687 28988 7205 29016
rect 6687 28985 6699 28988
rect 6641 28979 6699 28985
rect 7193 28985 7205 28988
rect 7239 29016 7251 29019
rect 7742 29016 7748 29028
rect 7239 28988 7748 29016
rect 7239 28985 7251 28988
rect 7193 28979 7251 28985
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 8849 29019 8907 29025
rect 8849 28985 8861 29019
rect 8895 29016 8907 29019
rect 9858 29016 9864 29028
rect 8895 28988 9864 29016
rect 8895 28985 8907 28988
rect 8849 28979 8907 28985
rect 9858 28976 9864 28988
rect 9916 28976 9922 29028
rect 3418 28908 3424 28960
rect 3476 28948 3482 28960
rect 3697 28951 3755 28957
rect 3697 28948 3709 28951
rect 3476 28920 3709 28948
rect 3476 28908 3482 28920
rect 3697 28917 3709 28920
rect 3743 28917 3755 28951
rect 6822 28948 6828 28960
rect 6783 28920 6828 28948
rect 3697 28911 3755 28917
rect 6822 28908 6828 28920
rect 6880 28908 6886 28960
rect 9674 28948 9680 28960
rect 9635 28920 9680 28948
rect 9674 28908 9680 28920
rect 9732 28908 9738 28960
rect 10778 28948 10784 28960
rect 10691 28920 10784 28948
rect 10778 28908 10784 28920
rect 10836 28948 10842 28960
rect 11422 28948 11428 28960
rect 10836 28920 11428 28948
rect 10836 28908 10842 28920
rect 11422 28908 11428 28920
rect 11480 28908 11486 28960
rect 12894 28908 12900 28960
rect 12952 28948 12958 28960
rect 13998 28948 14004 28960
rect 12952 28920 14004 28948
rect 12952 28908 12958 28920
rect 13998 28908 14004 28920
rect 14056 28908 14062 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 2774 28704 2780 28756
rect 2832 28744 2838 28756
rect 4341 28747 4399 28753
rect 2832 28716 2877 28744
rect 2832 28704 2838 28716
rect 4341 28713 4353 28747
rect 4387 28744 4399 28747
rect 4614 28744 4620 28756
rect 4387 28716 4620 28744
rect 4387 28713 4399 28716
rect 4341 28707 4399 28713
rect 4614 28704 4620 28716
rect 4672 28704 4678 28756
rect 4709 28747 4767 28753
rect 4709 28713 4721 28747
rect 4755 28744 4767 28747
rect 5166 28744 5172 28756
rect 4755 28716 5172 28744
rect 4755 28713 4767 28716
rect 4709 28707 4767 28713
rect 5166 28704 5172 28716
rect 5224 28704 5230 28756
rect 5902 28704 5908 28756
rect 5960 28744 5966 28756
rect 6181 28747 6239 28753
rect 6181 28744 6193 28747
rect 5960 28716 6193 28744
rect 5960 28704 5966 28716
rect 6181 28713 6193 28716
rect 6227 28713 6239 28747
rect 6181 28707 6239 28713
rect 6917 28747 6975 28753
rect 6917 28713 6929 28747
rect 6963 28744 6975 28747
rect 7190 28744 7196 28756
rect 6963 28716 7196 28744
rect 6963 28713 6975 28716
rect 6917 28707 6975 28713
rect 7190 28704 7196 28716
rect 7248 28744 7254 28756
rect 7466 28744 7472 28756
rect 7248 28716 7472 28744
rect 7248 28704 7254 28716
rect 7466 28704 7472 28716
rect 7524 28704 7530 28756
rect 7653 28747 7711 28753
rect 7653 28713 7665 28747
rect 7699 28744 7711 28747
rect 7834 28744 7840 28756
rect 7699 28716 7840 28744
rect 7699 28713 7711 28716
rect 7653 28707 7711 28713
rect 7834 28704 7840 28716
rect 7892 28704 7898 28756
rect 9858 28744 9864 28756
rect 9819 28716 9864 28744
rect 9858 28704 9864 28716
rect 9916 28704 9922 28756
rect 2501 28679 2559 28685
rect 2501 28645 2513 28679
rect 2547 28676 2559 28679
rect 2866 28676 2872 28688
rect 2547 28648 2872 28676
rect 2547 28645 2559 28648
rect 2501 28639 2559 28645
rect 2866 28636 2872 28648
rect 2924 28636 2930 28688
rect 5442 28636 5448 28688
rect 5500 28676 5506 28688
rect 6089 28679 6147 28685
rect 6089 28676 6101 28679
rect 5500 28648 6101 28676
rect 5500 28636 5506 28648
rect 6089 28645 6101 28648
rect 6135 28676 6147 28679
rect 6822 28676 6828 28688
rect 6135 28648 6828 28676
rect 6135 28645 6147 28648
rect 6089 28639 6147 28645
rect 6822 28636 6828 28648
rect 6880 28636 6886 28688
rect 7282 28676 7288 28688
rect 7243 28648 7288 28676
rect 7282 28636 7288 28648
rect 7340 28636 7346 28688
rect 11054 28636 11060 28688
rect 11112 28676 11118 28688
rect 11486 28679 11544 28685
rect 11486 28676 11498 28679
rect 11112 28648 11498 28676
rect 11112 28636 11118 28648
rect 11486 28645 11498 28648
rect 11532 28645 11544 28679
rect 11486 28639 11544 28645
rect 1397 28611 1455 28617
rect 1397 28577 1409 28611
rect 1443 28608 1455 28611
rect 1578 28608 1584 28620
rect 1443 28580 1584 28608
rect 1443 28577 1455 28580
rect 1397 28571 1455 28577
rect 1578 28568 1584 28580
rect 1636 28568 1642 28620
rect 8481 28611 8539 28617
rect 8481 28577 8493 28611
rect 8527 28608 8539 28611
rect 8846 28608 8852 28620
rect 8527 28580 8852 28608
rect 8527 28577 8539 28580
rect 8481 28571 8539 28577
rect 8846 28568 8852 28580
rect 8904 28568 8910 28620
rect 10594 28608 10600 28620
rect 10555 28580 10600 28608
rect 10594 28568 10600 28580
rect 10652 28568 10658 28620
rect 11241 28611 11299 28617
rect 11241 28577 11253 28611
rect 11287 28608 11299 28611
rect 11330 28608 11336 28620
rect 11287 28580 11336 28608
rect 11287 28577 11299 28580
rect 11241 28571 11299 28577
rect 5810 28500 5816 28552
rect 5868 28540 5874 28552
rect 6273 28543 6331 28549
rect 6273 28540 6285 28543
rect 5868 28512 6285 28540
rect 5868 28500 5874 28512
rect 6273 28509 6285 28512
rect 6319 28509 6331 28543
rect 6273 28503 6331 28509
rect 1581 28475 1639 28481
rect 1581 28441 1593 28475
rect 1627 28472 1639 28475
rect 3142 28472 3148 28484
rect 1627 28444 3148 28472
rect 1627 28441 1639 28444
rect 1581 28435 1639 28441
rect 3142 28432 3148 28444
rect 3200 28432 3206 28484
rect 3881 28475 3939 28481
rect 3881 28441 3893 28475
rect 3927 28472 3939 28475
rect 3927 28444 5212 28472
rect 3927 28441 3939 28444
rect 3881 28435 3939 28441
rect 5184 28416 5212 28444
rect 8570 28432 8576 28484
rect 8628 28472 8634 28484
rect 9217 28475 9275 28481
rect 9217 28472 9229 28475
rect 8628 28444 9229 28472
rect 8628 28432 8634 28444
rect 9217 28441 9229 28444
rect 9263 28472 9275 28475
rect 10413 28475 10471 28481
rect 10413 28472 10425 28475
rect 9263 28444 10425 28472
rect 9263 28441 9275 28444
rect 9217 28435 9275 28441
rect 10413 28441 10425 28444
rect 10459 28472 10471 28475
rect 11256 28472 11284 28571
rect 11330 28568 11336 28580
rect 11388 28568 11394 28620
rect 10459 28444 11284 28472
rect 10459 28441 10471 28444
rect 10413 28435 10471 28441
rect 3329 28407 3387 28413
rect 3329 28373 3341 28407
rect 3375 28404 3387 28407
rect 3418 28404 3424 28416
rect 3375 28376 3424 28404
rect 3375 28373 3387 28376
rect 3329 28367 3387 28373
rect 3418 28364 3424 28376
rect 3476 28364 3482 28416
rect 5166 28404 5172 28416
rect 5127 28376 5172 28404
rect 5166 28364 5172 28376
rect 5224 28404 5230 28416
rect 5350 28404 5356 28416
rect 5224 28376 5356 28404
rect 5224 28364 5230 28376
rect 5350 28364 5356 28376
rect 5408 28404 5414 28416
rect 5537 28407 5595 28413
rect 5537 28404 5549 28407
rect 5408 28376 5549 28404
rect 5408 28364 5414 28376
rect 5537 28373 5549 28376
rect 5583 28373 5595 28407
rect 5537 28367 5595 28373
rect 5626 28364 5632 28416
rect 5684 28404 5690 28416
rect 5721 28407 5779 28413
rect 5721 28404 5733 28407
rect 5684 28376 5733 28404
rect 5684 28364 5690 28376
rect 5721 28373 5733 28376
rect 5767 28373 5779 28407
rect 8294 28404 8300 28416
rect 8255 28376 8300 28404
rect 5721 28367 5779 28373
rect 8294 28364 8300 28376
rect 8352 28364 8358 28416
rect 8846 28404 8852 28416
rect 8807 28376 8852 28404
rect 8846 28364 8852 28376
rect 8904 28364 8910 28416
rect 11974 28364 11980 28416
rect 12032 28404 12038 28416
rect 12621 28407 12679 28413
rect 12621 28404 12633 28407
rect 12032 28376 12633 28404
rect 12032 28364 12038 28376
rect 12621 28373 12633 28376
rect 12667 28373 12679 28407
rect 12621 28367 12679 28373
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 5442 28200 5448 28212
rect 5403 28172 5448 28200
rect 5442 28160 5448 28172
rect 5500 28160 5506 28212
rect 5810 28200 5816 28212
rect 5771 28172 5816 28200
rect 5810 28160 5816 28172
rect 5868 28160 5874 28212
rect 5902 28160 5908 28212
rect 5960 28200 5966 28212
rect 6089 28203 6147 28209
rect 6089 28200 6101 28203
rect 5960 28172 6101 28200
rect 5960 28160 5966 28172
rect 6089 28169 6101 28172
rect 6135 28169 6147 28203
rect 6089 28163 6147 28169
rect 7558 28160 7564 28212
rect 7616 28200 7622 28212
rect 7834 28200 7840 28212
rect 7616 28172 7840 28200
rect 7616 28160 7622 28172
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 9858 28160 9864 28212
rect 9916 28200 9922 28212
rect 9953 28203 10011 28209
rect 9953 28200 9965 28203
rect 9916 28172 9965 28200
rect 9916 28160 9922 28172
rect 9953 28169 9965 28172
rect 9999 28169 10011 28203
rect 9953 28163 10011 28169
rect 11054 28160 11060 28212
rect 11112 28200 11118 28212
rect 11241 28203 11299 28209
rect 11241 28200 11253 28203
rect 11112 28172 11253 28200
rect 11112 28160 11118 28172
rect 11241 28169 11253 28172
rect 11287 28169 11299 28203
rect 11241 28163 11299 28169
rect 11422 28160 11428 28212
rect 11480 28200 11486 28212
rect 11609 28203 11667 28209
rect 11609 28200 11621 28203
rect 11480 28172 11621 28200
rect 11480 28160 11486 28172
rect 11609 28169 11621 28172
rect 11655 28169 11667 28203
rect 11609 28163 11667 28169
rect 2041 28067 2099 28073
rect 2041 28033 2053 28067
rect 2087 28064 2099 28067
rect 2406 28064 2412 28076
rect 2087 28036 2412 28064
rect 2087 28033 2099 28036
rect 2041 28027 2099 28033
rect 1397 27999 1455 28005
rect 1397 27965 1409 27999
rect 1443 27996 1455 27999
rect 1578 27996 1584 28008
rect 1443 27968 1584 27996
rect 1443 27965 1455 27968
rect 1397 27959 1455 27965
rect 1578 27956 1584 27968
rect 1636 27996 1642 28008
rect 2056 27996 2084 28027
rect 2406 28024 2412 28036
rect 2464 28024 2470 28076
rect 6641 28067 6699 28073
rect 6641 28033 6653 28067
rect 6687 28064 6699 28067
rect 7561 28067 7619 28073
rect 7561 28064 7573 28067
rect 6687 28036 7573 28064
rect 6687 28033 6699 28036
rect 6641 28027 6699 28033
rect 7561 28033 7573 28036
rect 7607 28064 7619 28067
rect 8389 28067 8447 28073
rect 8389 28064 8401 28067
rect 7607 28036 8401 28064
rect 7607 28033 7619 28036
rect 7561 28027 7619 28033
rect 8389 28033 8401 28036
rect 8435 28064 8447 28067
rect 8478 28064 8484 28076
rect 8435 28036 8484 28064
rect 8435 28033 8447 28036
rect 8389 28027 8447 28033
rect 8478 28024 8484 28036
rect 8536 28064 8542 28076
rect 8536 28036 8708 28064
rect 8536 28024 8542 28036
rect 8570 27996 8576 28008
rect 1636 27968 2084 27996
rect 8531 27968 8576 27996
rect 1636 27956 1642 27968
rect 8570 27956 8576 27968
rect 8628 27956 8634 28008
rect 8680 27996 8708 28036
rect 8829 27999 8887 28005
rect 8829 27996 8841 27999
rect 8680 27968 8841 27996
rect 8829 27965 8841 27968
rect 8875 27965 8887 27999
rect 8829 27959 8887 27965
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 2682 27860 2688 27872
rect 1627 27832 2688 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 2682 27820 2688 27832
rect 2740 27820 2746 27872
rect 7006 27860 7012 27872
rect 6967 27832 7012 27860
rect 7006 27820 7012 27832
rect 7064 27820 7070 27872
rect 7374 27860 7380 27872
rect 7335 27832 7380 27860
rect 7374 27820 7380 27832
rect 7432 27820 7438 27872
rect 7469 27863 7527 27869
rect 7469 27829 7481 27863
rect 7515 27860 7527 27863
rect 8110 27860 8116 27872
rect 7515 27832 8116 27860
rect 7515 27829 7527 27832
rect 7469 27823 7527 27829
rect 8110 27820 8116 27832
rect 8168 27820 8174 27872
rect 10594 27860 10600 27872
rect 10507 27832 10600 27860
rect 10594 27820 10600 27832
rect 10652 27860 10658 27872
rect 10962 27860 10968 27872
rect 10652 27832 10968 27860
rect 10652 27820 10658 27832
rect 10962 27820 10968 27832
rect 11020 27820 11026 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 3418 27616 3424 27668
rect 3476 27656 3482 27668
rect 4065 27659 4123 27665
rect 4065 27656 4077 27659
rect 3476 27628 4077 27656
rect 3476 27616 3482 27628
rect 4065 27625 4077 27628
rect 4111 27625 4123 27659
rect 7374 27656 7380 27668
rect 4065 27619 4123 27625
rect 6840 27628 7380 27656
rect 1670 27588 1676 27600
rect 1631 27560 1676 27588
rect 1670 27548 1676 27560
rect 1728 27548 1734 27600
rect 6089 27591 6147 27597
rect 6089 27557 6101 27591
rect 6135 27588 6147 27591
rect 6178 27588 6184 27600
rect 6135 27560 6184 27588
rect 6135 27557 6147 27560
rect 6089 27551 6147 27557
rect 6178 27548 6184 27560
rect 6236 27548 6242 27600
rect 6457 27591 6515 27597
rect 6457 27557 6469 27591
rect 6503 27588 6515 27591
rect 6840 27588 6868 27628
rect 7374 27616 7380 27628
rect 7432 27616 7438 27668
rect 8478 27656 8484 27668
rect 8439 27628 8484 27656
rect 8478 27616 8484 27628
rect 8536 27616 8542 27668
rect 9674 27656 9680 27668
rect 9635 27628 9680 27656
rect 9674 27616 9680 27628
rect 9732 27616 9738 27668
rect 11422 27616 11428 27668
rect 11480 27656 11486 27668
rect 11609 27659 11667 27665
rect 11609 27656 11621 27659
rect 11480 27628 11621 27656
rect 11480 27616 11486 27628
rect 11609 27625 11621 27628
rect 11655 27625 11667 27659
rect 11609 27619 11667 27625
rect 11974 27597 11980 27600
rect 6503 27560 6868 27588
rect 10781 27591 10839 27597
rect 6503 27557 6515 27560
rect 6457 27551 6515 27557
rect 10781 27557 10793 27591
rect 10827 27588 10839 27591
rect 11968 27588 11980 27597
rect 10827 27560 11980 27588
rect 10827 27557 10839 27560
rect 10781 27551 10839 27557
rect 11968 27551 11980 27560
rect 11974 27548 11980 27551
rect 12032 27548 12038 27600
rect 1394 27520 1400 27532
rect 1355 27492 1400 27520
rect 1394 27480 1400 27492
rect 1452 27480 1458 27532
rect 3510 27480 3516 27532
rect 3568 27520 3574 27532
rect 4433 27523 4491 27529
rect 4433 27520 4445 27523
rect 3568 27492 4445 27520
rect 3568 27480 3574 27492
rect 4433 27489 4445 27492
rect 4479 27520 4491 27523
rect 5534 27520 5540 27532
rect 4479 27492 5540 27520
rect 4479 27489 4491 27492
rect 4433 27483 4491 27489
rect 5534 27480 5540 27492
rect 5592 27480 5598 27532
rect 4522 27452 4528 27464
rect 4483 27424 4528 27452
rect 4522 27412 4528 27424
rect 4580 27412 4586 27464
rect 4709 27455 4767 27461
rect 4709 27421 4721 27455
rect 4755 27452 4767 27455
rect 5166 27452 5172 27464
rect 4755 27424 5172 27452
rect 4755 27421 4767 27424
rect 4709 27415 4767 27421
rect 5166 27412 5172 27424
rect 5224 27452 5230 27464
rect 5442 27452 5448 27464
rect 5224 27424 5448 27452
rect 5224 27412 5230 27424
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 6196 27452 6224 27548
rect 6730 27520 6736 27532
rect 6691 27492 6736 27520
rect 6730 27480 6736 27492
rect 6788 27480 6794 27532
rect 7368 27523 7426 27529
rect 7368 27489 7380 27523
rect 7414 27520 7426 27523
rect 7926 27520 7932 27532
rect 7414 27492 7932 27520
rect 7414 27489 7426 27492
rect 7368 27483 7426 27489
rect 7926 27480 7932 27492
rect 7984 27480 7990 27532
rect 10045 27523 10103 27529
rect 10045 27520 10057 27523
rect 9048 27492 10057 27520
rect 7101 27455 7159 27461
rect 7101 27452 7113 27455
rect 6196 27424 7113 27452
rect 7101 27421 7113 27424
rect 7147 27421 7159 27455
rect 7101 27415 7159 27421
rect 8478 27412 8484 27464
rect 8536 27452 8542 27464
rect 8754 27452 8760 27464
rect 8536 27424 8760 27452
rect 8536 27412 8542 27424
rect 8754 27412 8760 27424
rect 8812 27412 8818 27464
rect 6549 27387 6607 27393
rect 6549 27353 6561 27387
rect 6595 27384 6607 27387
rect 6638 27384 6644 27396
rect 6595 27356 6644 27384
rect 6595 27353 6607 27356
rect 6549 27347 6607 27353
rect 6638 27344 6644 27356
rect 6696 27344 6702 27396
rect 8754 27276 8760 27328
rect 8812 27316 8818 27328
rect 9048 27325 9076 27492
rect 10045 27489 10057 27492
rect 10091 27489 10103 27523
rect 11422 27520 11428 27532
rect 11383 27492 11428 27520
rect 10045 27483 10103 27489
rect 11422 27480 11428 27492
rect 11480 27480 11486 27532
rect 9490 27412 9496 27464
rect 9548 27452 9554 27464
rect 9674 27452 9680 27464
rect 9548 27424 9680 27452
rect 9548 27412 9554 27424
rect 9674 27412 9680 27424
rect 9732 27412 9738 27464
rect 10137 27455 10195 27461
rect 10137 27421 10149 27455
rect 10183 27421 10195 27455
rect 10137 27415 10195 27421
rect 9033 27319 9091 27325
rect 9033 27316 9045 27319
rect 8812 27288 9045 27316
rect 8812 27276 8818 27288
rect 9033 27285 9045 27288
rect 9079 27285 9091 27319
rect 9398 27316 9404 27328
rect 9359 27288 9404 27316
rect 9033 27279 9091 27285
rect 9398 27276 9404 27288
rect 9456 27316 9462 27328
rect 10152 27316 10180 27415
rect 10226 27412 10232 27464
rect 10284 27452 10290 27464
rect 11609 27455 11667 27461
rect 10284 27424 10329 27452
rect 10284 27412 10290 27424
rect 11609 27421 11621 27455
rect 11655 27452 11667 27455
rect 11701 27455 11759 27461
rect 11701 27452 11713 27455
rect 11655 27424 11713 27452
rect 11655 27421 11667 27424
rect 11609 27415 11667 27421
rect 11701 27421 11713 27424
rect 11747 27421 11759 27455
rect 11701 27415 11759 27421
rect 9456 27288 10180 27316
rect 9456 27276 9462 27288
rect 11146 27276 11152 27328
rect 11204 27316 11210 27328
rect 11241 27319 11299 27325
rect 11241 27316 11253 27319
rect 11204 27288 11253 27316
rect 11204 27276 11210 27288
rect 11241 27285 11253 27288
rect 11287 27285 11299 27319
rect 13078 27316 13084 27328
rect 13039 27288 13084 27316
rect 11241 27279 11299 27285
rect 13078 27276 13084 27288
rect 13136 27276 13142 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 1394 27072 1400 27124
rect 1452 27112 1458 27124
rect 1581 27115 1639 27121
rect 1581 27112 1593 27115
rect 1452 27084 1593 27112
rect 1452 27072 1458 27084
rect 1581 27081 1593 27084
rect 1627 27081 1639 27115
rect 3510 27112 3516 27124
rect 3471 27084 3516 27112
rect 1581 27075 1639 27081
rect 3510 27072 3516 27084
rect 3568 27072 3574 27124
rect 3973 27115 4031 27121
rect 3973 27081 3985 27115
rect 4019 27112 4031 27115
rect 4522 27112 4528 27124
rect 4019 27084 4528 27112
rect 4019 27081 4031 27084
rect 3973 27075 4031 27081
rect 4522 27072 4528 27084
rect 4580 27072 4586 27124
rect 5629 27115 5687 27121
rect 5629 27081 5641 27115
rect 5675 27112 5687 27115
rect 6730 27112 6736 27124
rect 5675 27084 6736 27112
rect 5675 27081 5687 27084
rect 5629 27075 5687 27081
rect 6730 27072 6736 27084
rect 6788 27072 6794 27124
rect 7190 27072 7196 27124
rect 7248 27072 7254 27124
rect 8570 27072 8576 27124
rect 8628 27112 8634 27124
rect 8757 27115 8815 27121
rect 8757 27112 8769 27115
rect 8628 27084 8769 27112
rect 8628 27072 8634 27084
rect 8757 27081 8769 27084
rect 8803 27112 8815 27115
rect 10410 27112 10416 27124
rect 8803 27084 9076 27112
rect 10371 27084 10416 27112
rect 8803 27081 8815 27084
rect 8757 27075 8815 27081
rect 3145 26979 3203 26985
rect 3145 26945 3157 26979
rect 3191 26976 3203 26979
rect 3970 26976 3976 26988
rect 3191 26948 3976 26976
rect 3191 26945 3203 26948
rect 3145 26939 3203 26945
rect 3970 26936 3976 26948
rect 4028 26976 4034 26988
rect 4525 26979 4583 26985
rect 4525 26976 4537 26979
rect 4028 26948 4537 26976
rect 4028 26936 4034 26948
rect 4525 26945 4537 26948
rect 4571 26945 4583 26979
rect 7208 26976 7236 27072
rect 8294 27004 8300 27056
rect 8352 27044 8358 27056
rect 8941 27047 8999 27053
rect 8941 27044 8953 27047
rect 8352 27016 8953 27044
rect 8352 27004 8358 27016
rect 8941 27013 8953 27016
rect 8987 27013 8999 27047
rect 8941 27007 8999 27013
rect 7377 26979 7435 26985
rect 7377 26976 7389 26979
rect 7208 26948 7389 26976
rect 4525 26939 4583 26945
rect 7377 26945 7389 26948
rect 7423 26976 7435 26979
rect 7466 26976 7472 26988
rect 7423 26948 7472 26976
rect 7423 26945 7435 26948
rect 7377 26939 7435 26945
rect 7466 26936 7472 26948
rect 7524 26936 7530 26988
rect 6641 26911 6699 26917
rect 6641 26877 6653 26911
rect 6687 26908 6699 26911
rect 9048 26908 9076 27084
rect 10410 27072 10416 27084
rect 10468 27072 10474 27124
rect 11422 27072 11428 27124
rect 11480 27112 11486 27124
rect 12069 27115 12127 27121
rect 12069 27112 12081 27115
rect 11480 27084 12081 27112
rect 11480 27072 11486 27084
rect 12069 27081 12081 27084
rect 12115 27081 12127 27115
rect 12069 27075 12127 27081
rect 11793 27047 11851 27053
rect 11793 27044 11805 27047
rect 11164 27016 11805 27044
rect 9490 26976 9496 26988
rect 9451 26948 9496 26976
rect 9490 26936 9496 26948
rect 9548 26936 9554 26988
rect 11054 26936 11060 26988
rect 11112 26976 11118 26988
rect 11164 26985 11192 27016
rect 11793 27013 11805 27016
rect 11839 27044 11851 27047
rect 11974 27044 11980 27056
rect 11839 27016 11980 27044
rect 11839 27013 11851 27016
rect 11793 27007 11851 27013
rect 11974 27004 11980 27016
rect 12032 27004 12038 27056
rect 11149 26979 11207 26985
rect 11149 26976 11161 26979
rect 11112 26948 11161 26976
rect 11112 26936 11118 26948
rect 11149 26945 11161 26948
rect 11195 26945 11207 26979
rect 11149 26939 11207 26945
rect 12526 26936 12532 26988
rect 12584 26976 12590 26988
rect 13354 26976 13360 26988
rect 12584 26948 13360 26976
rect 12584 26936 12590 26948
rect 13354 26936 13360 26948
rect 13412 26936 13418 26988
rect 9401 26911 9459 26917
rect 9401 26908 9413 26911
rect 6687 26880 7328 26908
rect 9048 26880 9413 26908
rect 6687 26877 6699 26880
rect 6641 26871 6699 26877
rect 7300 26852 7328 26880
rect 9401 26877 9413 26880
rect 9447 26877 9459 26911
rect 9401 26871 9459 26877
rect 10410 26868 10416 26920
rect 10468 26908 10474 26920
rect 10965 26911 11023 26917
rect 10965 26908 10977 26911
rect 10468 26880 10977 26908
rect 10468 26868 10474 26880
rect 10965 26877 10977 26880
rect 11011 26877 11023 26911
rect 10965 26871 11023 26877
rect 12802 26868 12808 26920
rect 12860 26908 12866 26920
rect 13722 26908 13728 26920
rect 12860 26880 13728 26908
rect 12860 26868 12866 26880
rect 13722 26868 13728 26880
rect 13780 26868 13786 26920
rect 3881 26843 3939 26849
rect 3881 26809 3893 26843
rect 3927 26840 3939 26843
rect 4062 26840 4068 26852
rect 3927 26812 4068 26840
rect 3927 26809 3939 26812
rect 3881 26803 3939 26809
rect 4062 26800 4068 26812
rect 4120 26840 4126 26852
rect 4433 26843 4491 26849
rect 4433 26840 4445 26843
rect 4120 26812 4445 26840
rect 4120 26800 4126 26812
rect 4433 26809 4445 26812
rect 4479 26840 4491 26843
rect 4982 26840 4988 26852
rect 4479 26812 4988 26840
rect 4479 26809 4491 26812
rect 4433 26803 4491 26809
rect 4982 26800 4988 26812
rect 5040 26800 5046 26852
rect 5721 26843 5779 26849
rect 5721 26809 5733 26843
rect 5767 26840 5779 26843
rect 6273 26843 6331 26849
rect 6273 26840 6285 26843
rect 5767 26812 6285 26840
rect 5767 26809 5779 26812
rect 5721 26803 5779 26809
rect 6273 26809 6285 26812
rect 6319 26840 6331 26843
rect 7193 26843 7251 26849
rect 7193 26840 7205 26843
rect 6319 26812 7205 26840
rect 6319 26809 6331 26812
rect 6273 26803 6331 26809
rect 7193 26809 7205 26812
rect 7239 26809 7251 26843
rect 7193 26803 7251 26809
rect 7282 26800 7288 26852
rect 7340 26840 7346 26852
rect 10873 26843 10931 26849
rect 10873 26840 10885 26843
rect 7340 26812 7385 26840
rect 9968 26812 10885 26840
rect 7340 26800 7346 26812
rect 4341 26775 4399 26781
rect 4341 26741 4353 26775
rect 4387 26772 4399 26775
rect 4614 26772 4620 26784
rect 4387 26744 4620 26772
rect 4387 26741 4399 26744
rect 4341 26735 4399 26741
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 5077 26775 5135 26781
rect 5077 26741 5089 26775
rect 5123 26772 5135 26775
rect 5442 26772 5448 26784
rect 5123 26744 5448 26772
rect 5123 26741 5135 26744
rect 5077 26735 5135 26741
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 6822 26772 6828 26784
rect 6783 26744 6828 26772
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 7926 26772 7932 26784
rect 7887 26744 7932 26772
rect 7926 26732 7932 26744
rect 7984 26732 7990 26784
rect 8386 26772 8392 26784
rect 8347 26744 8392 26772
rect 8386 26732 8392 26744
rect 8444 26772 8450 26784
rect 9309 26775 9367 26781
rect 9309 26772 9321 26775
rect 8444 26744 9321 26772
rect 8444 26732 8450 26744
rect 9309 26741 9321 26744
rect 9355 26741 9367 26775
rect 9309 26735 9367 26741
rect 9582 26732 9588 26784
rect 9640 26772 9646 26784
rect 9858 26772 9864 26784
rect 9640 26744 9864 26772
rect 9640 26732 9646 26744
rect 9858 26732 9864 26744
rect 9916 26772 9922 26784
rect 9968 26781 9996 26812
rect 10873 26809 10885 26812
rect 10919 26809 10931 26843
rect 10873 26803 10931 26809
rect 9953 26775 10011 26781
rect 9953 26772 9965 26775
rect 9916 26744 9965 26772
rect 9916 26732 9922 26744
rect 9953 26741 9965 26744
rect 9999 26741 10011 26775
rect 9953 26735 10011 26741
rect 10505 26775 10563 26781
rect 10505 26741 10517 26775
rect 10551 26772 10563 26775
rect 10778 26772 10784 26784
rect 10551 26744 10784 26772
rect 10551 26741 10563 26744
rect 10505 26735 10563 26741
rect 10778 26732 10784 26744
rect 10836 26732 10842 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 4522 26528 4528 26580
rect 4580 26568 4586 26580
rect 4617 26571 4675 26577
rect 4617 26568 4629 26571
rect 4580 26540 4629 26568
rect 4580 26528 4586 26540
rect 4617 26537 4629 26540
rect 4663 26537 4675 26571
rect 4617 26531 4675 26537
rect 5810 26528 5816 26580
rect 5868 26568 5874 26580
rect 6178 26568 6184 26580
rect 5868 26540 6184 26568
rect 5868 26528 5874 26540
rect 6178 26528 6184 26540
rect 6236 26568 6242 26580
rect 6641 26571 6699 26577
rect 6641 26568 6653 26571
rect 6236 26540 6653 26568
rect 6236 26528 6242 26540
rect 6641 26537 6653 26540
rect 6687 26537 6699 26571
rect 6641 26531 6699 26537
rect 7285 26571 7343 26577
rect 7285 26537 7297 26571
rect 7331 26568 7343 26571
rect 7466 26568 7472 26580
rect 7331 26540 7472 26568
rect 7331 26537 7343 26540
rect 7285 26531 7343 26537
rect 5528 26503 5586 26509
rect 5528 26469 5540 26503
rect 5574 26500 5586 26503
rect 7300 26500 7328 26531
rect 7466 26528 7472 26540
rect 7524 26568 7530 26580
rect 7561 26571 7619 26577
rect 7561 26568 7573 26571
rect 7524 26540 7573 26568
rect 7524 26528 7530 26540
rect 7561 26537 7573 26540
rect 7607 26537 7619 26571
rect 7561 26531 7619 26537
rect 8021 26571 8079 26577
rect 8021 26537 8033 26571
rect 8067 26568 8079 26571
rect 8754 26568 8760 26580
rect 8067 26540 8760 26568
rect 8067 26537 8079 26540
rect 8021 26531 8079 26537
rect 8754 26528 8760 26540
rect 8812 26528 8818 26580
rect 9125 26571 9183 26577
rect 9125 26537 9137 26571
rect 9171 26568 9183 26571
rect 9306 26568 9312 26580
rect 9171 26540 9312 26568
rect 9171 26537 9183 26540
rect 9125 26531 9183 26537
rect 9306 26528 9312 26540
rect 9364 26568 9370 26580
rect 9490 26568 9496 26580
rect 9364 26540 9496 26568
rect 9364 26528 9370 26540
rect 9490 26528 9496 26540
rect 9548 26528 9554 26580
rect 9953 26571 10011 26577
rect 9953 26537 9965 26571
rect 9999 26568 10011 26571
rect 10226 26568 10232 26580
rect 9999 26540 10232 26568
rect 9999 26537 10011 26540
rect 9953 26531 10011 26537
rect 10226 26528 10232 26540
rect 10284 26528 10290 26580
rect 11330 26528 11336 26580
rect 11388 26568 11394 26580
rect 11885 26571 11943 26577
rect 11885 26568 11897 26571
rect 11388 26540 11897 26568
rect 11388 26528 11394 26540
rect 11885 26537 11897 26540
rect 11931 26537 11943 26571
rect 11885 26531 11943 26537
rect 5574 26472 7328 26500
rect 5574 26469 5586 26472
rect 5528 26463 5586 26469
rect 8202 26392 8208 26444
rect 8260 26432 8266 26444
rect 8389 26435 8447 26441
rect 8389 26432 8401 26435
rect 8260 26404 8401 26432
rect 8260 26392 8266 26404
rect 8389 26401 8401 26404
rect 8435 26401 8447 26435
rect 8389 26395 8447 26401
rect 9674 26392 9680 26444
rect 9732 26432 9738 26444
rect 10873 26435 10931 26441
rect 10873 26432 10885 26435
rect 9732 26404 10885 26432
rect 9732 26392 9738 26404
rect 10873 26401 10885 26404
rect 10919 26401 10931 26435
rect 10873 26395 10931 26401
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26364 5319 26367
rect 5307 26336 5341 26364
rect 5307 26333 5319 26336
rect 5261 26327 5319 26333
rect 5169 26299 5227 26305
rect 5169 26296 5181 26299
rect 4080 26268 5181 26296
rect 4080 26240 4108 26268
rect 5169 26265 5181 26268
rect 5215 26296 5227 26299
rect 5276 26296 5304 26327
rect 8294 26324 8300 26376
rect 8352 26364 8358 26376
rect 8481 26367 8539 26373
rect 8481 26364 8493 26367
rect 8352 26336 8493 26364
rect 8352 26324 8358 26336
rect 8481 26333 8493 26336
rect 8527 26333 8539 26367
rect 8481 26327 8539 26333
rect 8665 26367 8723 26373
rect 8665 26333 8677 26367
rect 8711 26364 8723 26367
rect 9493 26367 9551 26373
rect 9493 26364 9505 26367
rect 8711 26336 9505 26364
rect 8711 26333 8723 26336
rect 8665 26327 8723 26333
rect 9493 26333 9505 26336
rect 9539 26364 9551 26367
rect 9582 26364 9588 26376
rect 9539 26336 9588 26364
rect 9539 26333 9551 26336
rect 9493 26327 9551 26333
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 9950 26324 9956 26376
rect 10008 26364 10014 26376
rect 10134 26364 10140 26376
rect 10008 26336 10140 26364
rect 10008 26324 10014 26336
rect 10134 26324 10140 26336
rect 10192 26364 10198 26376
rect 10965 26367 11023 26373
rect 10965 26364 10977 26367
rect 10192 26336 10977 26364
rect 10192 26324 10198 26336
rect 10965 26333 10977 26336
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 11054 26324 11060 26376
rect 11112 26364 11118 26376
rect 11112 26336 11157 26364
rect 11112 26324 11118 26336
rect 10229 26299 10287 26305
rect 10229 26296 10241 26299
rect 5215 26268 5304 26296
rect 5215 26265 5227 26268
rect 5169 26259 5227 26265
rect 4062 26188 4068 26240
rect 4120 26188 4126 26240
rect 4341 26231 4399 26237
rect 4341 26197 4353 26231
rect 4387 26228 4399 26231
rect 4522 26228 4528 26240
rect 4387 26200 4528 26228
rect 4387 26197 4399 26200
rect 4341 26191 4399 26197
rect 4522 26188 4528 26200
rect 4580 26188 4586 26240
rect 5276 26228 5304 26268
rect 9600 26268 10241 26296
rect 6730 26228 6736 26240
rect 5276 26200 6736 26228
rect 6730 26188 6736 26200
rect 6788 26188 6794 26240
rect 9490 26188 9496 26240
rect 9548 26228 9554 26240
rect 9600 26228 9628 26268
rect 10229 26265 10241 26268
rect 10275 26265 10287 26299
rect 11517 26299 11575 26305
rect 11517 26296 11529 26299
rect 10229 26259 10287 26265
rect 10980 26268 11529 26296
rect 10980 26240 11008 26268
rect 11517 26265 11529 26268
rect 11563 26265 11575 26299
rect 11517 26259 11575 26265
rect 9548 26200 9628 26228
rect 10505 26231 10563 26237
rect 9548 26188 9554 26200
rect 10505 26197 10517 26231
rect 10551 26228 10563 26231
rect 10962 26228 10968 26240
rect 10551 26200 10968 26228
rect 10551 26197 10563 26200
rect 10505 26191 10563 26197
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 3970 26024 3976 26036
rect 3931 25996 3976 26024
rect 3970 25984 3976 25996
rect 4028 25984 4034 26036
rect 5442 26024 5448 26036
rect 5403 25996 5448 26024
rect 5442 25984 5448 25996
rect 5500 25984 5506 26036
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 8018 26024 8024 26036
rect 7156 25996 8024 26024
rect 7156 25984 7162 25996
rect 8018 25984 8024 25996
rect 8076 26024 8082 26036
rect 8202 26024 8208 26036
rect 8076 25996 8208 26024
rect 8076 25984 8082 25996
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 8757 26027 8815 26033
rect 8757 25993 8769 26027
rect 8803 26024 8815 26027
rect 9398 26024 9404 26036
rect 8803 25996 9404 26024
rect 8803 25993 8815 25996
rect 8757 25987 8815 25993
rect 9398 25984 9404 25996
rect 9456 25984 9462 26036
rect 11054 25984 11060 26036
rect 11112 26024 11118 26036
rect 11609 26027 11667 26033
rect 11609 26024 11621 26027
rect 11112 25996 11621 26024
rect 11112 25984 11118 25996
rect 11609 25993 11621 25996
rect 11655 25993 11667 26027
rect 11609 25987 11667 25993
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 3988 25888 4016 25984
rect 10321 25959 10379 25965
rect 10321 25925 10333 25959
rect 10367 25956 10379 25959
rect 10870 25956 10876 25968
rect 10367 25928 10876 25956
rect 10367 25925 10379 25928
rect 10321 25919 10379 25925
rect 10870 25916 10876 25928
rect 10928 25916 10934 25968
rect 11977 25959 12035 25965
rect 11977 25956 11989 25959
rect 11072 25928 11989 25956
rect 7466 25888 7472 25900
rect 3988 25860 4200 25888
rect 7427 25860 7472 25888
rect 1397 25823 1455 25829
rect 1397 25789 1409 25823
rect 1443 25789 1455 25823
rect 1397 25783 1455 25789
rect 3605 25823 3663 25829
rect 3605 25789 3617 25823
rect 3651 25820 3663 25823
rect 4062 25820 4068 25832
rect 3651 25792 4068 25820
rect 3651 25789 3663 25792
rect 3605 25783 3663 25789
rect 1412 25684 1440 25783
rect 4062 25780 4068 25792
rect 4120 25780 4126 25832
rect 4172 25820 4200 25860
rect 7466 25848 7472 25860
rect 7524 25848 7530 25900
rect 9401 25891 9459 25897
rect 9401 25857 9413 25891
rect 9447 25857 9459 25891
rect 9401 25851 9459 25857
rect 4321 25823 4379 25829
rect 4321 25820 4333 25823
rect 4172 25792 4333 25820
rect 4321 25789 4333 25792
rect 4367 25820 4379 25823
rect 5442 25820 5448 25832
rect 4367 25792 5448 25820
rect 4367 25789 4379 25792
rect 4321 25783 4379 25789
rect 5442 25780 5448 25792
rect 5500 25780 5506 25832
rect 6641 25823 6699 25829
rect 6641 25789 6653 25823
rect 6687 25820 6699 25823
rect 6914 25820 6920 25832
rect 6687 25792 6920 25820
rect 6687 25789 6699 25792
rect 6641 25783 6699 25789
rect 6914 25780 6920 25792
rect 6972 25820 6978 25832
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 6972 25792 7205 25820
rect 6972 25780 6978 25792
rect 7193 25789 7205 25792
rect 7239 25820 7251 25823
rect 8202 25820 8208 25832
rect 7239 25792 8208 25820
rect 7239 25789 7251 25792
rect 7193 25783 7251 25789
rect 8202 25780 8208 25792
rect 8260 25780 8266 25832
rect 8481 25823 8539 25829
rect 8481 25789 8493 25823
rect 8527 25820 8539 25823
rect 9416 25820 9444 25851
rect 10778 25848 10784 25900
rect 10836 25888 10842 25900
rect 11072 25897 11100 25928
rect 11977 25925 11989 25928
rect 12023 25925 12035 25959
rect 11977 25919 12035 25925
rect 11057 25891 11115 25897
rect 11057 25888 11069 25891
rect 10836 25860 11069 25888
rect 10836 25848 10842 25860
rect 11057 25857 11069 25860
rect 11103 25857 11115 25891
rect 11057 25851 11115 25857
rect 11241 25891 11299 25897
rect 11241 25857 11253 25891
rect 11287 25888 11299 25891
rect 11330 25888 11336 25900
rect 11287 25860 11336 25888
rect 11287 25857 11299 25860
rect 11241 25851 11299 25857
rect 11330 25848 11336 25860
rect 11388 25848 11394 25900
rect 9490 25820 9496 25832
rect 8527 25792 9496 25820
rect 8527 25789 8539 25792
rect 8481 25783 8539 25789
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 10502 25820 10508 25832
rect 10463 25792 10508 25820
rect 10502 25780 10508 25792
rect 10560 25780 10566 25832
rect 10962 25820 10968 25832
rect 10923 25792 10968 25820
rect 10962 25780 10968 25792
rect 11020 25780 11026 25832
rect 6273 25755 6331 25761
rect 6273 25721 6285 25755
rect 6319 25752 6331 25755
rect 7282 25752 7288 25764
rect 6319 25724 7288 25752
rect 6319 25721 6331 25724
rect 6273 25715 6331 25721
rect 7282 25712 7288 25724
rect 7340 25712 7346 25764
rect 9125 25755 9183 25761
rect 9125 25721 9137 25755
rect 9171 25752 9183 25755
rect 9398 25752 9404 25764
rect 9171 25724 9404 25752
rect 9171 25721 9183 25724
rect 9125 25715 9183 25721
rect 9398 25712 9404 25724
rect 9456 25712 9462 25764
rect 2222 25684 2228 25696
rect 1412 25656 2228 25684
rect 2222 25644 2228 25656
rect 2280 25644 2286 25696
rect 6825 25687 6883 25693
rect 6825 25653 6837 25687
rect 6871 25684 6883 25687
rect 6914 25684 6920 25696
rect 6871 25656 6920 25684
rect 6871 25653 6883 25656
rect 6825 25647 6883 25653
rect 6914 25644 6920 25656
rect 6972 25644 6978 25696
rect 9217 25687 9275 25693
rect 9217 25653 9229 25687
rect 9263 25684 9275 25687
rect 9306 25684 9312 25696
rect 9263 25656 9312 25684
rect 9263 25653 9275 25656
rect 9217 25647 9275 25653
rect 9306 25644 9312 25656
rect 9364 25644 9370 25696
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 9769 25687 9827 25693
rect 9769 25684 9781 25687
rect 9732 25656 9781 25684
rect 9732 25644 9738 25656
rect 9769 25653 9781 25656
rect 9815 25653 9827 25687
rect 9769 25647 9827 25653
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 10137 25687 10195 25693
rect 10137 25684 10149 25687
rect 10008 25656 10149 25684
rect 10008 25644 10014 25656
rect 10137 25653 10149 25656
rect 10183 25653 10195 25687
rect 10594 25684 10600 25696
rect 10555 25656 10600 25684
rect 10137 25647 10195 25653
rect 10594 25644 10600 25656
rect 10652 25644 10658 25696
rect 12529 25687 12587 25693
rect 12529 25653 12541 25687
rect 12575 25684 12587 25687
rect 12710 25684 12716 25696
rect 12575 25656 12716 25684
rect 12575 25653 12587 25656
rect 12529 25647 12587 25653
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 5442 25480 5448 25492
rect 5403 25452 5448 25480
rect 5442 25440 5448 25452
rect 5500 25440 5506 25492
rect 6457 25483 6515 25489
rect 6457 25449 6469 25483
rect 6503 25480 6515 25483
rect 6638 25480 6644 25492
rect 6503 25452 6644 25480
rect 6503 25449 6515 25452
rect 6457 25443 6515 25449
rect 6638 25440 6644 25452
rect 6696 25480 6702 25492
rect 6825 25483 6883 25489
rect 6825 25480 6837 25483
rect 6696 25452 6837 25480
rect 6696 25440 6702 25452
rect 6825 25449 6837 25452
rect 6871 25449 6883 25483
rect 6825 25443 6883 25449
rect 8297 25483 8355 25489
rect 8297 25449 8309 25483
rect 8343 25480 8355 25483
rect 8662 25480 8668 25492
rect 8343 25452 8668 25480
rect 8343 25449 8355 25452
rect 8297 25443 8355 25449
rect 8662 25440 8668 25452
rect 8720 25480 8726 25492
rect 9214 25480 9220 25492
rect 8720 25452 9220 25480
rect 8720 25440 8726 25452
rect 9214 25440 9220 25452
rect 9272 25480 9278 25492
rect 9582 25480 9588 25492
rect 9272 25452 9588 25480
rect 9272 25440 9278 25452
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 10134 25440 10140 25492
rect 10192 25480 10198 25492
rect 10781 25483 10839 25489
rect 10781 25480 10793 25483
rect 10192 25452 10793 25480
rect 10192 25440 10198 25452
rect 10781 25449 10793 25452
rect 10827 25449 10839 25483
rect 10781 25443 10839 25449
rect 6089 25415 6147 25421
rect 6089 25381 6101 25415
rect 6135 25412 6147 25415
rect 7466 25412 7472 25424
rect 6135 25384 7472 25412
rect 6135 25381 6147 25384
rect 6089 25375 6147 25381
rect 7466 25372 7472 25384
rect 7524 25372 7530 25424
rect 10502 25372 10508 25424
rect 10560 25412 10566 25424
rect 11146 25412 11152 25424
rect 10560 25384 11152 25412
rect 10560 25372 10566 25384
rect 11146 25372 11152 25384
rect 11204 25412 11210 25424
rect 11793 25415 11851 25421
rect 11793 25412 11805 25415
rect 11204 25384 11805 25412
rect 11204 25372 11210 25384
rect 11793 25381 11805 25384
rect 11839 25381 11851 25415
rect 11793 25375 11851 25381
rect 4062 25344 4068 25356
rect 4023 25316 4068 25344
rect 4062 25304 4068 25316
rect 4120 25304 4126 25356
rect 4154 25304 4160 25356
rect 4212 25344 4218 25356
rect 4321 25347 4379 25353
rect 4321 25344 4333 25347
rect 4212 25316 4333 25344
rect 4212 25304 4218 25316
rect 4321 25313 4333 25316
rect 4367 25313 4379 25347
rect 4321 25307 4379 25313
rect 6733 25347 6791 25353
rect 6733 25313 6745 25347
rect 6779 25344 6791 25347
rect 6825 25347 6883 25353
rect 6825 25344 6837 25347
rect 6779 25316 6837 25344
rect 6779 25313 6791 25316
rect 6733 25307 6791 25313
rect 6825 25313 6837 25316
rect 6871 25313 6883 25347
rect 6825 25307 6883 25313
rect 7006 25304 7012 25356
rect 7064 25344 7070 25356
rect 7173 25347 7231 25353
rect 7173 25344 7185 25347
rect 7064 25316 7185 25344
rect 7064 25304 7070 25316
rect 7173 25313 7185 25316
rect 7219 25313 7231 25347
rect 7173 25307 7231 25313
rect 10321 25347 10379 25353
rect 10321 25313 10333 25347
rect 10367 25344 10379 25347
rect 12710 25344 12716 25356
rect 10367 25316 11008 25344
rect 12671 25316 12716 25344
rect 10367 25313 10379 25316
rect 10321 25307 10379 25313
rect 10980 25288 11008 25316
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 12805 25347 12863 25353
rect 12805 25313 12817 25347
rect 12851 25344 12863 25347
rect 13170 25344 13176 25356
rect 12851 25316 13176 25344
rect 12851 25313 12863 25316
rect 12805 25307 12863 25313
rect 13170 25304 13176 25316
rect 13228 25344 13234 25356
rect 13906 25344 13912 25356
rect 13228 25316 13912 25344
rect 13228 25304 13234 25316
rect 13906 25304 13912 25316
rect 13964 25304 13970 25356
rect 6917 25279 6975 25285
rect 6917 25276 6929 25279
rect 6748 25248 6929 25276
rect 6748 25152 6776 25248
rect 6917 25245 6929 25248
rect 6963 25245 6975 25279
rect 6917 25239 6975 25245
rect 8202 25236 8208 25288
rect 8260 25276 8266 25288
rect 8386 25276 8392 25288
rect 8260 25248 8392 25276
rect 8260 25236 8266 25248
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 10873 25279 10931 25285
rect 10873 25245 10885 25279
rect 10919 25245 10931 25279
rect 10873 25239 10931 25245
rect 10042 25168 10048 25220
rect 10100 25208 10106 25220
rect 10502 25208 10508 25220
rect 10100 25180 10508 25208
rect 10100 25168 10106 25180
rect 10502 25168 10508 25180
rect 10560 25208 10566 25220
rect 10888 25208 10916 25239
rect 10962 25236 10968 25288
rect 11020 25276 11026 25288
rect 12897 25279 12955 25285
rect 11020 25248 11065 25276
rect 11020 25236 11026 25248
rect 12897 25245 12909 25279
rect 12943 25245 12955 25279
rect 12897 25239 12955 25245
rect 10560 25180 10916 25208
rect 10560 25168 10566 25180
rect 11330 25168 11336 25220
rect 11388 25208 11394 25220
rect 11517 25211 11575 25217
rect 11517 25208 11529 25211
rect 11388 25180 11529 25208
rect 11388 25168 11394 25180
rect 11517 25177 11529 25180
rect 11563 25208 11575 25211
rect 12253 25211 12311 25217
rect 12253 25208 12265 25211
rect 11563 25180 12265 25208
rect 11563 25177 11575 25180
rect 11517 25171 11575 25177
rect 12253 25177 12265 25180
rect 12299 25208 12311 25211
rect 12912 25208 12940 25239
rect 13078 25208 13084 25220
rect 12299 25180 13084 25208
rect 12299 25177 12311 25180
rect 12253 25171 12311 25177
rect 13078 25168 13084 25180
rect 13136 25168 13142 25220
rect 6549 25143 6607 25149
rect 6549 25109 6561 25143
rect 6595 25140 6607 25143
rect 6730 25140 6736 25152
rect 6595 25112 6736 25140
rect 6595 25109 6607 25112
rect 6549 25103 6607 25109
rect 6730 25100 6736 25112
rect 6788 25140 6794 25152
rect 8386 25140 8392 25152
rect 6788 25112 8392 25140
rect 6788 25100 6794 25112
rect 8386 25100 8392 25112
rect 8444 25100 8450 25152
rect 9306 25100 9312 25152
rect 9364 25140 9370 25152
rect 9861 25143 9919 25149
rect 9861 25140 9873 25143
rect 9364 25112 9873 25140
rect 9364 25100 9370 25112
rect 9861 25109 9873 25112
rect 9907 25109 9919 25143
rect 10410 25140 10416 25152
rect 10371 25112 10416 25140
rect 9861 25103 9919 25109
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 12342 25140 12348 25152
rect 12303 25112 12348 25140
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 3789 24939 3847 24945
rect 3789 24905 3801 24939
rect 3835 24936 3847 24939
rect 4062 24936 4068 24948
rect 3835 24908 4068 24936
rect 3835 24905 3847 24908
rect 3789 24899 3847 24905
rect 4062 24896 4068 24908
rect 4120 24896 4126 24948
rect 5166 24936 5172 24948
rect 5127 24908 5172 24936
rect 5166 24896 5172 24908
rect 5224 24896 5230 24948
rect 6178 24936 6184 24948
rect 6139 24908 6184 24936
rect 6178 24896 6184 24908
rect 6236 24896 6242 24948
rect 6365 24939 6423 24945
rect 6365 24905 6377 24939
rect 6411 24936 6423 24939
rect 6641 24939 6699 24945
rect 6641 24936 6653 24939
rect 6411 24908 6653 24936
rect 6411 24905 6423 24908
rect 6365 24899 6423 24905
rect 6641 24905 6653 24908
rect 6687 24936 6699 24939
rect 7006 24936 7012 24948
rect 6687 24908 7012 24936
rect 6687 24905 6699 24908
rect 6641 24899 6699 24905
rect 7006 24896 7012 24908
rect 7064 24896 7070 24948
rect 9125 24939 9183 24945
rect 9125 24905 9137 24939
rect 9171 24936 9183 24939
rect 9306 24936 9312 24948
rect 9171 24908 9312 24936
rect 9171 24905 9183 24908
rect 9125 24899 9183 24905
rect 9306 24896 9312 24908
rect 9364 24896 9370 24948
rect 10042 24896 10048 24948
rect 10100 24936 10106 24948
rect 10137 24939 10195 24945
rect 10137 24936 10149 24939
rect 10100 24908 10149 24936
rect 10100 24896 10106 24908
rect 10137 24905 10149 24908
rect 10183 24905 10195 24939
rect 10137 24899 10195 24905
rect 12710 24896 12716 24948
rect 12768 24936 12774 24948
rect 13817 24939 13875 24945
rect 13817 24936 13829 24939
rect 12768 24908 13829 24936
rect 12768 24896 12774 24908
rect 13817 24905 13829 24908
rect 13863 24905 13875 24939
rect 13817 24899 13875 24905
rect 5997 24871 6055 24877
rect 5997 24837 6009 24871
rect 6043 24868 6055 24871
rect 6825 24871 6883 24877
rect 6825 24868 6837 24871
rect 6043 24840 6837 24868
rect 6043 24837 6055 24840
rect 5997 24831 6055 24837
rect 6825 24837 6837 24840
rect 6871 24837 6883 24871
rect 6825 24831 6883 24837
rect 12066 24828 12072 24880
rect 12124 24868 12130 24880
rect 12253 24871 12311 24877
rect 12253 24868 12265 24871
rect 12124 24840 12265 24868
rect 12124 24828 12130 24840
rect 12253 24837 12265 24840
rect 12299 24868 12311 24871
rect 13265 24871 13323 24877
rect 13265 24868 13277 24871
rect 12299 24840 13277 24868
rect 12299 24837 12311 24840
rect 12253 24831 12311 24837
rect 13265 24837 13277 24840
rect 13311 24837 13323 24871
rect 13265 24831 13323 24837
rect 5626 24800 5632 24812
rect 5587 24772 5632 24800
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24800 5871 24803
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 5859 24772 6377 24800
rect 5859 24769 5871 24772
rect 5813 24763 5871 24769
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 5077 24735 5135 24741
rect 5077 24701 5089 24735
rect 5123 24732 5135 24735
rect 5828 24732 5856 24763
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 6972 24772 7297 24800
rect 6972 24760 6978 24772
rect 7285 24769 7297 24772
rect 7331 24769 7343 24803
rect 7466 24800 7472 24812
rect 7427 24772 7472 24800
rect 7285 24763 7343 24769
rect 5123 24704 5856 24732
rect 7300 24732 7328 24763
rect 7466 24760 7472 24772
rect 7524 24760 7530 24812
rect 8294 24800 8300 24812
rect 8255 24772 8300 24800
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 8573 24803 8631 24809
rect 8573 24800 8585 24803
rect 8444 24772 8585 24800
rect 8444 24760 8450 24772
rect 8573 24769 8585 24772
rect 8619 24769 8631 24803
rect 8573 24763 8631 24769
rect 9582 24760 9588 24812
rect 9640 24800 9646 24812
rect 9677 24803 9735 24809
rect 9677 24800 9689 24803
rect 9640 24772 9689 24800
rect 9640 24760 9646 24772
rect 9677 24769 9689 24772
rect 9723 24769 9735 24803
rect 11330 24800 11336 24812
rect 11291 24772 11336 24800
rect 9677 24763 9735 24769
rect 11330 24760 11336 24772
rect 11388 24760 11394 24812
rect 13078 24800 13084 24812
rect 13039 24772 13084 24800
rect 13078 24760 13084 24772
rect 13136 24800 13142 24812
rect 14185 24803 14243 24809
rect 14185 24800 14197 24803
rect 13136 24772 14197 24800
rect 13136 24760 13142 24772
rect 14185 24769 14197 24772
rect 14231 24769 14243 24803
rect 14185 24763 14243 24769
rect 7837 24735 7895 24741
rect 7837 24732 7849 24735
rect 7300 24704 7849 24732
rect 5123 24701 5135 24704
rect 5077 24695 5135 24701
rect 7837 24701 7849 24704
rect 7883 24701 7895 24735
rect 8938 24732 8944 24744
rect 8899 24704 8944 24732
rect 7837 24695 7895 24701
rect 8938 24692 8944 24704
rect 8996 24692 9002 24744
rect 11057 24735 11115 24741
rect 11057 24732 11069 24735
rect 10336 24704 11069 24732
rect 4709 24667 4767 24673
rect 4709 24633 4721 24667
rect 4755 24664 4767 24667
rect 5537 24667 5595 24673
rect 5537 24664 5549 24667
rect 4755 24636 5549 24664
rect 4755 24633 4767 24636
rect 4709 24627 4767 24633
rect 5537 24633 5549 24636
rect 5583 24664 5595 24667
rect 5997 24667 6055 24673
rect 5997 24664 6009 24667
rect 5583 24636 6009 24664
rect 5583 24633 5595 24636
rect 5537 24627 5595 24633
rect 5997 24633 6009 24636
rect 6043 24633 6055 24667
rect 5997 24627 6055 24633
rect 6914 24624 6920 24676
rect 6972 24664 6978 24676
rect 7193 24667 7251 24673
rect 7193 24664 7205 24667
rect 6972 24636 7205 24664
rect 6972 24624 6978 24636
rect 7193 24633 7205 24636
rect 7239 24633 7251 24667
rect 8956 24664 8984 24692
rect 9585 24667 9643 24673
rect 9585 24664 9597 24667
rect 8956 24636 9597 24664
rect 7193 24627 7251 24633
rect 9585 24633 9597 24636
rect 9631 24633 9643 24667
rect 9585 24627 9643 24633
rect 10336 24608 10364 24704
rect 11057 24701 11069 24704
rect 11103 24701 11115 24735
rect 11057 24695 11115 24701
rect 10410 24624 10416 24676
rect 10468 24664 10474 24676
rect 11149 24667 11207 24673
rect 11149 24664 11161 24667
rect 10468 24636 11161 24664
rect 10468 24624 10474 24636
rect 11149 24633 11161 24636
rect 11195 24633 11207 24667
rect 11149 24627 11207 24633
rect 11330 24624 11336 24676
rect 11388 24664 11394 24676
rect 11885 24667 11943 24673
rect 11885 24664 11897 24667
rect 11388 24636 11897 24664
rect 11388 24624 11394 24636
rect 11885 24633 11897 24636
rect 11931 24664 11943 24667
rect 12250 24664 12256 24676
rect 11931 24636 12256 24664
rect 11931 24633 11943 24636
rect 11885 24627 11943 24633
rect 12250 24624 12256 24636
rect 12308 24664 12314 24676
rect 12897 24667 12955 24673
rect 12897 24664 12909 24667
rect 12308 24636 12909 24664
rect 12308 24624 12314 24636
rect 12897 24633 12909 24636
rect 12943 24633 12955 24667
rect 12897 24627 12955 24633
rect 13170 24624 13176 24676
rect 13228 24664 13234 24676
rect 13449 24667 13507 24673
rect 13449 24664 13461 24667
rect 13228 24636 13461 24664
rect 13228 24624 13234 24636
rect 13449 24633 13461 24636
rect 13495 24633 13507 24667
rect 13449 24627 13507 24633
rect 4154 24596 4160 24608
rect 4115 24568 4160 24596
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 9493 24599 9551 24605
rect 9493 24596 9505 24599
rect 9364 24568 9505 24596
rect 9364 24556 9370 24568
rect 9493 24565 9505 24568
rect 9539 24565 9551 24599
rect 9493 24559 9551 24565
rect 10318 24556 10324 24608
rect 10376 24596 10382 24608
rect 10505 24599 10563 24605
rect 10505 24596 10517 24599
rect 10376 24568 10517 24596
rect 10376 24556 10382 24568
rect 10505 24565 10517 24568
rect 10551 24565 10563 24599
rect 10686 24596 10692 24608
rect 10647 24568 10692 24596
rect 10505 24559 10563 24565
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 12710 24596 12716 24608
rect 12483 24568 12716 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 12805 24599 12863 24605
rect 12805 24565 12817 24599
rect 12851 24596 12863 24599
rect 13265 24599 13323 24605
rect 13265 24596 13277 24599
rect 12851 24568 13277 24596
rect 12851 24565 12863 24568
rect 12805 24559 12863 24565
rect 13265 24565 13277 24568
rect 13311 24596 13323 24599
rect 13722 24596 13728 24608
rect 13311 24568 13728 24596
rect 13311 24565 13323 24568
rect 13265 24559 13323 24565
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 5261 24395 5319 24401
rect 5261 24361 5273 24395
rect 5307 24392 5319 24395
rect 5626 24392 5632 24404
rect 5307 24364 5632 24392
rect 5307 24361 5319 24364
rect 5261 24355 5319 24361
rect 5626 24352 5632 24364
rect 5684 24352 5690 24404
rect 6914 24352 6920 24404
rect 6972 24392 6978 24404
rect 7561 24395 7619 24401
rect 7561 24392 7573 24395
rect 6972 24364 7573 24392
rect 6972 24352 6978 24364
rect 7561 24361 7573 24364
rect 7607 24361 7619 24395
rect 7561 24355 7619 24361
rect 8202 24352 8208 24404
rect 8260 24392 8266 24404
rect 9582 24392 9588 24404
rect 8260 24364 9588 24392
rect 8260 24352 8266 24364
rect 9582 24352 9588 24364
rect 9640 24352 9646 24404
rect 9953 24395 10011 24401
rect 9953 24361 9965 24395
rect 9999 24392 10011 24395
rect 10410 24392 10416 24404
rect 9999 24364 10416 24392
rect 9999 24361 10011 24364
rect 9953 24355 10011 24361
rect 10410 24352 10416 24364
rect 10468 24352 10474 24404
rect 10505 24395 10563 24401
rect 10505 24361 10517 24395
rect 10551 24392 10563 24395
rect 10594 24392 10600 24404
rect 10551 24364 10600 24392
rect 10551 24361 10563 24364
rect 10505 24355 10563 24361
rect 10594 24352 10600 24364
rect 10652 24352 10658 24404
rect 11422 24392 11428 24404
rect 11383 24364 11428 24392
rect 11422 24352 11428 24364
rect 11480 24352 11486 24404
rect 5896 24327 5954 24333
rect 5896 24293 5908 24327
rect 5942 24324 5954 24327
rect 6178 24324 6184 24336
rect 5942 24296 6184 24324
rect 5942 24293 5954 24296
rect 5896 24287 5954 24293
rect 6178 24284 6184 24296
rect 6236 24324 6242 24336
rect 7466 24324 7472 24336
rect 6236 24296 7472 24324
rect 6236 24284 6242 24296
rect 7466 24284 7472 24296
rect 7524 24284 7530 24336
rect 11440 24324 11468 24352
rect 11854 24327 11912 24333
rect 11854 24324 11866 24327
rect 11440 24296 11866 24324
rect 11854 24293 11866 24296
rect 11900 24293 11912 24327
rect 11854 24287 11912 24293
rect 4246 24216 4252 24268
rect 4304 24256 4310 24268
rect 6638 24256 6644 24268
rect 4304 24228 6644 24256
rect 4304 24216 4310 24228
rect 6638 24216 6644 24228
rect 6696 24216 6702 24268
rect 10413 24259 10471 24265
rect 10413 24225 10425 24259
rect 10459 24256 10471 24259
rect 10686 24256 10692 24268
rect 10459 24228 10692 24256
rect 10459 24225 10471 24228
rect 10413 24219 10471 24225
rect 10686 24216 10692 24228
rect 10744 24256 10750 24268
rect 11054 24256 11060 24268
rect 10744 24228 11060 24256
rect 10744 24216 10750 24228
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 5626 24188 5632 24200
rect 5587 24160 5632 24188
rect 5626 24148 5632 24160
rect 5684 24148 5690 24200
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24188 10655 24191
rect 10778 24188 10784 24200
rect 10643 24160 10784 24188
rect 10643 24157 10655 24160
rect 10597 24151 10655 24157
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 10870 24148 10876 24200
rect 10928 24188 10934 24200
rect 11146 24188 11152 24200
rect 10928 24160 11152 24188
rect 10928 24148 10934 24160
rect 11146 24148 11152 24160
rect 11204 24188 11210 24200
rect 11609 24191 11667 24197
rect 11609 24188 11621 24191
rect 11204 24160 11621 24188
rect 11204 24148 11210 24160
rect 11609 24157 11621 24160
rect 11655 24157 11667 24191
rect 11609 24151 11667 24157
rect 7006 24120 7012 24132
rect 6967 24092 7012 24120
rect 7006 24080 7012 24092
rect 7064 24080 7070 24132
rect 4522 24012 4528 24064
rect 4580 24052 4586 24064
rect 8202 24052 8208 24064
rect 4580 24024 8208 24052
rect 4580 24012 4586 24024
rect 8202 24012 8208 24024
rect 8260 24052 8266 24064
rect 9125 24055 9183 24061
rect 9125 24052 9137 24055
rect 8260 24024 9137 24052
rect 8260 24012 8266 24024
rect 9125 24021 9137 24024
rect 9171 24052 9183 24055
rect 9306 24052 9312 24064
rect 9171 24024 9312 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 10042 24052 10048 24064
rect 10003 24024 10048 24052
rect 10042 24012 10048 24024
rect 10100 24012 10106 24064
rect 10134 24012 10140 24064
rect 10192 24052 10198 24064
rect 11057 24055 11115 24061
rect 11057 24052 11069 24055
rect 10192 24024 11069 24052
rect 10192 24012 10198 24024
rect 11057 24021 11069 24024
rect 11103 24021 11115 24055
rect 12986 24052 12992 24064
rect 12947 24024 12992 24052
rect 11057 24015 11115 24021
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 5721 23851 5779 23857
rect 5721 23817 5733 23851
rect 5767 23848 5779 23851
rect 6178 23848 6184 23860
rect 5767 23820 6184 23848
rect 5767 23817 5779 23820
rect 5721 23811 5779 23817
rect 6178 23808 6184 23820
rect 6236 23808 6242 23860
rect 8662 23848 8668 23860
rect 8623 23820 8668 23848
rect 8662 23808 8668 23820
rect 8720 23808 8726 23860
rect 10778 23848 10784 23860
rect 10739 23820 10784 23848
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 11054 23848 11060 23860
rect 11015 23820 11060 23848
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 11422 23808 11428 23860
rect 11480 23848 11486 23860
rect 11609 23851 11667 23857
rect 11609 23848 11621 23851
rect 11480 23820 11621 23848
rect 11480 23808 11486 23820
rect 11609 23817 11621 23820
rect 11655 23817 11667 23851
rect 11609 23811 11667 23817
rect 8680 23712 8708 23808
rect 12986 23712 12992 23724
rect 8680 23684 8892 23712
rect 8754 23644 8760 23656
rect 8715 23616 8760 23644
rect 8754 23604 8760 23616
rect 8812 23604 8818 23656
rect 8864 23644 8892 23684
rect 12268 23684 12992 23712
rect 9013 23647 9071 23653
rect 9013 23644 9025 23647
rect 8864 23616 9025 23644
rect 9013 23613 9025 23616
rect 9059 23644 9071 23647
rect 9306 23644 9312 23656
rect 9059 23616 9312 23644
rect 9059 23613 9071 23616
rect 9013 23607 9071 23613
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 10778 23604 10784 23656
rect 10836 23644 10842 23656
rect 12158 23644 12164 23656
rect 10836 23616 12164 23644
rect 10836 23604 10842 23616
rect 12158 23604 12164 23616
rect 12216 23644 12222 23656
rect 12268 23644 12296 23684
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 12216 23616 12296 23644
rect 12216 23604 12222 23616
rect 12342 23604 12348 23656
rect 12400 23644 12406 23656
rect 12618 23644 12624 23656
rect 12400 23616 12624 23644
rect 12400 23604 12406 23616
rect 12618 23604 12624 23616
rect 12676 23604 12682 23656
rect 12710 23604 12716 23656
rect 12768 23644 12774 23656
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12768 23616 12909 23644
rect 12768 23604 12774 23616
rect 12897 23613 12909 23616
rect 12943 23644 12955 23647
rect 13449 23647 13507 23653
rect 13449 23644 13461 23647
rect 12943 23616 13461 23644
rect 12943 23613 12955 23616
rect 12897 23607 12955 23613
rect 13449 23613 13461 23616
rect 13495 23613 13507 23647
rect 13449 23607 13507 23613
rect 5626 23468 5632 23520
rect 5684 23508 5690 23520
rect 6089 23511 6147 23517
rect 6089 23508 6101 23511
rect 5684 23480 6101 23508
rect 5684 23468 5690 23480
rect 6089 23477 6101 23480
rect 6135 23508 6147 23511
rect 6730 23508 6736 23520
rect 6135 23480 6736 23508
rect 6135 23477 6147 23480
rect 6089 23471 6147 23477
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 9490 23468 9496 23520
rect 9548 23508 9554 23520
rect 10137 23511 10195 23517
rect 10137 23508 10149 23511
rect 9548 23480 10149 23508
rect 9548 23468 9554 23480
rect 10137 23477 10149 23480
rect 10183 23508 10195 23511
rect 10226 23508 10232 23520
rect 10183 23480 10232 23508
rect 10183 23477 10195 23480
rect 10137 23471 10195 23477
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 12492 23480 12537 23508
rect 12492 23468 12498 23480
rect 12618 23468 12624 23520
rect 12676 23508 12682 23520
rect 12805 23511 12863 23517
rect 12805 23508 12817 23511
rect 12676 23480 12817 23508
rect 12676 23468 12682 23480
rect 12805 23477 12817 23480
rect 12851 23508 12863 23511
rect 13817 23511 13875 23517
rect 13817 23508 13829 23511
rect 12851 23480 13829 23508
rect 12851 23477 12863 23480
rect 12805 23471 12863 23477
rect 13817 23477 13829 23480
rect 13863 23477 13875 23511
rect 13817 23471 13875 23477
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 4430 23264 4436 23316
rect 4488 23304 4494 23316
rect 4890 23304 4896 23316
rect 4488 23276 4896 23304
rect 4488 23264 4494 23276
rect 4890 23264 4896 23276
rect 4948 23304 4954 23316
rect 5169 23307 5227 23313
rect 5169 23304 5181 23307
rect 4948 23276 5181 23304
rect 4948 23264 4954 23276
rect 5169 23273 5181 23276
rect 5215 23273 5227 23307
rect 9306 23304 9312 23316
rect 9267 23276 9312 23304
rect 5169 23267 5227 23273
rect 9306 23264 9312 23276
rect 9364 23304 9370 23316
rect 9858 23304 9864 23316
rect 9364 23276 9864 23304
rect 9364 23264 9370 23276
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 10042 23264 10048 23316
rect 10100 23304 10106 23316
rect 10870 23304 10876 23316
rect 10100 23276 10876 23304
rect 10100 23264 10106 23276
rect 10870 23264 10876 23276
rect 10928 23304 10934 23316
rect 10965 23307 11023 23313
rect 10965 23304 10977 23307
rect 10928 23276 10977 23304
rect 10928 23264 10934 23276
rect 10965 23273 10977 23276
rect 11011 23273 11023 23307
rect 10965 23267 11023 23273
rect 11146 23264 11152 23316
rect 11204 23304 11210 23316
rect 11609 23307 11667 23313
rect 11609 23304 11621 23307
rect 11204 23276 11621 23304
rect 11204 23264 11210 23276
rect 11609 23273 11621 23276
rect 11655 23304 11667 23307
rect 12066 23304 12072 23316
rect 11655 23276 12072 23304
rect 11655 23273 11667 23276
rect 11609 23267 11667 23273
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 12342 23264 12348 23316
rect 12400 23264 12406 23316
rect 10137 23239 10195 23245
rect 10137 23205 10149 23239
rect 10183 23236 10195 23239
rect 10594 23236 10600 23248
rect 10183 23208 10600 23236
rect 10183 23205 10195 23208
rect 10137 23199 10195 23205
rect 10594 23196 10600 23208
rect 10652 23196 10658 23248
rect 11330 23236 11336 23248
rect 10888 23208 11336 23236
rect 9766 23128 9772 23180
rect 9824 23168 9830 23180
rect 10042 23168 10048 23180
rect 9824 23140 10048 23168
rect 9824 23128 9830 23140
rect 10042 23128 10048 23140
rect 10100 23128 10106 23180
rect 10888 23177 10916 23208
rect 11330 23196 11336 23208
rect 11388 23236 11394 23248
rect 12360 23236 12388 23264
rect 11388 23208 12388 23236
rect 11388 23196 11394 23208
rect 10873 23171 10931 23177
rect 10873 23137 10885 23171
rect 10919 23137 10931 23171
rect 12066 23168 12072 23180
rect 12027 23140 12072 23168
rect 10873 23131 10931 23137
rect 12066 23128 12072 23140
rect 12124 23128 12130 23180
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 12325 23171 12383 23177
rect 12325 23168 12337 23171
rect 12216 23140 12337 23168
rect 12216 23128 12222 23140
rect 12325 23137 12337 23140
rect 12371 23137 12383 23171
rect 12325 23131 12383 23137
rect 5261 23103 5319 23109
rect 5261 23069 5273 23103
rect 5307 23100 5319 23103
rect 5350 23100 5356 23112
rect 5307 23072 5356 23100
rect 5307 23069 5319 23072
rect 5261 23063 5319 23069
rect 5350 23060 5356 23072
rect 5408 23060 5414 23112
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 5491 23072 5856 23100
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 5828 22976 5856 23072
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 11149 23103 11207 23109
rect 11149 23100 11161 23103
rect 10652 23072 11161 23100
rect 10652 23060 10658 23072
rect 11149 23069 11161 23072
rect 11195 23100 11207 23103
rect 11195 23072 12020 23100
rect 11195 23069 11207 23072
rect 11149 23063 11207 23069
rect 10502 23032 10508 23044
rect 10463 23004 10508 23032
rect 10502 22992 10508 23004
rect 10560 22992 10566 23044
rect 2498 22924 2504 22976
rect 2556 22964 2562 22976
rect 2593 22967 2651 22973
rect 2593 22964 2605 22967
rect 2556 22936 2605 22964
rect 2556 22924 2562 22936
rect 2593 22933 2605 22936
rect 2639 22964 2651 22967
rect 2774 22964 2780 22976
rect 2639 22936 2780 22964
rect 2639 22933 2651 22936
rect 2593 22927 2651 22933
rect 2774 22924 2780 22936
rect 2832 22924 2838 22976
rect 4798 22964 4804 22976
rect 4759 22936 4804 22964
rect 4798 22924 4804 22936
rect 4856 22924 4862 22976
rect 5810 22964 5816 22976
rect 5771 22936 5816 22964
rect 5810 22924 5816 22936
rect 5868 22924 5874 22976
rect 7650 22964 7656 22976
rect 7611 22936 7656 22964
rect 7650 22924 7656 22936
rect 7708 22924 7714 22976
rect 8754 22924 8760 22976
rect 8812 22964 8818 22976
rect 8849 22967 8907 22973
rect 8849 22964 8861 22967
rect 8812 22936 8861 22964
rect 8812 22924 8818 22936
rect 8849 22933 8861 22936
rect 8895 22964 8907 22967
rect 9306 22964 9312 22976
rect 8895 22936 9312 22964
rect 8895 22933 8907 22936
rect 8849 22927 8907 22933
rect 9306 22924 9312 22936
rect 9364 22924 9370 22976
rect 11992 22964 12020 23072
rect 12342 22964 12348 22976
rect 11992 22936 12348 22964
rect 12342 22924 12348 22936
rect 12400 22964 12406 22976
rect 13449 22967 13507 22973
rect 13449 22964 13461 22967
rect 12400 22936 13461 22964
rect 12400 22924 12406 22936
rect 13449 22933 13461 22936
rect 13495 22933 13507 22967
rect 13449 22927 13507 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 4890 22760 4896 22772
rect 4851 22732 4896 22760
rect 4890 22720 4896 22732
rect 4948 22720 4954 22772
rect 5350 22720 5356 22772
rect 5408 22760 5414 22772
rect 6273 22763 6331 22769
rect 6273 22760 6285 22763
rect 5408 22732 6285 22760
rect 5408 22720 5414 22732
rect 6273 22729 6285 22732
rect 6319 22760 6331 22763
rect 7190 22760 7196 22772
rect 6319 22732 7196 22760
rect 6319 22729 6331 22732
rect 6273 22723 6331 22729
rect 7190 22720 7196 22732
rect 7248 22720 7254 22772
rect 7374 22720 7380 22772
rect 7432 22760 7438 22772
rect 7561 22763 7619 22769
rect 7561 22760 7573 22763
rect 7432 22732 7573 22760
rect 7432 22720 7438 22732
rect 7561 22729 7573 22732
rect 7607 22729 7619 22763
rect 7561 22723 7619 22729
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 9125 22763 9183 22769
rect 9125 22760 9137 22763
rect 8352 22732 9137 22760
rect 8352 22720 8358 22732
rect 9125 22729 9137 22732
rect 9171 22729 9183 22763
rect 9125 22723 9183 22729
rect 9309 22763 9367 22769
rect 9309 22729 9321 22763
rect 9355 22760 9367 22763
rect 9398 22760 9404 22772
rect 9355 22732 9404 22760
rect 9355 22729 9367 22732
rect 9309 22723 9367 22729
rect 4614 22652 4620 22704
rect 4672 22692 4678 22704
rect 5368 22692 5396 22720
rect 4672 22664 5396 22692
rect 7469 22695 7527 22701
rect 4672 22652 4678 22664
rect 7469 22661 7481 22695
rect 7515 22692 7527 22695
rect 7926 22692 7932 22704
rect 7515 22664 7932 22692
rect 7515 22661 7527 22664
rect 7469 22655 7527 22661
rect 7926 22652 7932 22664
rect 7984 22692 7990 22704
rect 7984 22664 8156 22692
rect 7984 22652 7990 22664
rect 2498 22624 2504 22636
rect 2459 22596 2504 22624
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 4246 22584 4252 22636
rect 4304 22624 4310 22636
rect 5721 22627 5779 22633
rect 5721 22624 5733 22627
rect 4304 22596 5733 22624
rect 4304 22584 4310 22596
rect 5721 22593 5733 22596
rect 5767 22624 5779 22627
rect 5810 22624 5816 22636
rect 5767 22596 5816 22624
rect 5767 22593 5779 22596
rect 5721 22587 5779 22593
rect 5810 22584 5816 22596
rect 5868 22624 5874 22636
rect 6549 22627 6607 22633
rect 6549 22624 6561 22627
rect 5868 22596 6561 22624
rect 5868 22584 5874 22596
rect 6549 22593 6561 22596
rect 6595 22624 6607 22627
rect 6914 22624 6920 22636
rect 6595 22596 6920 22624
rect 6595 22593 6607 22596
rect 6549 22587 6607 22593
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 7650 22584 7656 22636
rect 7708 22624 7714 22636
rect 8128 22633 8156 22664
rect 8021 22627 8079 22633
rect 8021 22624 8033 22627
rect 7708 22596 8033 22624
rect 7708 22584 7714 22596
rect 8021 22593 8033 22596
rect 8067 22593 8079 22627
rect 8021 22587 8079 22593
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22624 8171 22627
rect 8294 22624 8300 22636
rect 8159 22596 8300 22624
rect 8159 22593 8171 22596
rect 8113 22587 8171 22593
rect 8294 22584 8300 22596
rect 8352 22584 8358 22636
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22556 4583 22559
rect 5534 22556 5540 22568
rect 4571 22528 5540 22556
rect 4571 22525 4583 22528
rect 4525 22519 4583 22525
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 9140 22556 9168 22723
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 10594 22760 10600 22772
rect 10555 22732 10600 22760
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 10870 22760 10876 22772
rect 10831 22732 10876 22760
rect 10870 22720 10876 22732
rect 10928 22720 10934 22772
rect 11330 22760 11336 22772
rect 11291 22732 11336 22760
rect 11330 22720 11336 22732
rect 11388 22720 11394 22772
rect 11422 22720 11428 22772
rect 11480 22720 11486 22772
rect 12158 22760 12164 22772
rect 12119 22732 12164 22760
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 9858 22624 9864 22636
rect 9819 22596 9864 22624
rect 9858 22584 9864 22596
rect 9916 22584 9922 22636
rect 11440 22568 11468 22720
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9140 22528 9781 22556
rect 9769 22525 9781 22528
rect 9815 22556 9827 22559
rect 10318 22556 10324 22568
rect 9815 22528 10324 22556
rect 9815 22525 9827 22528
rect 9769 22519 9827 22525
rect 10318 22516 10324 22528
rect 10376 22516 10382 22568
rect 11422 22516 11428 22568
rect 11480 22516 11486 22568
rect 2409 22491 2467 22497
rect 2409 22457 2421 22491
rect 2455 22488 2467 22491
rect 2768 22491 2826 22497
rect 2768 22488 2780 22491
rect 2455 22460 2780 22488
rect 2455 22457 2467 22460
rect 2409 22451 2467 22457
rect 2768 22457 2780 22460
rect 2814 22488 2826 22491
rect 4062 22488 4068 22500
rect 2814 22460 4068 22488
rect 2814 22457 2826 22460
rect 2768 22451 2826 22457
rect 4062 22448 4068 22460
rect 4120 22448 4126 22500
rect 2958 22380 2964 22432
rect 3016 22420 3022 22432
rect 3881 22423 3939 22429
rect 3881 22420 3893 22423
rect 3016 22392 3893 22420
rect 3016 22380 3022 22392
rect 3881 22389 3893 22392
rect 3927 22420 3939 22423
rect 4154 22420 4160 22432
rect 3927 22392 4160 22420
rect 3927 22389 3939 22392
rect 3881 22383 3939 22389
rect 4154 22380 4160 22392
rect 4212 22380 4218 22432
rect 5166 22420 5172 22432
rect 5127 22392 5172 22420
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 5629 22423 5687 22429
rect 5629 22389 5641 22423
rect 5675 22420 5687 22423
rect 5902 22420 5908 22432
rect 5675 22392 5908 22420
rect 5675 22389 5687 22392
rect 5629 22383 5687 22389
rect 5902 22380 5908 22392
rect 5960 22380 5966 22432
rect 7101 22423 7159 22429
rect 7101 22389 7113 22423
rect 7147 22420 7159 22423
rect 7926 22420 7932 22432
rect 7147 22392 7932 22420
rect 7147 22389 7159 22392
rect 7101 22383 7159 22389
rect 7926 22380 7932 22392
rect 7984 22380 7990 22432
rect 9490 22380 9496 22432
rect 9548 22420 9554 22432
rect 9677 22423 9735 22429
rect 9677 22420 9689 22423
rect 9548 22392 9689 22420
rect 9548 22380 9554 22392
rect 9677 22389 9689 22392
rect 9723 22389 9735 22423
rect 9677 22383 9735 22389
rect 12066 22380 12072 22432
rect 12124 22420 12130 22432
rect 12618 22420 12624 22432
rect 12124 22392 12624 22420
rect 12124 22380 12130 22392
rect 12618 22380 12624 22392
rect 12676 22380 12682 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 8294 22176 8300 22228
rect 8352 22216 8358 22228
rect 8481 22219 8539 22225
rect 8481 22216 8493 22219
rect 8352 22188 8493 22216
rect 8352 22176 8358 22188
rect 8481 22185 8493 22188
rect 8527 22185 8539 22219
rect 9674 22216 9680 22228
rect 9635 22188 9680 22216
rect 8481 22179 8539 22185
rect 9674 22176 9680 22188
rect 9732 22176 9738 22228
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 10042 22216 10048 22228
rect 9824 22188 10048 22216
rect 9824 22176 9830 22188
rect 10042 22176 10048 22188
rect 10100 22176 10106 22228
rect 10137 22219 10195 22225
rect 10137 22185 10149 22219
rect 10183 22216 10195 22219
rect 12894 22216 12900 22228
rect 10183 22188 12900 22216
rect 10183 22185 10195 22188
rect 10137 22179 10195 22185
rect 4154 22108 4160 22160
rect 4212 22148 4218 22160
rect 4310 22151 4368 22157
rect 4310 22148 4322 22151
rect 4212 22120 4322 22148
rect 4212 22108 4218 22120
rect 4310 22117 4322 22120
rect 4356 22117 4368 22151
rect 4310 22111 4368 22117
rect 8202 22108 8208 22160
rect 8260 22148 8266 22160
rect 8260 22120 8340 22148
rect 8260 22108 8266 22120
rect 2317 22083 2375 22089
rect 2317 22049 2329 22083
rect 2363 22080 2375 22083
rect 2777 22083 2835 22089
rect 2777 22080 2789 22083
rect 2363 22052 2789 22080
rect 2363 22049 2375 22052
rect 2317 22043 2375 22049
rect 2777 22049 2789 22052
rect 2823 22049 2835 22083
rect 2777 22043 2835 22049
rect 2869 22083 2927 22089
rect 2869 22049 2881 22083
rect 2915 22080 2927 22083
rect 3234 22080 3240 22092
rect 2915 22052 3240 22080
rect 2915 22049 2927 22052
rect 2869 22043 2927 22049
rect 2792 21944 2820 22043
rect 3234 22040 3240 22052
rect 3292 22040 3298 22092
rect 6270 22080 6276 22092
rect 4080 22052 6276 22080
rect 2958 22012 2964 22024
rect 2919 21984 2964 22012
rect 2958 21972 2964 21984
rect 3016 21972 3022 22024
rect 4080 22021 4108 22052
rect 5644 22024 5672 22052
rect 6270 22040 6276 22052
rect 6328 22080 6334 22092
rect 6730 22080 6736 22092
rect 6328 22052 6736 22080
rect 6328 22040 6334 22052
rect 6730 22040 6736 22052
rect 6788 22080 6794 22092
rect 7374 22089 7380 22092
rect 7101 22083 7159 22089
rect 7101 22080 7113 22083
rect 6788 22052 7113 22080
rect 6788 22040 6794 22052
rect 7101 22049 7113 22052
rect 7147 22049 7159 22083
rect 7368 22080 7380 22089
rect 7335 22052 7380 22080
rect 7101 22043 7159 22049
rect 7368 22043 7380 22052
rect 7374 22040 7380 22043
rect 7432 22040 7438 22092
rect 8312 22024 8340 22120
rect 9950 22108 9956 22160
rect 10008 22148 10014 22160
rect 10152 22148 10180 22179
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 10008 22120 10180 22148
rect 10008 22108 10014 22120
rect 10042 22080 10048 22092
rect 10003 22052 10048 22080
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 12342 22089 12348 22092
rect 12336 22080 12348 22089
rect 12303 22052 12348 22080
rect 12336 22043 12348 22052
rect 12342 22040 12348 22043
rect 12400 22040 12406 22092
rect 4065 22015 4123 22021
rect 4065 22012 4077 22015
rect 3804 21984 4077 22012
rect 3326 21944 3332 21956
rect 2792 21916 3332 21944
rect 3326 21904 3332 21916
rect 3384 21904 3390 21956
rect 2130 21836 2136 21888
rect 2188 21876 2194 21888
rect 2409 21879 2467 21885
rect 2409 21876 2421 21879
rect 2188 21848 2421 21876
rect 2188 21836 2194 21848
rect 2409 21845 2421 21848
rect 2455 21845 2467 21879
rect 2409 21839 2467 21845
rect 2774 21836 2780 21888
rect 2832 21876 2838 21888
rect 3804 21885 3832 21984
rect 4065 21981 4077 21984
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 5626 21972 5632 22024
rect 5684 21972 5690 22024
rect 8294 21972 8300 22024
rect 8352 21972 8358 22024
rect 10226 21972 10232 22024
rect 10284 22012 10290 22024
rect 10284 21984 10329 22012
rect 10284 21972 10290 21984
rect 11514 21972 11520 22024
rect 11572 22012 11578 22024
rect 12069 22015 12127 22021
rect 12069 22012 12081 22015
rect 11572 21984 12081 22012
rect 11572 21972 11578 21984
rect 12069 21981 12081 21984
rect 12115 21981 12127 22015
rect 12069 21975 12127 21981
rect 3789 21879 3847 21885
rect 3789 21876 3801 21879
rect 2832 21848 3801 21876
rect 2832 21836 2838 21848
rect 3789 21845 3801 21848
rect 3835 21845 3847 21879
rect 5442 21876 5448 21888
rect 5403 21848 5448 21876
rect 3789 21839 3847 21845
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 5902 21836 5908 21888
rect 5960 21876 5966 21888
rect 6089 21879 6147 21885
rect 6089 21876 6101 21879
rect 5960 21848 6101 21876
rect 5960 21836 5966 21848
rect 6089 21845 6101 21848
rect 6135 21876 6147 21879
rect 6730 21876 6736 21888
rect 6135 21848 6736 21876
rect 6135 21845 6147 21848
rect 6089 21839 6147 21845
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 8662 21836 8668 21888
rect 8720 21876 8726 21888
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 8720 21848 9413 21876
rect 8720 21836 8726 21848
rect 9401 21845 9413 21848
rect 9447 21876 9459 21879
rect 9490 21876 9496 21888
rect 9447 21848 9496 21876
rect 9447 21845 9459 21848
rect 9401 21839 9459 21845
rect 9490 21836 9496 21848
rect 9548 21876 9554 21888
rect 10594 21876 10600 21888
rect 9548 21848 10600 21876
rect 9548 21836 9554 21848
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 13446 21876 13452 21888
rect 13407 21848 13452 21876
rect 13446 21836 13452 21848
rect 13504 21836 13510 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 5166 21632 5172 21684
rect 5224 21672 5230 21684
rect 5353 21675 5411 21681
rect 5353 21672 5365 21675
rect 5224 21644 5365 21672
rect 5224 21632 5230 21644
rect 5353 21641 5365 21644
rect 5399 21641 5411 21675
rect 6270 21672 6276 21684
rect 6231 21644 6276 21672
rect 5353 21635 5411 21641
rect 6270 21632 6276 21644
rect 6328 21632 6334 21684
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 7837 21675 7895 21681
rect 7837 21672 7849 21675
rect 7708 21644 7849 21672
rect 7708 21632 7714 21644
rect 7837 21641 7849 21644
rect 7883 21641 7895 21675
rect 7837 21635 7895 21641
rect 9769 21675 9827 21681
rect 9769 21641 9781 21675
rect 9815 21672 9827 21675
rect 9950 21672 9956 21684
rect 9815 21644 9956 21672
rect 9815 21641 9827 21644
rect 9769 21635 9827 21641
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10284 21644 10425 21672
rect 10284 21632 10290 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 10413 21635 10471 21641
rect 12161 21675 12219 21681
rect 12161 21641 12173 21675
rect 12207 21672 12219 21675
rect 12342 21672 12348 21684
rect 12207 21644 12348 21672
rect 12207 21641 12219 21644
rect 12161 21635 12219 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 12618 21672 12624 21684
rect 12579 21644 12624 21672
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 13630 21672 13636 21684
rect 13591 21644 13636 21672
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 3234 21564 3240 21616
rect 3292 21604 3298 21616
rect 3973 21607 4031 21613
rect 3973 21604 3985 21607
rect 3292 21576 3985 21604
rect 3292 21564 3298 21576
rect 3973 21573 3985 21576
rect 4019 21573 4031 21607
rect 5184 21604 5212 21632
rect 3973 21567 4031 21573
rect 4448 21576 5212 21604
rect 4448 21545 4476 21576
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21536 3111 21539
rect 4433 21539 4491 21545
rect 3099 21508 3556 21536
rect 3099 21505 3111 21508
rect 3053 21499 3111 21505
rect 2317 21471 2375 21477
rect 2317 21437 2329 21471
rect 2363 21468 2375 21471
rect 2866 21468 2872 21480
rect 2363 21440 2872 21468
rect 2363 21437 2375 21440
rect 2317 21431 2375 21437
rect 2866 21428 2872 21440
rect 2924 21428 2930 21480
rect 3528 21477 3556 21508
rect 4433 21505 4445 21539
rect 4479 21505 4491 21539
rect 4433 21499 4491 21505
rect 4522 21496 4528 21548
rect 4580 21536 4586 21548
rect 4985 21539 5043 21545
rect 4985 21536 4997 21539
rect 4580 21508 4997 21536
rect 4580 21496 4586 21508
rect 4985 21505 4997 21508
rect 5031 21536 5043 21539
rect 5442 21536 5448 21548
rect 5031 21508 5448 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21536 6699 21539
rect 7374 21536 7380 21548
rect 6687 21508 7380 21536
rect 6687 21505 6699 21508
rect 6641 21499 6699 21505
rect 7374 21496 7380 21508
rect 7432 21536 7438 21548
rect 8481 21539 8539 21545
rect 8481 21536 8493 21539
rect 7432 21508 8493 21536
rect 7432 21496 7438 21508
rect 8481 21505 8493 21508
rect 8527 21536 8539 21539
rect 10244 21536 10272 21632
rect 8527 21508 10272 21536
rect 8527 21505 8539 21508
rect 8481 21499 8539 21505
rect 3513 21471 3571 21477
rect 3513 21437 3525 21471
rect 3559 21468 3571 21471
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 3559 21440 3893 21468
rect 3559 21437 3571 21440
rect 3513 21431 3571 21437
rect 3881 21437 3893 21440
rect 3927 21468 3939 21471
rect 4246 21468 4252 21480
rect 3927 21440 4252 21468
rect 3927 21437 3939 21440
rect 3881 21431 3939 21437
rect 4246 21428 4252 21440
rect 4304 21428 4310 21480
rect 8202 21428 8208 21480
rect 8260 21468 8266 21480
rect 8297 21471 8355 21477
rect 8297 21468 8309 21471
rect 8260 21440 8309 21468
rect 8260 21428 8266 21440
rect 8297 21437 8309 21440
rect 8343 21437 8355 21471
rect 8297 21431 8355 21437
rect 12158 21428 12164 21480
rect 12216 21468 12222 21480
rect 13446 21468 13452 21480
rect 12216 21440 13452 21468
rect 12216 21428 12222 21440
rect 13446 21428 13452 21440
rect 13504 21468 13510 21480
rect 14001 21471 14059 21477
rect 14001 21468 14013 21471
rect 13504 21440 14013 21468
rect 13504 21428 13510 21440
rect 14001 21437 14013 21440
rect 14047 21437 14059 21471
rect 14001 21431 14059 21437
rect 1949 21403 2007 21409
rect 1949 21369 1961 21403
rect 1995 21400 2007 21403
rect 2777 21403 2835 21409
rect 2777 21400 2789 21403
rect 1995 21372 2789 21400
rect 1995 21369 2007 21372
rect 1949 21363 2007 21369
rect 2777 21369 2789 21372
rect 2823 21400 2835 21403
rect 5537 21403 5595 21409
rect 5537 21400 5549 21403
rect 2823 21372 5549 21400
rect 2823 21369 2835 21372
rect 2777 21363 2835 21369
rect 5537 21369 5549 21372
rect 5583 21369 5595 21403
rect 5537 21363 5595 21369
rect 2406 21332 2412 21344
rect 2367 21304 2412 21332
rect 2406 21292 2412 21304
rect 2464 21292 2470 21344
rect 2866 21332 2872 21344
rect 2827 21304 2872 21332
rect 2866 21292 2872 21304
rect 2924 21292 2930 21344
rect 4154 21292 4160 21344
rect 4212 21332 4218 21344
rect 4341 21335 4399 21341
rect 4341 21332 4353 21335
rect 4212 21304 4353 21332
rect 4212 21292 4218 21304
rect 4341 21301 4353 21304
rect 4387 21301 4399 21335
rect 4341 21295 4399 21301
rect 4982 21292 4988 21344
rect 5040 21332 5046 21344
rect 5350 21332 5356 21344
rect 5040 21304 5356 21332
rect 5040 21292 5046 21304
rect 5350 21292 5356 21304
rect 5408 21292 5414 21344
rect 7745 21335 7803 21341
rect 7745 21301 7757 21335
rect 7791 21332 7803 21335
rect 7926 21332 7932 21344
rect 7791 21304 7932 21332
rect 7791 21301 7803 21304
rect 7745 21295 7803 21301
rect 7926 21292 7932 21304
rect 7984 21332 7990 21344
rect 8110 21332 8116 21344
rect 7984 21304 8116 21332
rect 7984 21292 7990 21304
rect 8110 21292 8116 21304
rect 8168 21332 8174 21344
rect 8205 21335 8263 21341
rect 8205 21332 8217 21335
rect 8168 21304 8217 21332
rect 8168 21292 8174 21304
rect 8205 21301 8217 21304
rect 8251 21301 8263 21335
rect 10042 21332 10048 21344
rect 10003 21304 10048 21332
rect 8205 21295 8263 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 11514 21292 11520 21344
rect 11572 21332 11578 21344
rect 12618 21332 12624 21344
rect 11572 21304 12624 21332
rect 11572 21292 11578 21304
rect 12618 21292 12624 21304
rect 12676 21292 12682 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 2958 21128 2964 21140
rect 2919 21100 2964 21128
rect 2958 21088 2964 21100
rect 3016 21088 3022 21140
rect 3234 21128 3240 21140
rect 3195 21100 3240 21128
rect 3234 21088 3240 21100
rect 3292 21088 3298 21140
rect 3326 21088 3332 21140
rect 3384 21128 3390 21140
rect 4065 21131 4123 21137
rect 4065 21128 4077 21131
rect 3384 21100 4077 21128
rect 3384 21088 3390 21100
rect 4065 21097 4077 21100
rect 4111 21097 4123 21131
rect 4430 21128 4436 21140
rect 4391 21100 4436 21128
rect 4065 21091 4123 21097
rect 4430 21088 4436 21100
rect 4488 21088 4494 21140
rect 4525 21131 4583 21137
rect 4525 21097 4537 21131
rect 4571 21128 4583 21131
rect 4798 21128 4804 21140
rect 4571 21100 4804 21128
rect 4571 21097 4583 21100
rect 4525 21091 4583 21097
rect 2314 21020 2320 21072
rect 2372 21060 2378 21072
rect 2409 21063 2467 21069
rect 2409 21060 2421 21063
rect 2372 21032 2421 21060
rect 2372 21020 2378 21032
rect 2409 21029 2421 21032
rect 2455 21029 2467 21063
rect 2409 21023 2467 21029
rect 3970 21020 3976 21072
rect 4028 21060 4034 21072
rect 4540 21060 4568 21091
rect 4798 21088 4804 21100
rect 4856 21088 4862 21140
rect 6914 21088 6920 21140
rect 6972 21128 6978 21140
rect 7193 21131 7251 21137
rect 7193 21128 7205 21131
rect 6972 21100 7205 21128
rect 6972 21088 6978 21100
rect 7193 21097 7205 21100
rect 7239 21097 7251 21131
rect 7193 21091 7251 21097
rect 7929 21131 7987 21137
rect 7929 21097 7941 21131
rect 7975 21128 7987 21131
rect 8202 21128 8208 21140
rect 7975 21100 8208 21128
rect 7975 21097 7987 21100
rect 7929 21091 7987 21097
rect 8202 21088 8208 21100
rect 8260 21088 8266 21140
rect 8297 21131 8355 21137
rect 8297 21097 8309 21131
rect 8343 21128 8355 21131
rect 10042 21128 10048 21140
rect 8343 21100 10048 21128
rect 8343 21097 8355 21100
rect 8297 21091 8355 21097
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 4028 21032 4568 21060
rect 4028 21020 4034 21032
rect 5994 21020 6000 21072
rect 6052 21069 6058 21072
rect 6052 21063 6116 21069
rect 6052 21029 6070 21063
rect 6104 21029 6116 21063
rect 6052 21023 6116 21029
rect 6052 21020 6058 21023
rect 2130 20992 2136 21004
rect 2091 20964 2136 20992
rect 2130 20952 2136 20964
rect 2188 20952 2194 21004
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 5813 20995 5871 21001
rect 5813 20992 5825 20995
rect 5684 20964 5825 20992
rect 5684 20952 5690 20964
rect 5813 20961 5825 20964
rect 5859 20961 5871 20995
rect 5813 20955 5871 20961
rect 10496 20995 10554 21001
rect 10496 20961 10508 20995
rect 10542 20992 10554 20995
rect 10962 20992 10968 21004
rect 10542 20964 10968 20992
rect 10542 20961 10554 20964
rect 10496 20955 10554 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 4062 20884 4068 20936
rect 4120 20924 4126 20936
rect 4522 20924 4528 20936
rect 4120 20896 4528 20924
rect 4120 20884 4126 20896
rect 4522 20884 4528 20896
rect 4580 20924 4586 20936
rect 4617 20927 4675 20933
rect 4617 20924 4629 20927
rect 4580 20896 4629 20924
rect 4580 20884 4586 20896
rect 4617 20893 4629 20896
rect 4663 20893 4675 20927
rect 4617 20887 4675 20893
rect 9306 20884 9312 20936
rect 9364 20924 9370 20936
rect 9401 20927 9459 20933
rect 9401 20924 9413 20927
rect 9364 20896 9413 20924
rect 9364 20884 9370 20896
rect 9401 20893 9413 20896
rect 9447 20924 9459 20927
rect 10226 20924 10232 20936
rect 9447 20896 10232 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 10226 20884 10232 20896
rect 10284 20884 10290 20936
rect 3881 20859 3939 20865
rect 3881 20825 3893 20859
rect 3927 20856 3939 20859
rect 4154 20856 4160 20868
rect 3927 20828 4160 20856
rect 3927 20825 3939 20828
rect 3881 20819 3939 20825
rect 4154 20816 4160 20828
rect 4212 20816 4218 20868
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 11609 20791 11667 20797
rect 11609 20788 11621 20791
rect 11204 20760 11621 20788
rect 11204 20748 11210 20760
rect 11609 20757 11621 20760
rect 11655 20757 11667 20791
rect 11609 20751 11667 20757
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 2130 20584 2136 20596
rect 2091 20556 2136 20584
rect 2130 20544 2136 20556
rect 2188 20544 2194 20596
rect 3329 20587 3387 20593
rect 3329 20553 3341 20587
rect 3375 20584 3387 20587
rect 3970 20584 3976 20596
rect 3375 20556 3976 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 4154 20544 4160 20596
rect 4212 20584 4218 20596
rect 4525 20587 4583 20593
rect 4525 20584 4537 20587
rect 4212 20556 4537 20584
rect 4212 20544 4218 20556
rect 4525 20553 4537 20556
rect 4571 20553 4583 20587
rect 4525 20547 4583 20553
rect 5626 20544 5632 20596
rect 5684 20584 5690 20596
rect 6181 20587 6239 20593
rect 6181 20584 6193 20587
rect 5684 20556 6193 20584
rect 5684 20544 5690 20556
rect 6181 20553 6193 20556
rect 6227 20553 6239 20587
rect 6181 20547 6239 20553
rect 3697 20519 3755 20525
rect 3697 20485 3709 20519
rect 3743 20516 3755 20519
rect 4062 20516 4068 20528
rect 3743 20488 4068 20516
rect 3743 20485 3755 20488
rect 3697 20479 3755 20485
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20448 4031 20451
rect 4246 20448 4252 20460
rect 4019 20420 4252 20448
rect 4019 20417 4031 20420
rect 3973 20411 4031 20417
rect 4246 20408 4252 20420
rect 4304 20448 4310 20460
rect 5077 20451 5135 20457
rect 5077 20448 5089 20451
rect 4304 20420 5089 20448
rect 4304 20408 4310 20420
rect 5077 20417 5089 20420
rect 5123 20417 5135 20451
rect 6196 20448 6224 20547
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11241 20587 11299 20593
rect 11241 20584 11253 20587
rect 11112 20556 11253 20584
rect 11112 20544 11118 20556
rect 11241 20553 11253 20556
rect 11287 20553 11299 20587
rect 11241 20547 11299 20553
rect 6822 20448 6828 20460
rect 6196 20420 6828 20448
rect 5077 20411 5135 20417
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 9306 20448 9312 20460
rect 9267 20420 9312 20448
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 4433 20315 4491 20321
rect 4433 20281 4445 20315
rect 4479 20312 4491 20315
rect 4893 20315 4951 20321
rect 4893 20312 4905 20315
rect 4479 20284 4905 20312
rect 4479 20281 4491 20284
rect 4433 20275 4491 20281
rect 4893 20281 4905 20284
rect 4939 20312 4951 20315
rect 5258 20312 5264 20324
rect 4939 20284 5264 20312
rect 4939 20281 4951 20284
rect 4893 20275 4951 20281
rect 5258 20272 5264 20284
rect 5316 20312 5322 20324
rect 5810 20312 5816 20324
rect 5316 20284 5816 20312
rect 5316 20272 5322 20284
rect 5810 20272 5816 20284
rect 5868 20272 5874 20324
rect 7098 20321 7104 20324
rect 6641 20315 6699 20321
rect 6641 20281 6653 20315
rect 6687 20312 6699 20315
rect 7070 20315 7104 20321
rect 7070 20312 7082 20315
rect 6687 20284 7082 20312
rect 6687 20281 6699 20284
rect 6641 20275 6699 20281
rect 7070 20281 7082 20284
rect 7156 20312 7162 20324
rect 9217 20315 9275 20321
rect 7156 20284 7218 20312
rect 7070 20275 7104 20281
rect 7098 20272 7104 20275
rect 7156 20272 7162 20284
rect 9217 20281 9229 20315
rect 9263 20312 9275 20315
rect 9576 20315 9634 20321
rect 9576 20312 9588 20315
rect 9263 20284 9588 20312
rect 9263 20281 9275 20284
rect 9217 20275 9275 20281
rect 9576 20281 9588 20284
rect 9622 20312 9634 20315
rect 11146 20312 11152 20324
rect 9622 20284 11152 20312
rect 9622 20281 9634 20284
rect 9576 20275 9634 20281
rect 11146 20272 11152 20284
rect 11204 20272 11210 20324
rect 4522 20204 4528 20256
rect 4580 20244 4586 20256
rect 4982 20244 4988 20256
rect 4580 20216 4988 20244
rect 4580 20204 4586 20216
rect 4982 20204 4988 20216
rect 5040 20204 5046 20256
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 5994 20244 6000 20256
rect 5951 20216 6000 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 8202 20244 8208 20256
rect 8163 20216 8208 20244
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 10686 20244 10692 20256
rect 10647 20216 10692 20244
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 11514 20204 11520 20256
rect 11572 20244 11578 20256
rect 11609 20247 11667 20253
rect 11609 20244 11621 20247
rect 11572 20216 11621 20244
rect 11572 20204 11578 20216
rect 11609 20213 11621 20216
rect 11655 20213 11667 20247
rect 11609 20207 11667 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 4430 20000 4436 20052
rect 4488 20040 4494 20052
rect 4893 20043 4951 20049
rect 4893 20040 4905 20043
rect 4488 20012 4905 20040
rect 4488 20000 4494 20012
rect 4893 20009 4905 20012
rect 4939 20009 4951 20043
rect 4893 20003 4951 20009
rect 5905 20043 5963 20049
rect 5905 20009 5917 20043
rect 5951 20040 5963 20043
rect 6730 20040 6736 20052
rect 5951 20012 6736 20040
rect 5951 20009 5963 20012
rect 5905 20003 5963 20009
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 6822 20000 6828 20052
rect 6880 20040 6886 20052
rect 6917 20043 6975 20049
rect 6917 20040 6929 20043
rect 6880 20012 6929 20040
rect 6880 20000 6886 20012
rect 6917 20009 6929 20012
rect 6963 20009 6975 20043
rect 6917 20003 6975 20009
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9306 20040 9312 20052
rect 9171 20012 9312 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9306 20000 9312 20012
rect 9364 20000 9370 20052
rect 10318 20040 10324 20052
rect 10279 20012 10324 20040
rect 10318 20000 10324 20012
rect 10376 20000 10382 20052
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11112 20012 11897 20040
rect 11112 20000 11118 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 5994 19932 6000 19984
rect 6052 19972 6058 19984
rect 10772 19975 10830 19981
rect 6052 19944 6592 19972
rect 6052 19932 6058 19944
rect 6270 19904 6276 19916
rect 6231 19876 6276 19904
rect 6270 19864 6276 19876
rect 6328 19864 6334 19916
rect 6362 19864 6368 19916
rect 6420 19904 6426 19916
rect 6420 19876 6465 19904
rect 6420 19864 6426 19876
rect 6564 19845 6592 19944
rect 10772 19941 10784 19975
rect 10818 19972 10830 19975
rect 10962 19972 10968 19984
rect 10818 19944 10968 19972
rect 10818 19941 10830 19944
rect 10772 19935 10830 19941
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 10226 19864 10232 19916
rect 10284 19904 10290 19916
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 10284 19876 10517 19904
rect 10284 19864 10290 19876
rect 10505 19873 10517 19876
rect 10551 19904 10563 19907
rect 11514 19904 11520 19916
rect 10551 19876 11520 19904
rect 10551 19873 10563 19876
rect 10505 19867 10563 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19836 6607 19839
rect 8202 19836 8208 19848
rect 6595 19808 8208 19836
rect 6595 19805 6607 19808
rect 6549 19799 6607 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 12434 19796 12440 19848
rect 12492 19836 12498 19848
rect 12989 19839 13047 19845
rect 12989 19836 13001 19839
rect 12492 19808 13001 19836
rect 12492 19796 12498 19808
rect 12989 19805 13001 19808
rect 13035 19805 13047 19839
rect 12989 19799 13047 19805
rect 2590 19700 2596 19712
rect 2551 19672 2596 19700
rect 2590 19660 2596 19672
rect 2648 19660 2654 19712
rect 4430 19660 4436 19712
rect 4488 19700 4494 19712
rect 4525 19703 4583 19709
rect 4525 19700 4537 19703
rect 4488 19672 4537 19700
rect 4488 19660 4494 19672
rect 4525 19669 4537 19672
rect 4571 19669 4583 19703
rect 8662 19700 8668 19712
rect 8623 19672 8668 19700
rect 4525 19663 4583 19669
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 9493 19703 9551 19709
rect 9493 19669 9505 19703
rect 9539 19700 9551 19703
rect 9674 19700 9680 19712
rect 9539 19672 9680 19700
rect 9539 19669 9551 19672
rect 9493 19663 9551 19669
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 9858 19700 9864 19712
rect 9819 19672 9864 19700
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19700 12590 19712
rect 13538 19700 13544 19712
rect 12584 19672 13544 19700
rect 12584 19660 12590 19672
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 5629 19499 5687 19505
rect 5629 19465 5641 19499
rect 5675 19496 5687 19499
rect 5994 19496 6000 19508
rect 5675 19468 6000 19496
rect 5675 19465 5687 19468
rect 5629 19459 5687 19465
rect 5994 19456 6000 19468
rect 6052 19456 6058 19508
rect 9858 19388 9864 19440
rect 9916 19428 9922 19440
rect 10321 19431 10379 19437
rect 10321 19428 10333 19431
rect 9916 19400 10333 19428
rect 9916 19388 9922 19400
rect 10321 19397 10333 19400
rect 10367 19397 10379 19431
rect 10321 19391 10379 19397
rect 2590 19360 2596 19372
rect 2551 19332 2596 19360
rect 2590 19320 2596 19332
rect 2648 19320 2654 19372
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 9600 19332 10057 19360
rect 6362 19292 6368 19304
rect 6012 19264 6368 19292
rect 2501 19227 2559 19233
rect 2501 19193 2513 19227
rect 2547 19224 2559 19227
rect 2838 19227 2896 19233
rect 2838 19224 2850 19227
rect 2547 19196 2850 19224
rect 2547 19193 2559 19196
rect 2501 19187 2559 19193
rect 2838 19193 2850 19196
rect 2884 19224 2896 19227
rect 3510 19224 3516 19236
rect 2884 19196 3516 19224
rect 2884 19193 2896 19196
rect 2838 19187 2896 19193
rect 3510 19184 3516 19196
rect 3568 19184 3574 19236
rect 6012 19168 6040 19264
rect 6362 19252 6368 19264
rect 6420 19252 6426 19304
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 9600 19292 9628 19332
rect 10045 19329 10057 19332
rect 10091 19360 10103 19363
rect 10686 19360 10692 19372
rect 10091 19332 10692 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 10965 19363 11023 19369
rect 10965 19329 10977 19363
rect 11011 19360 11023 19363
rect 11146 19360 11152 19372
rect 11011 19332 11152 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12584 19332 12909 19360
rect 12584 19320 12590 19332
rect 12897 19329 12909 19332
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 9548 19264 9628 19292
rect 9769 19295 9827 19301
rect 9548 19252 9554 19264
rect 9769 19261 9781 19295
rect 9815 19292 9827 19295
rect 9858 19292 9864 19304
rect 9815 19264 9864 19292
rect 9815 19261 9827 19264
rect 9769 19255 9827 19261
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11333 19295 11391 19301
rect 11333 19292 11345 19295
rect 11112 19264 11345 19292
rect 11112 19252 11118 19264
rect 11333 19261 11345 19264
rect 11379 19292 11391 19295
rect 12618 19292 12624 19304
rect 11379 19264 12624 19292
rect 11379 19261 11391 19264
rect 11333 19255 11391 19261
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 6270 19184 6276 19236
rect 6328 19184 6334 19236
rect 7469 19227 7527 19233
rect 7469 19193 7481 19227
rect 7515 19224 7527 19227
rect 7561 19227 7619 19233
rect 7561 19224 7573 19227
rect 7515 19196 7573 19224
rect 7515 19193 7527 19196
rect 7469 19187 7527 19193
rect 7561 19193 7573 19196
rect 7607 19224 7619 19227
rect 7834 19224 7840 19236
rect 7607 19196 7840 19224
rect 7607 19193 7619 19196
rect 7561 19187 7619 19193
rect 7834 19184 7840 19196
rect 7892 19184 7898 19236
rect 10781 19227 10839 19233
rect 10781 19224 10793 19227
rect 10336 19196 10793 19224
rect 3970 19156 3976 19168
rect 3931 19128 3976 19156
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 5994 19156 6000 19168
rect 5955 19128 6000 19156
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 6288 19156 6316 19184
rect 10336 19168 10364 19196
rect 10781 19193 10793 19196
rect 10827 19193 10839 19227
rect 10781 19187 10839 19193
rect 12066 19184 12072 19236
rect 12124 19224 12130 19236
rect 12161 19227 12219 19233
rect 12161 19224 12173 19227
rect 12124 19196 12173 19224
rect 12124 19184 12130 19196
rect 12161 19193 12173 19196
rect 12207 19193 12219 19227
rect 13004 19224 13032 19323
rect 12161 19187 12219 19193
rect 12268 19196 13032 19224
rect 6365 19159 6423 19165
rect 6365 19156 6377 19159
rect 6288 19128 6377 19156
rect 6365 19125 6377 19128
rect 6411 19156 6423 19159
rect 6822 19156 6828 19168
rect 6411 19128 6828 19156
rect 6411 19125 6423 19128
rect 6365 19119 6423 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 8846 19156 8852 19168
rect 8444 19128 8852 19156
rect 8444 19116 8450 19128
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 9398 19156 9404 19168
rect 9359 19128 9404 19156
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 9732 19128 9873 19156
rect 9732 19116 9738 19128
rect 9861 19125 9873 19128
rect 9907 19125 9919 19159
rect 9861 19119 9919 19125
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10318 19156 10324 19168
rect 10100 19128 10324 19156
rect 10100 19116 10106 19128
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11793 19159 11851 19165
rect 11793 19156 11805 19159
rect 11112 19128 11805 19156
rect 11112 19116 11118 19128
rect 11793 19125 11805 19128
rect 11839 19156 11851 19159
rect 12268 19156 12296 19196
rect 11839 19128 12296 19156
rect 11839 19125 11851 19128
rect 11793 19119 11851 19125
rect 12342 19116 12348 19168
rect 12400 19156 12406 19168
rect 12437 19159 12495 19165
rect 12437 19156 12449 19159
rect 12400 19128 12449 19156
rect 12400 19116 12406 19128
rect 12437 19125 12449 19128
rect 12483 19125 12495 19159
rect 12437 19119 12495 19125
rect 12710 19116 12716 19168
rect 12768 19156 12774 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12768 19128 12817 19156
rect 12768 19116 12774 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 12805 19119 12863 19125
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 2590 18952 2596 18964
rect 2551 18924 2596 18952
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 6178 18912 6184 18964
rect 6236 18952 6242 18964
rect 6273 18955 6331 18961
rect 6273 18952 6285 18955
rect 6236 18924 6285 18952
rect 6236 18912 6242 18924
rect 6273 18921 6285 18924
rect 6319 18921 6331 18955
rect 7098 18952 7104 18964
rect 7059 18924 7104 18952
rect 6273 18915 6331 18921
rect 7098 18912 7104 18924
rect 7156 18952 7162 18964
rect 7650 18952 7656 18964
rect 7156 18924 7656 18952
rect 7156 18912 7162 18924
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 7929 18955 7987 18961
rect 7929 18921 7941 18955
rect 7975 18952 7987 18955
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 7975 18924 8493 18952
rect 7975 18921 7987 18924
rect 7929 18915 7987 18921
rect 8481 18921 8493 18924
rect 8527 18952 8539 18955
rect 9677 18955 9735 18961
rect 9677 18952 9689 18955
rect 8527 18924 9689 18952
rect 8527 18921 8539 18924
rect 8481 18915 8539 18921
rect 9677 18921 9689 18924
rect 9723 18921 9735 18955
rect 11146 18952 11152 18964
rect 11107 18924 11152 18952
rect 9677 18915 9735 18921
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 12066 18912 12072 18964
rect 12124 18952 12130 18964
rect 12710 18952 12716 18964
rect 12124 18924 12716 18952
rect 12124 18912 12130 18924
rect 12710 18912 12716 18924
rect 12768 18952 12774 18964
rect 13446 18952 13452 18964
rect 12768 18924 13452 18952
rect 12768 18912 12774 18924
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 1670 18884 1676 18896
rect 1631 18856 1676 18884
rect 1670 18844 1676 18856
rect 1728 18844 1734 18896
rect 5994 18844 6000 18896
rect 6052 18884 6058 18896
rect 6546 18884 6552 18896
rect 6052 18856 6552 18884
rect 6052 18844 6058 18856
rect 6546 18844 6552 18856
rect 6604 18844 6610 18896
rect 9490 18884 9496 18896
rect 9451 18856 9496 18884
rect 9490 18844 9496 18856
rect 9548 18844 9554 18896
rect 10045 18887 10103 18893
rect 10045 18853 10057 18887
rect 10091 18884 10103 18887
rect 10134 18884 10140 18896
rect 10091 18856 10140 18884
rect 10091 18853 10103 18856
rect 10045 18847 10103 18853
rect 10134 18844 10140 18856
rect 10192 18884 10198 18896
rect 11330 18884 11336 18896
rect 10192 18856 11336 18884
rect 10192 18844 10198 18856
rect 11330 18844 11336 18856
rect 11388 18844 11394 18896
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18785 1455 18819
rect 1397 18779 1455 18785
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18816 6239 18819
rect 6730 18816 6736 18828
rect 6227 18788 6736 18816
rect 6227 18785 6239 18788
rect 6181 18779 6239 18785
rect 1412 18748 1440 18779
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 8018 18776 8024 18828
rect 8076 18816 8082 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 8076 18788 8401 18816
rect 8076 18776 8082 18788
rect 8389 18785 8401 18788
rect 8435 18816 8447 18819
rect 8478 18816 8484 18828
rect 8435 18788 8484 18816
rect 8435 18785 8447 18788
rect 8389 18779 8447 18785
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 1670 18748 1676 18760
rect 1412 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 5994 18708 6000 18760
rect 6052 18748 6058 18760
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 6052 18720 6377 18748
rect 6052 18708 6058 18720
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 8570 18748 8576 18760
rect 8483 18720 8576 18748
rect 6365 18711 6423 18717
rect 8570 18708 8576 18720
rect 8628 18748 8634 18760
rect 9508 18748 9536 18844
rect 9858 18776 9864 18828
rect 9916 18776 9922 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11773 18819 11831 18825
rect 11773 18816 11785 18819
rect 11112 18788 11785 18816
rect 11112 18776 11118 18788
rect 11773 18785 11785 18788
rect 11819 18785 11831 18819
rect 11773 18779 11831 18785
rect 8628 18720 9536 18748
rect 9876 18748 9904 18776
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 9876 18720 10149 18748
rect 8628 18708 8634 18720
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 8021 18683 8079 18689
rect 8021 18649 8033 18683
rect 8067 18680 8079 18683
rect 8662 18680 8668 18692
rect 8067 18652 8668 18680
rect 8067 18649 8079 18652
rect 8021 18643 8079 18649
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 5534 18612 5540 18624
rect 5307 18584 5540 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 5810 18612 5816 18624
rect 5771 18584 5816 18612
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 7558 18612 7564 18624
rect 7519 18584 7564 18612
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 9125 18615 9183 18621
rect 9125 18581 9137 18615
rect 9171 18612 9183 18615
rect 9490 18612 9496 18624
rect 9171 18584 9496 18612
rect 9171 18581 9183 18584
rect 9125 18575 9183 18581
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 10152 18612 10180 18711
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 10321 18751 10379 18757
rect 10321 18748 10333 18751
rect 10284 18720 10333 18748
rect 10284 18708 10290 18720
rect 10321 18717 10333 18720
rect 10367 18748 10379 18751
rect 11146 18748 11152 18760
rect 10367 18720 11152 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 11514 18748 11520 18760
rect 11475 18720 11520 18748
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 10318 18612 10324 18624
rect 10152 18584 10324 18612
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 10686 18612 10692 18624
rect 10647 18584 10692 18612
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 12897 18615 12955 18621
rect 12897 18612 12909 18615
rect 12676 18584 12909 18612
rect 12676 18572 12682 18584
rect 12897 18581 12909 18584
rect 12943 18612 12955 18615
rect 12986 18612 12992 18624
rect 12943 18584 12992 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 3510 18368 3516 18420
rect 3568 18408 3574 18420
rect 3881 18411 3939 18417
rect 3881 18408 3893 18411
rect 3568 18380 3893 18408
rect 3568 18368 3574 18380
rect 3881 18377 3893 18380
rect 3927 18408 3939 18411
rect 4062 18408 4068 18420
rect 3927 18380 4068 18408
rect 3927 18377 3939 18380
rect 3881 18371 3939 18377
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18408 5135 18411
rect 5350 18408 5356 18420
rect 5123 18380 5356 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 6178 18408 6184 18420
rect 6139 18380 6184 18408
rect 6178 18368 6184 18380
rect 6236 18368 6242 18420
rect 8570 18408 8576 18420
rect 8531 18380 8576 18408
rect 8570 18368 8576 18380
rect 8628 18368 8634 18420
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 10318 18408 10324 18420
rect 9815 18380 10324 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 10318 18368 10324 18380
rect 10376 18408 10382 18420
rect 10962 18408 10968 18420
rect 10376 18380 10968 18408
rect 10376 18368 10382 18380
rect 10962 18368 10968 18380
rect 11020 18368 11026 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 11572 18380 13829 18408
rect 11572 18368 11578 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 13817 18371 13875 18377
rect 1670 18340 1676 18352
rect 1631 18312 1676 18340
rect 1670 18300 1676 18312
rect 1728 18300 1734 18352
rect 7098 18340 7104 18352
rect 7059 18312 7104 18340
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 8665 18343 8723 18349
rect 8665 18340 8677 18343
rect 7576 18312 8677 18340
rect 7576 18284 7604 18312
rect 8665 18309 8677 18312
rect 8711 18309 8723 18343
rect 8665 18303 8723 18309
rect 12066 18300 12072 18352
rect 12124 18340 12130 18352
rect 12161 18343 12219 18349
rect 12161 18340 12173 18343
rect 12124 18312 12173 18340
rect 12124 18300 12130 18312
rect 12161 18309 12173 18312
rect 12207 18340 12219 18343
rect 12894 18340 12900 18352
rect 12207 18312 12900 18340
rect 12207 18309 12219 18312
rect 12161 18303 12219 18309
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 5813 18275 5871 18281
rect 5813 18272 5825 18275
rect 4755 18244 5825 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 5813 18241 5825 18244
rect 5859 18272 5871 18275
rect 5994 18272 6000 18284
rect 5859 18244 6000 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 5994 18232 6000 18244
rect 6052 18232 6058 18284
rect 7558 18272 7564 18284
rect 7519 18244 7564 18272
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 7650 18232 7656 18284
rect 7708 18272 7714 18284
rect 7708 18244 7753 18272
rect 7708 18232 7714 18244
rect 8754 18232 8760 18284
rect 8812 18272 8818 18284
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 8812 18244 9229 18272
rect 8812 18232 8818 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 10870 18272 10876 18284
rect 10831 18244 10876 18272
rect 9217 18235 9275 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 12434 18232 12440 18284
rect 12492 18272 12498 18284
rect 13078 18272 13084 18284
rect 12492 18244 12848 18272
rect 13039 18244 13084 18272
rect 12492 18232 12498 18244
rect 2501 18207 2559 18213
rect 2501 18173 2513 18207
rect 2547 18204 2559 18207
rect 2590 18204 2596 18216
rect 2547 18176 2596 18204
rect 2547 18173 2559 18176
rect 2501 18167 2559 18173
rect 2590 18164 2596 18176
rect 2648 18164 2654 18216
rect 5350 18164 5356 18216
rect 5408 18204 5414 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 5408 18176 5641 18204
rect 5408 18164 5414 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 8662 18164 8668 18216
rect 8720 18204 8726 18216
rect 9033 18207 9091 18213
rect 9033 18204 9045 18207
rect 8720 18176 9045 18204
rect 8720 18164 8726 18176
rect 9033 18173 9045 18176
rect 9079 18173 9091 18207
rect 9033 18167 9091 18173
rect 9125 18207 9183 18213
rect 9125 18173 9137 18207
rect 9171 18204 9183 18207
rect 9398 18204 9404 18216
rect 9171 18176 9404 18204
rect 9171 18173 9183 18176
rect 9125 18167 9183 18173
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 10594 18204 10600 18216
rect 9548 18176 10600 18204
rect 9548 18164 9554 18176
rect 10594 18164 10600 18176
rect 10652 18204 10658 18216
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 10652 18176 10793 18204
rect 10652 18164 10658 18176
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12452 18204 12480 18232
rect 12820 18213 12848 18244
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 11931 18176 12480 18204
rect 12805 18207 12863 18213
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12805 18173 12817 18207
rect 12851 18173 12863 18207
rect 12805 18167 12863 18173
rect 2409 18139 2467 18145
rect 2409 18105 2421 18139
rect 2455 18136 2467 18139
rect 2746 18139 2804 18145
rect 2746 18136 2758 18139
rect 2455 18108 2758 18136
rect 2455 18105 2467 18108
rect 2409 18099 2467 18105
rect 2746 18105 2758 18108
rect 2792 18136 2804 18139
rect 4338 18136 4344 18148
rect 2792 18108 4344 18136
rect 2792 18105 2804 18108
rect 2746 18099 2804 18105
rect 4338 18096 4344 18108
rect 4396 18096 4402 18148
rect 5534 18136 5540 18148
rect 5495 18108 5540 18136
rect 5534 18096 5540 18108
rect 5592 18096 5598 18148
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 11146 18136 11152 18148
rect 10735 18108 11152 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 11146 18096 11152 18108
rect 11204 18136 11210 18148
rect 13449 18139 13507 18145
rect 13449 18136 13461 18139
rect 11204 18108 13461 18136
rect 11204 18096 11210 18108
rect 13449 18105 13461 18108
rect 13495 18105 13507 18139
rect 13449 18099 13507 18105
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18068 5227 18071
rect 5442 18068 5448 18080
rect 5215 18040 5448 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 6641 18071 6699 18077
rect 6641 18037 6653 18071
rect 6687 18068 6699 18071
rect 6730 18068 6736 18080
rect 6687 18040 6736 18068
rect 6687 18037 6699 18040
rect 6641 18031 6699 18037
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 8205 18071 8263 18077
rect 8205 18037 8217 18071
rect 8251 18068 8263 18071
rect 8478 18068 8484 18080
rect 8251 18040 8484 18068
rect 8251 18037 8263 18040
rect 8205 18031 8263 18037
rect 8478 18028 8484 18040
rect 8536 18068 8542 18080
rect 8662 18068 8668 18080
rect 8536 18040 8668 18068
rect 8536 18028 8542 18040
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 10134 18068 10140 18080
rect 10095 18040 10140 18068
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11425 18071 11483 18077
rect 11425 18068 11437 18071
rect 11112 18040 11437 18068
rect 11112 18028 11118 18040
rect 11425 18037 11437 18040
rect 11471 18037 11483 18071
rect 11425 18031 11483 18037
rect 12342 18028 12348 18080
rect 12400 18068 12406 18080
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 12400 18040 12449 18068
rect 12400 18028 12406 18040
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12894 18068 12900 18080
rect 12855 18040 12900 18068
rect 12437 18031 12495 18037
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 5166 17864 5172 17876
rect 3476 17836 5172 17864
rect 3476 17824 3482 17836
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 8205 17867 8263 17873
rect 8205 17864 8217 17867
rect 7708 17836 8217 17864
rect 7708 17824 7714 17836
rect 8205 17833 8217 17836
rect 8251 17833 8263 17867
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 8205 17827 8263 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 9916 17836 10149 17864
rect 9916 17824 9922 17836
rect 10137 17833 10149 17836
rect 10183 17833 10195 17867
rect 10137 17827 10195 17833
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 10870 17864 10876 17876
rect 10827 17836 10876 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11517 17867 11575 17873
rect 11517 17833 11529 17867
rect 11563 17864 11575 17867
rect 11977 17867 12035 17873
rect 11977 17864 11989 17867
rect 11563 17836 11989 17864
rect 11563 17833 11575 17836
rect 11517 17827 11575 17833
rect 11977 17833 11989 17836
rect 12023 17864 12035 17867
rect 12342 17864 12348 17876
rect 12023 17836 12348 17864
rect 12023 17833 12035 17836
rect 11977 17827 12035 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 3970 17756 3976 17808
rect 4028 17796 4034 17808
rect 4402 17799 4460 17805
rect 4402 17796 4414 17799
rect 4028 17768 4414 17796
rect 4028 17756 4034 17768
rect 4402 17765 4414 17768
rect 4448 17765 4460 17799
rect 9490 17796 9496 17808
rect 9403 17768 9496 17796
rect 4402 17759 4460 17765
rect 9490 17756 9496 17768
rect 9548 17796 9554 17808
rect 10226 17796 10232 17808
rect 9548 17768 10232 17796
rect 9548 17756 9554 17768
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 12066 17796 12072 17808
rect 11979 17768 12072 17796
rect 12066 17756 12072 17768
rect 12124 17796 12130 17808
rect 12250 17796 12256 17808
rect 12124 17768 12256 17796
rect 12124 17756 12130 17768
rect 12250 17756 12256 17768
rect 12308 17756 12314 17808
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 2774 17728 2780 17740
rect 2363 17700 2780 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 2774 17688 2780 17700
rect 2832 17728 2838 17740
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17660 3111 17663
rect 3326 17660 3332 17672
rect 3099 17632 3332 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 3326 17620 3332 17632
rect 3384 17660 3390 17672
rect 3988 17660 4016 17756
rect 7092 17731 7150 17737
rect 7092 17697 7104 17731
rect 7138 17728 7150 17731
rect 7374 17728 7380 17740
rect 7138 17700 7380 17728
rect 7138 17697 7150 17700
rect 7092 17691 7150 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 9306 17688 9312 17740
rect 9364 17728 9370 17740
rect 9766 17728 9772 17740
rect 9364 17700 9772 17728
rect 9364 17688 9370 17700
rect 9766 17688 9772 17700
rect 9824 17728 9830 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9824 17700 10057 17728
rect 9824 17688 9830 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 3384 17632 4016 17660
rect 4157 17663 4215 17669
rect 3384 17620 3390 17632
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 6822 17660 6828 17672
rect 6783 17632 6828 17660
rect 4157 17623 4215 17629
rect 2590 17552 2596 17604
rect 2648 17592 2654 17604
rect 3418 17592 3424 17604
rect 2648 17564 3424 17592
rect 2648 17552 2654 17564
rect 3418 17552 3424 17564
rect 3476 17592 3482 17604
rect 4172 17592 4200 17623
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 10244 17669 10272 17756
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 12250 17660 12256 17672
rect 12163 17632 12256 17660
rect 10229 17623 10287 17629
rect 12250 17620 12256 17632
rect 12308 17660 12314 17672
rect 12986 17660 12992 17672
rect 12308 17632 12992 17660
rect 12308 17620 12314 17632
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 3476 17564 4200 17592
rect 3476 17552 3482 17564
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 11609 17595 11667 17601
rect 11609 17592 11621 17595
rect 11204 17564 11621 17592
rect 11204 17552 11210 17564
rect 11609 17561 11621 17564
rect 11655 17561 11667 17595
rect 13078 17592 13084 17604
rect 11609 17555 11667 17561
rect 12728 17564 13084 17592
rect 12728 17536 12756 17564
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 1854 17484 1860 17536
rect 1912 17524 1918 17536
rect 2409 17527 2467 17533
rect 2409 17524 2421 17527
rect 1912 17496 2421 17524
rect 1912 17484 1918 17496
rect 2409 17493 2421 17496
rect 2455 17493 2467 17527
rect 3510 17524 3516 17536
rect 3471 17496 3516 17524
rect 2409 17487 2467 17493
rect 3510 17484 3516 17496
rect 3568 17484 3574 17536
rect 5537 17527 5595 17533
rect 5537 17493 5549 17527
rect 5583 17524 5595 17527
rect 5994 17524 6000 17536
rect 5583 17496 6000 17524
rect 5583 17493 5595 17496
rect 5537 17487 5595 17493
rect 5994 17484 6000 17496
rect 6052 17524 6058 17536
rect 6089 17527 6147 17533
rect 6089 17524 6101 17527
rect 6052 17496 6101 17524
rect 6052 17484 6058 17496
rect 6089 17493 6101 17496
rect 6135 17493 6147 17527
rect 6089 17487 6147 17493
rect 6733 17527 6791 17533
rect 6733 17493 6745 17527
rect 6779 17524 6791 17527
rect 7466 17524 7472 17536
rect 6779 17496 7472 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 8754 17524 8760 17536
rect 8715 17496 8760 17524
rect 8754 17484 8760 17496
rect 8812 17484 8818 17536
rect 11054 17524 11060 17536
rect 11015 17496 11060 17524
rect 11054 17484 11060 17496
rect 11112 17524 11118 17536
rect 12710 17524 12716 17536
rect 11112 17496 12716 17524
rect 11112 17484 11118 17496
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 12802 17484 12808 17536
rect 12860 17524 12866 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 12860 17496 13001 17524
rect 12860 17484 12866 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 3421 17323 3479 17329
rect 3421 17320 3433 17323
rect 2832 17292 3433 17320
rect 2832 17280 2838 17292
rect 3421 17289 3433 17292
rect 3467 17289 3479 17323
rect 4890 17320 4896 17332
rect 4851 17292 4896 17320
rect 3421 17283 3479 17289
rect 4890 17280 4896 17292
rect 4948 17280 4954 17332
rect 7466 17280 7472 17332
rect 7524 17320 7530 17332
rect 8113 17323 8171 17329
rect 8113 17320 8125 17323
rect 7524 17292 8125 17320
rect 7524 17280 7530 17292
rect 8113 17289 8125 17292
rect 8159 17289 8171 17323
rect 8113 17283 8171 17289
rect 9401 17323 9459 17329
rect 9401 17289 9413 17323
rect 9447 17320 9459 17323
rect 9490 17320 9496 17332
rect 9447 17292 9496 17320
rect 9447 17289 9459 17292
rect 9401 17283 9459 17289
rect 9490 17280 9496 17292
rect 9548 17280 9554 17332
rect 9769 17323 9827 17329
rect 9769 17289 9781 17323
rect 9815 17320 9827 17323
rect 9858 17320 9864 17332
rect 9815 17292 9864 17320
rect 9815 17289 9827 17292
rect 9769 17283 9827 17289
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10686 17320 10692 17332
rect 10599 17292 10692 17320
rect 10686 17280 10692 17292
rect 10744 17320 10750 17332
rect 11146 17320 11152 17332
rect 10744 17292 11152 17320
rect 10744 17280 10750 17292
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 11885 17323 11943 17329
rect 11885 17289 11897 17323
rect 11931 17320 11943 17323
rect 12250 17320 12256 17332
rect 11931 17292 12256 17320
rect 11931 17289 11943 17292
rect 11885 17283 11943 17289
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12492 17292 12537 17320
rect 12492 17280 12498 17292
rect 2501 17255 2559 17261
rect 2501 17221 2513 17255
rect 2547 17252 2559 17255
rect 3326 17252 3332 17264
rect 2547 17224 3332 17252
rect 2547 17221 2559 17224
rect 2501 17215 2559 17221
rect 3326 17212 3332 17224
rect 3384 17212 3390 17264
rect 4985 17255 5043 17261
rect 4985 17252 4997 17255
rect 3896 17224 4997 17252
rect 1578 17184 1584 17196
rect 1539 17156 1584 17184
rect 1578 17144 1584 17156
rect 1636 17144 1642 17196
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 3896 17193 3924 17224
rect 4985 17221 4997 17224
rect 5031 17221 5043 17255
rect 4985 17215 5043 17221
rect 6086 17212 6092 17264
rect 6144 17252 6150 17264
rect 6730 17252 6736 17264
rect 6144 17224 6736 17252
rect 6144 17212 6150 17224
rect 6730 17212 6736 17224
rect 6788 17212 6794 17264
rect 10781 17255 10839 17261
rect 10781 17221 10793 17255
rect 10827 17252 10839 17255
rect 12802 17252 12808 17264
rect 10827 17224 12808 17252
rect 10827 17221 10839 17224
rect 10781 17215 10839 17221
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 3881 17187 3939 17193
rect 3881 17184 3893 17187
rect 3568 17156 3893 17184
rect 3568 17144 3574 17156
rect 3881 17153 3893 17156
rect 3927 17153 3939 17187
rect 4062 17184 4068 17196
rect 4023 17156 4068 17184
rect 3881 17147 3939 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4338 17144 4344 17196
rect 4396 17184 4402 17196
rect 5537 17187 5595 17193
rect 5537 17184 5549 17187
rect 4396 17156 5549 17184
rect 4396 17144 4402 17156
rect 5537 17153 5549 17156
rect 5583 17153 5595 17187
rect 7374 17184 7380 17196
rect 7287 17156 7380 17184
rect 5537 17147 5595 17153
rect 7374 17144 7380 17156
rect 7432 17184 7438 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7432 17156 8033 17184
rect 7432 17144 7438 17156
rect 8021 17153 8033 17156
rect 8067 17184 8079 17187
rect 8754 17184 8760 17196
rect 8067 17156 8760 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11020 17156 11345 17184
rect 11020 17144 11026 17156
rect 11333 17153 11345 17156
rect 11379 17153 11391 17187
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 11333 17147 11391 17153
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 1394 17116 1400 17128
rect 1355 17088 1400 17116
rect 1394 17076 1400 17088
rect 1452 17076 1458 17128
rect 4890 17076 4896 17128
rect 4948 17116 4954 17128
rect 5353 17119 5411 17125
rect 5353 17116 5365 17119
rect 4948 17088 5365 17116
rect 4948 17076 4954 17088
rect 5353 17085 5365 17088
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 10778 17116 10784 17128
rect 10468 17088 10784 17116
rect 10468 17076 10474 17088
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 11112 17088 11253 17116
rect 11112 17076 11118 17088
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 12802 17116 12808 17128
rect 12763 17088 12808 17116
rect 11241 17079 11299 17085
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 2961 17051 3019 17057
rect 2961 17017 2973 17051
rect 3007 17048 3019 17051
rect 3789 17051 3847 17057
rect 3789 17048 3801 17051
rect 3007 17020 3801 17048
rect 3007 17017 3019 17020
rect 2961 17011 3019 17017
rect 3789 17017 3801 17020
rect 3835 17048 3847 17051
rect 4154 17048 4160 17060
rect 3835 17020 4160 17048
rect 3835 17017 3847 17020
rect 3789 17011 3847 17017
rect 4154 17008 4160 17020
rect 4212 17008 4218 17060
rect 4522 17008 4528 17060
rect 4580 17048 4586 17060
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 4580 17020 6837 17048
rect 4580 17008 4586 17020
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 9490 17008 9496 17060
rect 9548 17048 9554 17060
rect 9766 17048 9772 17060
rect 9548 17020 9772 17048
rect 9548 17008 9554 17020
rect 9766 17008 9772 17020
rect 9824 17048 9830 17060
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 9824 17020 10057 17048
rect 9824 17008 9830 17020
rect 10045 17017 10057 17020
rect 10091 17017 10103 17051
rect 10045 17011 10103 17017
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 4304 16952 4445 16980
rect 4304 16940 4310 16952
rect 4433 16949 4445 16952
rect 4479 16980 4491 16983
rect 5442 16980 5448 16992
rect 4479 16952 5448 16980
rect 4479 16949 4491 16952
rect 4433 16943 4491 16949
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 6086 16940 6092 16992
rect 6144 16980 6150 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6144 16952 6561 16980
rect 6144 16940 6150 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 8478 16980 8484 16992
rect 8439 16952 8484 16980
rect 6549 16943 6607 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 8573 16983 8631 16989
rect 8573 16949 8585 16983
rect 8619 16980 8631 16983
rect 8846 16980 8852 16992
rect 8619 16952 8852 16980
rect 8619 16949 8631 16952
rect 8573 16943 8631 16949
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16980 12958 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 12952 16952 13461 16980
rect 12952 16940 12958 16952
rect 13449 16949 13461 16952
rect 13495 16949 13507 16983
rect 13449 16943 13507 16949
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 1581 16779 1639 16785
rect 1581 16776 1593 16779
rect 1452 16748 1593 16776
rect 1452 16736 1458 16748
rect 1581 16745 1593 16748
rect 1627 16745 1639 16779
rect 1581 16739 1639 16745
rect 2317 16779 2375 16785
rect 2317 16745 2329 16779
rect 2363 16776 2375 16779
rect 2409 16779 2467 16785
rect 2409 16776 2421 16779
rect 2363 16748 2421 16776
rect 2363 16745 2375 16748
rect 2317 16739 2375 16745
rect 2409 16745 2421 16748
rect 2455 16776 2467 16779
rect 2866 16776 2872 16788
rect 2455 16748 2872 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 3697 16779 3755 16785
rect 3697 16776 3709 16779
rect 3476 16748 3709 16776
rect 3476 16736 3482 16748
rect 3697 16745 3709 16748
rect 3743 16776 3755 16779
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3743 16748 3801 16776
rect 3743 16745 3755 16748
rect 3697 16739 3755 16745
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 4154 16776 4160 16788
rect 4115 16748 4160 16776
rect 3789 16739 3847 16745
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 4522 16776 4528 16788
rect 4483 16748 4528 16776
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 4617 16779 4675 16785
rect 4617 16745 4629 16779
rect 4663 16776 4675 16779
rect 4798 16776 4804 16788
rect 4663 16748 4804 16776
rect 4663 16745 4675 16748
rect 4617 16739 4675 16745
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 5534 16776 5540 16788
rect 5495 16748 5540 16776
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 6086 16776 6092 16788
rect 5736 16748 6092 16776
rect 3513 16711 3571 16717
rect 3513 16677 3525 16711
rect 3559 16708 3571 16711
rect 4062 16708 4068 16720
rect 3559 16680 4068 16708
rect 3559 16677 3571 16680
rect 3513 16671 3571 16677
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3234 16640 3240 16652
rect 2823 16612 3240 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 2866 16572 2872 16584
rect 2827 16544 2872 16572
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 3053 16575 3111 16581
rect 3053 16572 3065 16575
rect 3016 16544 3065 16572
rect 3016 16532 3022 16544
rect 3053 16541 3065 16544
rect 3099 16572 3111 16575
rect 3528 16572 3556 16671
rect 4062 16668 4068 16680
rect 4120 16668 4126 16720
rect 5736 16649 5764 16748
rect 6086 16736 6092 16748
rect 6144 16776 6150 16788
rect 6822 16776 6828 16788
rect 6144 16748 6828 16776
rect 6144 16736 6150 16748
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7837 16779 7895 16785
rect 7837 16745 7849 16779
rect 7883 16776 7895 16779
rect 8018 16776 8024 16788
rect 7883 16748 8024 16776
rect 7883 16745 7895 16748
rect 7837 16739 7895 16745
rect 8018 16736 8024 16748
rect 8076 16776 8082 16788
rect 8478 16776 8484 16788
rect 8076 16748 8484 16776
rect 8076 16736 8082 16748
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 9398 16776 9404 16788
rect 8803 16748 9404 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 10410 16776 10416 16788
rect 10371 16748 10416 16776
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 11885 16779 11943 16785
rect 11885 16745 11897 16779
rect 11931 16776 11943 16779
rect 12066 16776 12072 16788
rect 11931 16748 12072 16776
rect 11931 16745 11943 16748
rect 11885 16739 11943 16745
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 12768 16748 13369 16776
rect 12768 16736 12774 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 13357 16739 13415 16745
rect 5994 16717 6000 16720
rect 5988 16708 6000 16717
rect 5907 16680 6000 16708
rect 5988 16671 6000 16680
rect 6052 16708 6058 16720
rect 6178 16708 6184 16720
rect 6052 16680 6184 16708
rect 5994 16668 6000 16671
rect 6052 16668 6058 16680
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 10873 16711 10931 16717
rect 10873 16708 10885 16711
rect 10336 16680 10885 16708
rect 10336 16652 10364 16680
rect 10873 16677 10885 16680
rect 10919 16677 10931 16711
rect 10873 16671 10931 16677
rect 3697 16643 3755 16649
rect 3697 16609 3709 16643
rect 3743 16640 3755 16643
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 3743 16612 5733 16640
rect 3743 16609 3755 16612
rect 3697 16603 3755 16609
rect 5721 16609 5733 16612
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8846 16640 8852 16652
rect 8251 16612 8852 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 8846 16600 8852 16612
rect 8904 16600 8910 16652
rect 10318 16640 10324 16652
rect 10279 16612 10324 16640
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10781 16643 10839 16649
rect 10781 16609 10793 16643
rect 10827 16609 10839 16643
rect 10781 16603 10839 16609
rect 3099 16544 3556 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4709 16575 4767 16581
rect 4709 16572 4721 16575
rect 4396 16544 4721 16572
rect 4396 16532 4402 16544
rect 4709 16541 4721 16544
rect 4755 16572 4767 16575
rect 4982 16572 4988 16584
rect 4755 16544 4988 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4982 16532 4988 16544
rect 5040 16572 5046 16584
rect 5169 16575 5227 16581
rect 5169 16572 5181 16575
rect 5040 16544 5181 16572
rect 5040 16532 5046 16544
rect 5169 16541 5181 16544
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10042 16572 10048 16584
rect 9999 16544 10048 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10042 16532 10048 16544
rect 10100 16572 10106 16584
rect 10796 16572 10824 16603
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 11112 16612 11437 16640
rect 11112 16600 11118 16612
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 12066 16600 12072 16652
rect 12124 16640 12130 16652
rect 12233 16643 12291 16649
rect 12233 16640 12245 16643
rect 12124 16612 12245 16640
rect 12124 16600 12130 16612
rect 12233 16609 12245 16612
rect 12279 16609 12291 16643
rect 12233 16603 12291 16609
rect 10962 16572 10968 16584
rect 10100 16544 10824 16572
rect 10923 16544 10968 16572
rect 10100 16532 10106 16544
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11882 16532 11888 16584
rect 11940 16572 11946 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11940 16544 11989 16572
rect 11940 16532 11946 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 5994 16396 6000 16448
rect 6052 16436 6058 16448
rect 7101 16439 7159 16445
rect 7101 16436 7113 16439
rect 6052 16408 7113 16436
rect 6052 16396 6058 16408
rect 7101 16405 7113 16408
rect 7147 16405 7159 16439
rect 7101 16399 7159 16405
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 12894 16436 12900 16448
rect 11204 16408 12900 16436
rect 11204 16396 11210 16408
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 4522 16232 4528 16244
rect 4483 16204 4528 16232
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 4982 16232 4988 16244
rect 4943 16204 4988 16232
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 6546 16192 6552 16244
rect 6604 16232 6610 16244
rect 6822 16232 6828 16244
rect 6604 16204 6828 16232
rect 6604 16192 6610 16204
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7009 16235 7067 16241
rect 7009 16232 7021 16235
rect 6972 16204 7021 16232
rect 6972 16192 6978 16204
rect 7009 16201 7021 16204
rect 7055 16201 7067 16235
rect 7009 16195 7067 16201
rect 8754 16192 8760 16244
rect 8812 16232 8818 16244
rect 9125 16235 9183 16241
rect 9125 16232 9137 16235
rect 8812 16204 9137 16232
rect 8812 16192 8818 16204
rect 9125 16201 9137 16204
rect 9171 16201 9183 16235
rect 9125 16195 9183 16201
rect 10781 16235 10839 16241
rect 10781 16201 10793 16235
rect 10827 16232 10839 16235
rect 11054 16232 11060 16244
rect 10827 16204 11060 16232
rect 10827 16201 10839 16204
rect 10781 16195 10839 16201
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 12066 16232 12072 16244
rect 12027 16204 12072 16232
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 4798 16164 4804 16176
rect 4295 16136 4804 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 9953 16167 10011 16173
rect 9953 16133 9965 16167
rect 9999 16164 10011 16167
rect 10962 16164 10968 16176
rect 9999 16136 10968 16164
rect 9999 16133 10011 16136
rect 9953 16127 10011 16133
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 2958 16096 2964 16108
rect 2547 16068 2964 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 2958 16056 2964 16068
rect 3016 16056 3022 16108
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 5629 16099 5687 16105
rect 5629 16096 5641 16099
rect 5592 16068 5641 16096
rect 5592 16056 5598 16068
rect 5629 16065 5641 16068
rect 5675 16065 5687 16099
rect 5629 16059 5687 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 5994 16096 6000 16108
rect 5859 16068 6000 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16096 7711 16099
rect 11425 16099 11483 16105
rect 7699 16068 7880 16096
rect 7699 16065 7711 16068
rect 7653 16059 7711 16065
rect 7742 16028 7748 16040
rect 7703 16000 7748 16028
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 7852 16028 7880 16068
rect 11425 16065 11437 16099
rect 11471 16096 11483 16099
rect 12066 16096 12072 16108
rect 11471 16068 12072 16096
rect 11471 16065 11483 16068
rect 11425 16059 11483 16065
rect 12066 16056 12072 16068
rect 12124 16056 12130 16108
rect 8012 16031 8070 16037
rect 8012 16028 8024 16031
rect 7852 16000 8024 16028
rect 8012 15997 8024 16000
rect 8058 16028 8070 16031
rect 8570 16028 8576 16040
rect 8058 16000 8576 16028
rect 8058 15997 8070 16000
rect 8012 15991 8070 15997
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 9732 16000 10333 16028
rect 9732 15988 9738 16000
rect 10321 15997 10333 16000
rect 10367 16028 10379 16031
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10367 16000 11161 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 11149 15997 11161 16000
rect 11195 16028 11207 16031
rect 11330 16028 11336 16040
rect 11195 16000 11336 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 11882 15988 11888 16040
rect 11940 15988 11946 16040
rect 5537 15963 5595 15969
rect 5537 15929 5549 15963
rect 5583 15960 5595 15963
rect 5810 15960 5816 15972
rect 5583 15932 5816 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 5810 15920 5816 15932
rect 5868 15960 5874 15972
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 5868 15932 6561 15960
rect 5868 15920 5874 15932
rect 6549 15929 6561 15932
rect 6595 15929 6607 15963
rect 10594 15960 10600 15972
rect 10555 15932 10600 15960
rect 6549 15923 6607 15929
rect 10594 15920 10600 15932
rect 10652 15960 10658 15972
rect 11241 15963 11299 15969
rect 11241 15960 11253 15963
rect 10652 15932 11253 15960
rect 10652 15920 10658 15932
rect 11241 15929 11253 15932
rect 11287 15929 11299 15963
rect 11241 15923 11299 15929
rect 2590 15852 2596 15904
rect 2648 15892 2654 15904
rect 2866 15892 2872 15904
rect 2648 15864 2872 15892
rect 2648 15852 2654 15864
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 3234 15892 3240 15904
rect 3147 15864 3240 15892
rect 3234 15852 3240 15864
rect 3292 15892 3298 15904
rect 4062 15892 4068 15904
rect 3292 15864 4068 15892
rect 3292 15852 3298 15864
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5442 15892 5448 15904
rect 5215 15864 5448 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 6178 15892 6184 15904
rect 6139 15864 6184 15892
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 11330 15852 11336 15904
rect 11388 15892 11394 15904
rect 11900 15892 11928 15988
rect 12621 15895 12679 15901
rect 12621 15892 12633 15895
rect 11388 15864 12633 15892
rect 11388 15852 11394 15864
rect 12621 15861 12633 15864
rect 12667 15861 12679 15895
rect 12621 15855 12679 15861
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15688 5319 15691
rect 5994 15688 6000 15700
rect 5307 15660 6000 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 7742 15688 7748 15700
rect 7703 15660 7748 15688
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 8018 15688 8024 15700
rect 7979 15660 8024 15688
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 9033 15691 9091 15697
rect 9033 15688 9045 15691
rect 8628 15660 9045 15688
rect 8628 15648 8634 15660
rect 9033 15657 9045 15660
rect 9079 15657 9091 15691
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 9033 15651 9091 15657
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10505 15691 10563 15697
rect 10505 15657 10517 15691
rect 10551 15688 10563 15691
rect 10686 15688 10692 15700
rect 10551 15660 10692 15688
rect 10551 15657 10563 15660
rect 10505 15651 10563 15657
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 11149 15691 11207 15697
rect 11149 15657 11161 15691
rect 11195 15688 11207 15691
rect 12066 15688 12072 15700
rect 11195 15660 12072 15688
rect 11195 15657 11207 15660
rect 11149 15651 11207 15657
rect 11164 15620 11192 15651
rect 12066 15648 12072 15660
rect 12124 15688 12130 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 12124 15660 13001 15688
rect 12124 15648 12130 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 12989 15651 13047 15657
rect 11072 15592 11192 15620
rect 5902 15512 5908 15564
rect 5960 15552 5966 15564
rect 5997 15555 6055 15561
rect 5997 15552 6009 15555
rect 5960 15524 6009 15552
rect 5960 15512 5966 15524
rect 5997 15521 6009 15524
rect 6043 15552 6055 15555
rect 7282 15552 7288 15564
rect 6043 15524 7288 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 8386 15552 8392 15564
rect 8347 15524 8392 15552
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 10410 15552 10416 15564
rect 8536 15524 8581 15552
rect 10371 15524 10416 15552
rect 8536 15512 8542 15524
rect 10410 15512 10416 15524
rect 10468 15512 10474 15564
rect 5166 15444 5172 15496
rect 5224 15484 5230 15496
rect 6086 15484 6092 15496
rect 5224 15456 6092 15484
rect 5224 15444 5230 15456
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 6273 15487 6331 15493
rect 6273 15484 6285 15487
rect 6236 15456 6285 15484
rect 6236 15444 6242 15456
rect 6273 15453 6285 15456
rect 6319 15484 6331 15487
rect 6362 15484 6368 15496
rect 6319 15456 6368 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8496 15484 8524 15512
rect 11072 15496 11100 15592
rect 11146 15512 11152 15564
rect 11204 15552 11210 15564
rect 11865 15555 11923 15561
rect 11865 15552 11877 15555
rect 11204 15524 11877 15552
rect 11204 15512 11210 15524
rect 11865 15521 11877 15524
rect 11911 15521 11923 15555
rect 11865 15515 11923 15521
rect 8260 15456 8524 15484
rect 8260 15444 8266 15456
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 10689 15487 10747 15493
rect 8628 15456 8673 15484
rect 8628 15444 8634 15456
rect 10689 15453 10701 15487
rect 10735 15484 10747 15487
rect 11054 15484 11060 15496
rect 10735 15456 11060 15484
rect 10735 15453 10747 15456
rect 10689 15447 10747 15453
rect 8478 15376 8484 15428
rect 8536 15416 8542 15428
rect 9582 15416 9588 15428
rect 8536 15388 9588 15416
rect 8536 15376 8542 15388
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 9953 15419 10011 15425
rect 9953 15385 9965 15419
rect 9999 15416 10011 15419
rect 10704 15416 10732 15447
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 11609 15487 11667 15493
rect 11609 15484 11621 15487
rect 11388 15456 11621 15484
rect 11388 15444 11394 15456
rect 11609 15453 11621 15456
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 9999 15388 10732 15416
rect 9999 15385 10011 15388
rect 9953 15379 10011 15385
rect 5626 15348 5632 15360
rect 5587 15320 5632 15348
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 5902 15104 5908 15156
rect 5960 15144 5966 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5960 15116 6009 15144
rect 5960 15104 5966 15116
rect 5997 15113 6009 15116
rect 6043 15113 6055 15147
rect 6362 15144 6368 15156
rect 6323 15116 6368 15144
rect 5997 15107 6055 15113
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 8113 15147 8171 15153
rect 8113 15113 8125 15147
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8573 15147 8631 15153
rect 8573 15144 8585 15147
rect 8352 15116 8585 15144
rect 8352 15104 8358 15116
rect 8573 15113 8585 15116
rect 8619 15144 8631 15147
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8619 15116 8677 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8846 15144 8852 15156
rect 8807 15116 8852 15144
rect 8665 15107 8723 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 10376 15116 10425 15144
rect 10376 15104 10382 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 10413 15107 10471 15113
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 9953 15079 10011 15085
rect 9953 15076 9965 15079
rect 9824 15048 9965 15076
rect 9824 15036 9830 15048
rect 9953 15045 9965 15048
rect 9999 15076 10011 15079
rect 10686 15076 10692 15088
rect 9999 15048 10692 15076
rect 9999 15045 10011 15048
rect 9953 15039 10011 15045
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 1578 15008 1584 15020
rect 1539 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 8570 15008 8576 15020
rect 8352 14980 8576 15008
rect 8352 14968 8358 14980
rect 8570 14968 8576 14980
rect 8628 15008 8634 15020
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 8628 14980 9413 15008
rect 8628 14968 8634 14980
rect 9401 14977 9413 14980
rect 9447 14977 9459 15011
rect 11054 15008 11060 15020
rect 11015 14980 11060 15008
rect 9401 14971 9459 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1762 14940 1768 14952
rect 1443 14912 1768 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 6086 14940 6092 14952
rect 5767 14912 6092 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 6086 14900 6092 14912
rect 6144 14940 6150 14952
rect 8846 14940 8852 14952
rect 6144 14912 8852 14940
rect 6144 14900 6150 14912
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9364 14912 9409 14940
rect 9364 14900 9370 14912
rect 8573 14875 8631 14881
rect 8573 14841 8585 14875
rect 8619 14872 8631 14875
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 8619 14844 9229 14872
rect 8619 14841 8631 14844
rect 8573 14835 8631 14841
rect 9217 14841 9229 14844
rect 9263 14872 9275 14875
rect 9582 14872 9588 14884
rect 9263 14844 9588 14872
rect 9263 14841 9275 14844
rect 9217 14835 9275 14841
rect 9582 14832 9588 14844
rect 9640 14832 9646 14884
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 10060 14844 10793 14872
rect 10060 14816 10088 14844
rect 10781 14841 10793 14844
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 11330 14832 11336 14884
rect 11388 14872 11394 14884
rect 11977 14875 12035 14881
rect 11977 14872 11989 14875
rect 11388 14844 11989 14872
rect 11388 14832 11394 14844
rect 11977 14841 11989 14844
rect 12023 14841 12035 14875
rect 11977 14835 12035 14841
rect 2498 14804 2504 14816
rect 2459 14776 2504 14804
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 10226 14804 10232 14816
rect 10187 14776 10232 14804
rect 10226 14764 10232 14776
rect 10284 14804 10290 14816
rect 10873 14807 10931 14813
rect 10873 14804 10885 14807
rect 10284 14776 10885 14804
rect 10284 14764 10290 14776
rect 10873 14773 10885 14776
rect 10919 14773 10931 14807
rect 10873 14767 10931 14773
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11609 14807 11667 14813
rect 11609 14804 11621 14807
rect 11204 14776 11621 14804
rect 11204 14764 11210 14776
rect 11609 14773 11621 14776
rect 11655 14773 11667 14807
rect 11609 14767 11667 14773
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2590 14600 2596 14612
rect 2455 14572 2596 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 3418 14600 3424 14612
rect 3379 14572 3424 14600
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 4062 14600 4068 14612
rect 4023 14572 4068 14600
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 4706 14600 4712 14612
rect 4479 14572 4712 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 5626 14560 5632 14612
rect 5684 14600 5690 14612
rect 6089 14603 6147 14609
rect 6089 14600 6101 14603
rect 5684 14572 6101 14600
rect 5684 14560 5690 14572
rect 6089 14569 6101 14572
rect 6135 14569 6147 14603
rect 8294 14600 8300 14612
rect 8255 14572 8300 14600
rect 6089 14563 6147 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9306 14600 9312 14612
rect 8987 14572 9312 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 5810 14532 5816 14544
rect 5592 14504 5816 14532
rect 5592 14492 5598 14504
rect 5810 14492 5816 14504
rect 5868 14532 5874 14544
rect 5997 14535 6055 14541
rect 5997 14532 6009 14535
rect 5868 14504 6009 14532
rect 5868 14492 5874 14504
rect 5997 14501 6009 14504
rect 6043 14501 6055 14535
rect 5997 14495 6055 14501
rect 7650 14492 7656 14544
rect 7708 14532 7714 14544
rect 8956 14532 8984 14563
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9674 14600 9680 14612
rect 9635 14572 9680 14600
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 11149 14603 11207 14609
rect 11149 14600 11161 14603
rect 11112 14572 11161 14600
rect 11112 14560 11118 14572
rect 11149 14569 11161 14572
rect 11195 14569 11207 14603
rect 11149 14563 11207 14569
rect 13538 14532 13544 14544
rect 7708 14504 8984 14532
rect 13499 14504 13544 14532
rect 7708 14492 7714 14504
rect 13538 14492 13544 14504
rect 13596 14492 13602 14544
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 3234 14464 3240 14476
rect 2832 14436 2877 14464
rect 3068 14436 3240 14464
rect 2832 14424 2838 14436
rect 2498 14356 2504 14408
rect 2556 14396 2562 14408
rect 3068 14405 3096 14436
rect 3234 14424 3240 14436
rect 3292 14464 3298 14476
rect 4338 14464 4344 14476
rect 3292 14436 4344 14464
rect 3292 14424 3298 14436
rect 4338 14424 4344 14436
rect 4396 14464 4402 14476
rect 4396 14436 4660 14464
rect 4396 14424 4402 14436
rect 2869 14399 2927 14405
rect 2869 14396 2881 14399
rect 2556 14368 2881 14396
rect 2556 14356 2562 14368
rect 2869 14365 2881 14368
rect 2915 14365 2927 14399
rect 2869 14359 2927 14365
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14365 3111 14399
rect 3053 14359 3111 14365
rect 3881 14399 3939 14405
rect 3881 14365 3893 14399
rect 3927 14396 3939 14399
rect 4062 14396 4068 14408
rect 3927 14368 4068 14396
rect 3927 14365 3939 14368
rect 3881 14359 3939 14365
rect 1946 14288 1952 14340
rect 2004 14328 2010 14340
rect 3068 14328 3096 14359
rect 4062 14356 4068 14368
rect 4120 14396 4126 14408
rect 4632 14405 4660 14436
rect 7190 14424 7196 14476
rect 7248 14464 7254 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 7248 14436 7573 14464
rect 7248 14424 7254 14436
rect 7561 14433 7573 14436
rect 7607 14464 7619 14467
rect 8018 14464 8024 14476
rect 7607 14436 8024 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 13262 14464 13268 14476
rect 13223 14436 13268 14464
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4120 14368 4537 14396
rect 4120 14356 4126 14368
rect 4525 14365 4537 14368
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14396 4675 14399
rect 4982 14396 4988 14408
rect 4663 14368 4988 14396
rect 4663 14365 4675 14368
rect 4617 14359 4675 14365
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 6086 14356 6092 14408
rect 6144 14396 6150 14408
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 6144 14368 6193 14396
rect 6144 14356 6150 14368
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 7653 14399 7711 14405
rect 7653 14396 7665 14399
rect 7524 14368 7665 14396
rect 7524 14356 7530 14368
rect 7653 14365 7665 14368
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14396 7895 14399
rect 8570 14396 8576 14408
rect 7883 14368 8576 14396
rect 7883 14365 7895 14368
rect 7837 14359 7895 14365
rect 7006 14328 7012 14340
rect 2004 14300 3096 14328
rect 6919 14300 7012 14328
rect 2004 14288 2010 14300
rect 7006 14288 7012 14300
rect 7064 14328 7070 14340
rect 7852 14328 7880 14359
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 7064 14300 7880 14328
rect 7064 14288 7070 14300
rect 10226 14288 10232 14340
rect 10284 14328 10290 14340
rect 10428 14328 10456 14356
rect 10781 14331 10839 14337
rect 10781 14328 10793 14331
rect 10284 14300 10793 14328
rect 10284 14288 10290 14300
rect 10781 14297 10793 14300
rect 10827 14297 10839 14331
rect 10781 14291 10839 14297
rect 1673 14263 1731 14269
rect 1673 14229 1685 14263
rect 1719 14260 1731 14263
rect 1762 14260 1768 14272
rect 1719 14232 1768 14260
rect 1719 14229 1731 14232
rect 1673 14223 1731 14229
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 2222 14260 2228 14272
rect 2183 14232 2228 14260
rect 2222 14220 2228 14232
rect 2280 14220 2286 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5629 14263 5687 14269
rect 5629 14260 5641 14263
rect 5592 14232 5641 14260
rect 5592 14220 5598 14232
rect 5629 14229 5641 14232
rect 5675 14229 5687 14263
rect 5629 14223 5687 14229
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7282 14260 7288 14272
rect 7239 14232 7288 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 8110 14260 8116 14272
rect 7800 14232 8116 14260
rect 7800 14220 7806 14232
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10413 14263 10471 14269
rect 10413 14260 10425 14263
rect 10100 14232 10425 14260
rect 10100 14220 10106 14232
rect 10413 14229 10425 14232
rect 10459 14229 10471 14263
rect 10413 14223 10471 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14056 1731 14059
rect 1946 14056 1952 14068
rect 1719 14028 1952 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14056 2191 14059
rect 2498 14056 2504 14068
rect 2179 14028 2504 14056
rect 2179 14025 2191 14028
rect 2133 14019 2191 14025
rect 2498 14016 2504 14028
rect 2556 14016 2562 14068
rect 3234 14056 3240 14068
rect 3195 14028 3240 14056
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 4706 14056 4712 14068
rect 3651 14028 4712 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 5040 14028 5089 14056
rect 5040 14016 5046 14028
rect 5077 14025 5089 14028
rect 5123 14025 5135 14059
rect 5077 14019 5135 14025
rect 5721 14059 5779 14065
rect 5721 14025 5733 14059
rect 5767 14056 5779 14059
rect 5810 14056 5816 14068
rect 5767 14028 5816 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 6086 14056 6092 14068
rect 6047 14028 6092 14056
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 8018 14056 8024 14068
rect 6687 14028 8024 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 3418 13948 3424 14000
rect 3476 13988 3482 14000
rect 3476 13960 3740 13988
rect 3476 13948 3482 13960
rect 2222 13880 2228 13932
rect 2280 13920 2286 13932
rect 3712 13929 3740 13960
rect 2685 13923 2743 13929
rect 2685 13920 2697 13923
rect 2280 13892 2697 13920
rect 2280 13880 2286 13892
rect 2685 13889 2697 13892
rect 2731 13920 2743 13923
rect 3697 13923 3755 13929
rect 2731 13892 3556 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13852 2099 13855
rect 2590 13852 2596 13864
rect 2087 13824 2596 13852
rect 2087 13821 2099 13824
rect 2041 13815 2099 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3418 13852 3424 13864
rect 2700 13824 3424 13852
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 2501 13719 2559 13725
rect 2501 13716 2513 13719
rect 2464 13688 2513 13716
rect 2464 13676 2470 13688
rect 2501 13685 2513 13688
rect 2547 13685 2559 13719
rect 2501 13679 2559 13685
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 2700 13716 2728 13824
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 3528 13796 3556 13892
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 6914 13920 6920 13932
rect 6875 13892 6920 13920
rect 3697 13883 3755 13889
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 3510 13744 3516 13796
rect 3568 13784 3574 13796
rect 3942 13787 4000 13793
rect 3942 13784 3954 13787
rect 3568 13756 3954 13784
rect 3568 13744 3574 13756
rect 3942 13753 3954 13756
rect 3988 13753 4000 13787
rect 3942 13747 4000 13753
rect 6086 13744 6092 13796
rect 6144 13784 6150 13796
rect 6932 13784 6960 13880
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 7173 13855 7231 13861
rect 7173 13852 7185 13855
rect 7064 13824 7185 13852
rect 7064 13812 7070 13824
rect 7173 13821 7185 13824
rect 7219 13821 7231 13855
rect 7173 13815 7231 13821
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8628 13824 8861 13852
rect 8628 13812 8634 13824
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 8849 13815 8907 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 6144 13756 6960 13784
rect 6144 13744 6150 13756
rect 8294 13716 8300 13728
rect 2648 13688 2728 13716
rect 8255 13688 8300 13716
rect 2648 13676 2654 13688
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 2314 13512 2320 13524
rect 2271 13484 2320 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2314 13472 2320 13484
rect 2372 13472 2378 13524
rect 2774 13512 2780 13524
rect 2424 13484 2780 13512
rect 2424 13249 2452 13484
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 4062 13512 4068 13524
rect 4023 13484 4068 13512
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 6144 13484 6653 13512
rect 6144 13472 6150 13484
rect 6472 13456 6500 13484
rect 6641 13481 6653 13484
rect 6687 13481 6699 13515
rect 6641 13475 6699 13481
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8110 13512 8116 13524
rect 7892 13484 8116 13512
rect 7892 13472 7898 13484
rect 8110 13472 8116 13484
rect 8168 13512 8174 13524
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 8168 13484 8217 13512
rect 8168 13472 8174 13484
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 8205 13475 8263 13481
rect 4522 13444 4528 13456
rect 4483 13416 4528 13444
rect 4522 13404 4528 13416
rect 4580 13404 4586 13456
rect 6454 13404 6460 13456
rect 6512 13404 6518 13456
rect 7466 13404 7472 13456
rect 7524 13444 7530 13456
rect 11968 13447 12026 13453
rect 7524 13416 7604 13444
rect 7524 13404 7530 13416
rect 2590 13336 2596 13388
rect 2648 13376 2654 13388
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2648 13348 2789 13376
rect 2648 13336 2654 13348
rect 2777 13345 2789 13348
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 2866 13336 2872 13388
rect 2924 13376 2930 13388
rect 3605 13379 3663 13385
rect 3605 13376 3617 13379
rect 2924 13348 3617 13376
rect 2924 13336 2930 13348
rect 3605 13345 3617 13348
rect 3651 13345 3663 13379
rect 3605 13339 3663 13345
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4706 13376 4712 13388
rect 4479 13348 4712 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 7190 13376 7196 13388
rect 7151 13348 7196 13376
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 7576 13376 7604 13416
rect 11968 13413 11980 13447
rect 12014 13444 12026 13447
rect 12066 13444 12072 13456
rect 12014 13416 12072 13444
rect 12014 13413 12026 13416
rect 11968 13407 12026 13413
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 7834 13376 7840 13388
rect 7576 13348 7840 13376
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 10042 13336 10048 13388
rect 10100 13376 10106 13388
rect 10321 13379 10379 13385
rect 10321 13376 10333 13379
rect 10100 13348 10333 13376
rect 10100 13336 10106 13348
rect 10321 13345 10333 13348
rect 10367 13345 10379 13379
rect 10321 13339 10379 13345
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 3099 13280 4629 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 1857 13243 1915 13249
rect 1857 13209 1869 13243
rect 1903 13240 1915 13243
rect 2409 13243 2467 13249
rect 2409 13240 2421 13243
rect 1903 13212 2421 13240
rect 1903 13209 1915 13212
rect 1857 13203 1915 13209
rect 2409 13209 2421 13212
rect 2455 13209 2467 13243
rect 2409 13203 2467 13209
rect 3528 13184 3556 13280
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 7282 13308 7288 13320
rect 7243 13280 7288 13308
rect 4617 13271 4675 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 8754 13308 8760 13320
rect 7524 13280 8760 13308
rect 7524 13268 7530 13280
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 10008 13280 10425 13308
rect 10008 13268 10014 13280
rect 10413 13277 10425 13280
rect 10459 13277 10471 13311
rect 10594 13308 10600 13320
rect 10555 13280 10600 13308
rect 10413 13271 10471 13277
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11701 13311 11759 13317
rect 11701 13308 11713 13311
rect 11388 13280 11713 13308
rect 11388 13268 11394 13280
rect 11701 13277 11713 13280
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 3605 13243 3663 13249
rect 3605 13209 3617 13243
rect 3651 13240 3663 13243
rect 3651 13212 5304 13240
rect 3651 13209 3663 13212
rect 3605 13203 3663 13209
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 3697 13175 3755 13181
rect 3697 13172 3709 13175
rect 3568 13144 3709 13172
rect 3568 13132 3574 13144
rect 3697 13141 3709 13144
rect 3743 13141 3755 13175
rect 5166 13172 5172 13184
rect 5127 13144 5172 13172
rect 3697 13135 3755 13141
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5276 13172 5304 13212
rect 5810 13200 5816 13252
rect 5868 13240 5874 13252
rect 6825 13243 6883 13249
rect 6825 13240 6837 13243
rect 5868 13212 6837 13240
rect 5868 13200 5874 13212
rect 6825 13209 6837 13212
rect 6871 13209 6883 13243
rect 7834 13240 7840 13252
rect 7795 13212 7840 13240
rect 6825 13203 6883 13209
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 9306 13172 9312 13184
rect 5276 13144 9312 13172
rect 9306 13132 9312 13144
rect 9364 13172 9370 13184
rect 9766 13172 9772 13184
rect 9364 13144 9772 13172
rect 9364 13132 9370 13144
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13172 10011 13175
rect 10502 13172 10508 13184
rect 9999 13144 10508 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 10962 13172 10968 13184
rect 10923 13144 10968 13172
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 13078 13172 13084 13184
rect 13039 13144 13084 13172
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12968 2191 12971
rect 2866 12968 2872 12980
rect 2179 12940 2872 12968
rect 2179 12937 2191 12940
rect 2133 12931 2191 12937
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 4249 12971 4307 12977
rect 4249 12937 4261 12971
rect 4295 12968 4307 12971
rect 4522 12968 4528 12980
rect 4295 12940 4528 12968
rect 4295 12937 4307 12940
rect 4249 12931 4307 12937
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 7377 12971 7435 12977
rect 7377 12968 7389 12971
rect 7340 12940 7389 12968
rect 7340 12928 7346 12940
rect 7377 12937 7389 12940
rect 7423 12937 7435 12971
rect 7377 12931 7435 12937
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10505 12971 10563 12977
rect 10505 12968 10517 12971
rect 9732 12940 10517 12968
rect 9732 12928 9738 12940
rect 10505 12937 10517 12940
rect 10551 12937 10563 12971
rect 10505 12931 10563 12937
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 11514 12968 11520 12980
rect 10652 12940 11520 12968
rect 10652 12928 10658 12940
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 7101 12903 7159 12909
rect 7101 12869 7113 12903
rect 7147 12900 7159 12903
rect 7466 12900 7472 12912
rect 7147 12872 7472 12900
rect 7147 12869 7159 12872
rect 7101 12863 7159 12869
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 10413 12903 10471 12909
rect 10413 12869 10425 12903
rect 10459 12900 10471 12903
rect 10459 12872 11192 12900
rect 10459 12869 10471 12872
rect 10413 12863 10471 12869
rect 11164 12844 11192 12872
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 11388 12872 12633 12900
rect 11388 12860 11394 12872
rect 12621 12869 12633 12872
rect 12667 12869 12679 12903
rect 12621 12863 12679 12869
rect 2222 12832 2228 12844
rect 2183 12804 2228 12832
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5224 12804 5549 12832
rect 5224 12792 5230 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7892 12804 7941 12832
rect 7892 12792 7898 12804
rect 7929 12801 7941 12804
rect 7975 12832 7987 12835
rect 10962 12832 10968 12844
rect 7975 12804 8156 12832
rect 10923 12804 10968 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12764 5506 12776
rect 5997 12767 6055 12773
rect 5997 12764 6009 12767
rect 5500 12736 6009 12764
rect 5500 12724 5506 12736
rect 5997 12733 6009 12736
rect 6043 12733 6055 12767
rect 5997 12727 6055 12733
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12733 8079 12767
rect 8128 12764 8156 12804
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 8294 12773 8300 12776
rect 8288 12764 8300 12773
rect 8128 12736 8300 12764
rect 8021 12727 8079 12733
rect 8288 12727 8300 12736
rect 2498 12705 2504 12708
rect 1765 12699 1823 12705
rect 1765 12665 1777 12699
rect 1811 12696 1823 12699
rect 2470 12699 2504 12705
rect 2470 12696 2482 12699
rect 1811 12668 2482 12696
rect 1811 12665 1823 12668
rect 1765 12659 1823 12665
rect 2470 12665 2482 12668
rect 2556 12696 2562 12708
rect 2556 12668 2618 12696
rect 2470 12659 2504 12665
rect 2498 12656 2504 12659
rect 2556 12656 2562 12668
rect 4522 12656 4528 12708
rect 4580 12696 4586 12708
rect 5074 12696 5080 12708
rect 4580 12668 5080 12696
rect 4580 12656 4586 12668
rect 5074 12656 5080 12668
rect 5132 12656 5138 12708
rect 5353 12699 5411 12705
rect 5353 12665 5365 12699
rect 5399 12696 5411 12699
rect 5534 12696 5540 12708
rect 5399 12668 5540 12696
rect 5399 12665 5411 12668
rect 5353 12659 5411 12665
rect 5534 12656 5540 12668
rect 5592 12696 5598 12708
rect 6365 12699 6423 12705
rect 6365 12696 6377 12699
rect 5592 12668 6377 12696
rect 5592 12656 5598 12668
rect 6365 12665 6377 12668
rect 6411 12665 6423 12699
rect 6365 12659 6423 12665
rect 6454 12656 6460 12708
rect 6512 12656 6518 12708
rect 8036 12696 8064 12727
rect 8294 12724 8300 12727
rect 8352 12724 8358 12776
rect 8110 12696 8116 12708
rect 8036 12668 8116 12696
rect 8110 12656 8116 12668
rect 8168 12696 8174 12708
rect 8386 12696 8392 12708
rect 8168 12668 8392 12696
rect 8168 12656 8174 12668
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 9490 12696 9496 12708
rect 8680 12668 9496 12696
rect 2958 12588 2964 12640
rect 3016 12628 3022 12640
rect 3510 12628 3516 12640
rect 3016 12600 3516 12628
rect 3016 12588 3022 12600
rect 3510 12588 3516 12600
rect 3568 12628 3574 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3568 12600 3617 12628
rect 3568 12588 3574 12600
rect 3605 12597 3617 12600
rect 3651 12597 3663 12631
rect 3605 12591 3663 12597
rect 4617 12631 4675 12637
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 4706 12628 4712 12640
rect 4663 12600 4712 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5442 12588 5448 12640
rect 5500 12628 5506 12640
rect 6472 12628 6500 12656
rect 8680 12640 8708 12668
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 5500 12600 6500 12628
rect 5500 12588 5506 12600
rect 8662 12588 8668 12640
rect 8720 12588 8726 12640
rect 8754 12588 8760 12640
rect 8812 12628 8818 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8812 12600 9413 12628
rect 8812 12588 8818 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 10042 12628 10048 12640
rect 10003 12600 10048 12628
rect 9401 12591 9459 12597
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 10870 12628 10876 12640
rect 10831 12600 10876 12628
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 11977 12631 12035 12637
rect 11977 12597 11989 12631
rect 12023 12628 12035 12631
rect 12066 12628 12072 12640
rect 12023 12600 12072 12628
rect 12023 12597 12035 12600
rect 11977 12591 12035 12597
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 5166 12384 5172 12436
rect 5224 12424 5230 12436
rect 5626 12424 5632 12436
rect 5224 12396 5632 12424
rect 5224 12384 5230 12396
rect 5626 12384 5632 12396
rect 5684 12424 5690 12436
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 5684 12396 6561 12424
rect 5684 12384 5690 12396
rect 6549 12393 6561 12396
rect 6595 12393 6607 12427
rect 7098 12424 7104 12436
rect 7059 12396 7104 12424
rect 6549 12387 6607 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7248 12396 7481 12424
rect 7248 12384 7254 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 7469 12387 7527 12393
rect 8389 12427 8447 12433
rect 8389 12393 8401 12427
rect 8435 12424 8447 12427
rect 8662 12424 8668 12436
rect 8435 12396 8668 12424
rect 8435 12393 8447 12396
rect 8389 12387 8447 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9950 12424 9956 12436
rect 9911 12396 9956 12424
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 10045 12427 10103 12433
rect 10045 12393 10057 12427
rect 10091 12424 10103 12427
rect 10962 12424 10968 12436
rect 10091 12396 10968 12424
rect 10091 12393 10103 12396
rect 10045 12387 10103 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 13078 12424 13084 12436
rect 12032 12396 13084 12424
rect 12032 12384 12038 12396
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 1670 12356 1676 12368
rect 1631 12328 1676 12356
rect 1670 12316 1676 12328
rect 1728 12316 1734 12368
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 5414 12359 5472 12365
rect 5414 12356 5426 12359
rect 3292 12328 5426 12356
rect 3292 12316 3298 12328
rect 5414 12325 5426 12328
rect 5460 12356 5472 12359
rect 5718 12356 5724 12368
rect 5460 12328 5724 12356
rect 5460 12325 5472 12328
rect 5414 12319 5472 12325
rect 5718 12316 5724 12328
rect 5776 12356 5782 12368
rect 6178 12356 6184 12368
rect 5776 12328 6184 12356
rect 5776 12316 5782 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 8110 12316 8116 12368
rect 8168 12356 8174 12368
rect 11422 12356 11428 12368
rect 8168 12328 11428 12356
rect 8168 12316 8174 12328
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 11854 12359 11912 12365
rect 11854 12356 11866 12359
rect 11572 12328 11866 12356
rect 11572 12316 11578 12328
rect 11854 12325 11866 12328
rect 11900 12325 11912 12359
rect 11854 12319 11912 12325
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 10410 12288 10416 12300
rect 7975 12260 8616 12288
rect 10371 12260 10416 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 2958 12220 2964 12232
rect 2915 12192 2964 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 2958 12180 2964 12192
rect 3016 12220 3022 12232
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 3016 12192 4261 12220
rect 3016 12180 3022 12192
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 5166 12220 5172 12232
rect 4249 12183 4307 12189
rect 4908 12192 5172 12220
rect 4908 12161 4936 12192
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 8202 12220 8208 12232
rect 7800 12192 8208 12220
rect 7800 12180 7806 12192
rect 8202 12180 8208 12192
rect 8260 12220 8266 12232
rect 8588 12229 8616 12260
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 8260 12192 8493 12220
rect 8260 12180 8266 12192
rect 8481 12189 8493 12192
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 10042 12220 10048 12232
rect 8619 12192 10048 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10686 12220 10692 12232
rect 10647 12192 10692 12220
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11054 12180 11060 12232
rect 11112 12180 11118 12232
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 11606 12220 11612 12232
rect 11388 12192 11612 12220
rect 11388 12180 11394 12192
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 4893 12155 4951 12161
rect 4893 12121 4905 12155
rect 4939 12121 4951 12155
rect 4893 12115 4951 12121
rect 8021 12155 8079 12161
rect 8021 12121 8033 12155
rect 8067 12152 8079 12155
rect 9950 12152 9956 12164
rect 8067 12124 9956 12152
rect 8067 12121 8079 12124
rect 8021 12115 8079 12121
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 11072 12152 11100 12180
rect 11422 12152 11428 12164
rect 11072 12124 11428 12152
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 2406 12084 2412 12096
rect 2367 12056 2412 12084
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 3234 12084 3240 12096
rect 3195 12056 3240 12084
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 4798 12084 4804 12096
rect 4759 12056 4804 12084
rect 4798 12044 4804 12056
rect 4856 12084 4862 12096
rect 4982 12084 4988 12096
rect 4856 12056 4988 12084
rect 4856 12044 4862 12056
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5442 12084 5448 12096
rect 5224 12056 5448 12084
rect 5224 12044 5230 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 11146 12084 11152 12096
rect 11107 12056 11152 12084
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12084 11575 12087
rect 11790 12084 11796 12096
rect 11563 12056 11796 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 12986 12084 12992 12096
rect 12947 12056 12992 12084
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 2314 11840 2320 11892
rect 2372 11880 2378 11892
rect 2501 11883 2559 11889
rect 2501 11880 2513 11883
rect 2372 11852 2513 11880
rect 2372 11840 2378 11852
rect 2501 11849 2513 11852
rect 2547 11849 2559 11883
rect 5718 11880 5724 11892
rect 5679 11852 5724 11880
rect 2501 11843 2559 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7282 11880 7288 11892
rect 7055 11852 7288 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 10042 11880 10048 11892
rect 10003 11852 10048 11880
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10560 11852 10977 11880
rect 10560 11840 10566 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 12437 11883 12495 11889
rect 12437 11880 12449 11883
rect 11204 11852 12449 11880
rect 11204 11840 11210 11852
rect 12437 11849 12449 11852
rect 12483 11849 12495 11883
rect 12437 11843 12495 11849
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 13354 11880 13360 11892
rect 12676 11852 13360 11880
rect 12676 11840 12682 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 2225 11815 2283 11821
rect 2225 11812 2237 11815
rect 1412 11784 2237 11812
rect 1412 11685 1440 11784
rect 2225 11781 2237 11784
rect 2271 11812 2283 11815
rect 4709 11815 4767 11821
rect 4709 11812 4721 11815
rect 2271 11784 4721 11812
rect 2271 11781 2283 11784
rect 2225 11775 2283 11781
rect 4709 11781 4721 11784
rect 4755 11781 4767 11815
rect 10686 11812 10692 11824
rect 10647 11784 10692 11812
rect 4709 11775 4767 11781
rect 10686 11772 10692 11784
rect 10744 11812 10750 11824
rect 12066 11812 12072 11824
rect 10744 11784 12072 11812
rect 10744 11772 10750 11784
rect 12066 11772 12072 11784
rect 12124 11812 12130 11824
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 12124 11784 12173 11812
rect 12124 11772 12130 11784
rect 12161 11781 12173 11784
rect 12207 11812 12219 11815
rect 12207 11784 13032 11812
rect 12207 11781 12219 11784
rect 12161 11775 12219 11781
rect 13004 11756 13032 11784
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 3234 11704 3240 11756
rect 3292 11744 3298 11756
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 3292 11716 3709 11744
rect 3292 11704 3298 11716
rect 3697 11713 3709 11716
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 4798 11704 4804 11756
rect 4856 11744 4862 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4856 11716 5181 11744
rect 4856 11704 4862 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 6687 11716 7665 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7653 11713 7665 11716
rect 7699 11744 7711 11747
rect 7834 11744 7840 11756
rect 7699 11716 7840 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11645 1455 11679
rect 3602 11676 3608 11688
rect 3563 11648 3608 11676
rect 1397 11639 1455 11645
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11676 4675 11679
rect 5276 11676 5304 11707
rect 7834 11704 7840 11716
rect 7892 11744 7898 11756
rect 8018 11744 8024 11756
rect 7892 11716 8024 11744
rect 7892 11704 7898 11716
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 8444 11716 8677 11744
rect 8444 11704 8450 11716
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 11514 11704 11520 11756
rect 11572 11744 11578 11756
rect 11609 11747 11667 11753
rect 11609 11744 11621 11747
rect 11572 11716 11621 11744
rect 11572 11704 11578 11716
rect 11609 11713 11621 11716
rect 11655 11713 11667 11747
rect 11609 11707 11667 11713
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 13044 11716 13093 11744
rect 13044 11704 13050 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 5350 11676 5356 11688
rect 4663 11648 5356 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7377 11679 7435 11685
rect 7377 11676 7389 11679
rect 7156 11648 7389 11676
rect 7156 11636 7162 11648
rect 7377 11645 7389 11648
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 8921 11679 8979 11685
rect 8921 11676 8933 11679
rect 8812 11648 8933 11676
rect 8812 11636 8818 11648
rect 8921 11645 8933 11648
rect 8967 11645 8979 11679
rect 8921 11639 8979 11645
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11333 11679 11391 11685
rect 11333 11676 11345 11679
rect 11112 11648 11345 11676
rect 11112 11636 11118 11648
rect 11333 11645 11345 11648
rect 11379 11676 11391 11679
rect 11790 11676 11796 11688
rect 11379 11648 11796 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 3053 11611 3111 11617
rect 3053 11577 3065 11611
rect 3099 11608 3111 11611
rect 4249 11611 4307 11617
rect 3099 11580 3556 11608
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 3528 11552 3556 11580
rect 4249 11577 4261 11611
rect 4295 11608 4307 11611
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4295 11580 5089 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 5077 11577 5089 11580
rect 5123 11608 5135 11611
rect 5442 11608 5448 11620
rect 5123 11580 5448 11608
rect 5123 11577 5135 11580
rect 5077 11571 5135 11577
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 11606 11568 11612 11620
rect 11664 11568 11670 11620
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 13354 11608 13360 11620
rect 12584 11580 13360 11608
rect 12584 11568 12590 11580
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 3142 11540 3148 11552
rect 3103 11512 3148 11540
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7469 11543 7527 11549
rect 7469 11540 7481 11543
rect 7156 11512 7481 11540
rect 7156 11500 7162 11512
rect 7469 11509 7481 11512
rect 7515 11509 7527 11543
rect 7469 11503 7527 11509
rect 8113 11543 8171 11549
rect 8113 11509 8125 11543
rect 8159 11540 8171 11543
rect 8202 11540 8208 11552
rect 8159 11512 8208 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8481 11543 8539 11549
rect 8481 11509 8493 11543
rect 8527 11540 8539 11543
rect 8662 11540 8668 11552
rect 8527 11512 8668 11540
rect 8527 11509 8539 11512
rect 8481 11503 8539 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 9824 11512 11161 11540
rect 9824 11500 9830 11512
rect 11149 11509 11161 11512
rect 11195 11540 11207 11543
rect 11238 11540 11244 11552
rect 11195 11512 11244 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11238 11500 11244 11512
rect 11296 11540 11302 11552
rect 11624 11540 11652 11568
rect 12802 11540 12808 11552
rect 11296 11512 11652 11540
rect 12763 11512 12808 11540
rect 11296 11500 11302 11512
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 12986 11540 12992 11552
rect 12943 11512 12992 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 12986 11500 12992 11512
rect 13044 11540 13050 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13044 11512 13461 11540
rect 13044 11500 13050 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1762 11336 1768 11348
rect 1719 11308 1768 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 3602 11336 3608 11348
rect 3283 11308 3608 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5074 11336 5080 11348
rect 5031 11308 5080 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 5224 11308 5273 11336
rect 5224 11296 5230 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5261 11299 5319 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5902 11336 5908 11348
rect 5863 11308 5908 11336
rect 5902 11296 5908 11308
rect 5960 11296 5966 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 7248 11308 7481 11336
rect 7248 11296 7254 11308
rect 7469 11305 7481 11308
rect 7515 11305 7527 11339
rect 8754 11336 8760 11348
rect 8715 11308 8760 11336
rect 7469 11299 7527 11305
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11336 11115 11339
rect 11514 11336 11520 11348
rect 11103 11308 11520 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12802 11336 12808 11348
rect 12207 11308 12808 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12802 11296 12808 11308
rect 12860 11336 12866 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 12860 11308 13185 11336
rect 12860 11296 12866 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13173 11299 13231 11305
rect 7650 11228 7656 11280
rect 7708 11268 7714 11280
rect 7926 11268 7932 11280
rect 7708 11240 7932 11268
rect 7708 11228 7714 11240
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 8386 11228 8392 11280
rect 8444 11268 8450 11280
rect 9033 11271 9091 11277
rect 9033 11268 9045 11271
rect 8444 11240 9045 11268
rect 8444 11228 8450 11240
rect 9033 11237 9045 11240
rect 9079 11237 9091 11271
rect 9033 11231 9091 11237
rect 9493 11271 9551 11277
rect 9493 11237 9505 11271
rect 9539 11268 9551 11271
rect 10410 11268 10416 11280
rect 9539 11240 10416 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 5810 11200 5816 11212
rect 5771 11172 5816 11200
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 7834 11200 7840 11212
rect 7795 11172 7840 11200
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 9048 11200 9076 11231
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 11238 11228 11244 11280
rect 11296 11268 11302 11280
rect 11609 11271 11667 11277
rect 11609 11268 11621 11271
rect 11296 11240 11621 11268
rect 11296 11228 11302 11240
rect 11609 11237 11621 11240
rect 11655 11237 11667 11271
rect 12618 11268 12624 11280
rect 12579 11240 12624 11268
rect 11609 11231 11667 11237
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9048 11172 9689 11200
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9950 11209 9956 11212
rect 9944 11200 9956 11209
rect 9911 11172 9956 11200
rect 9944 11163 9956 11172
rect 9950 11160 9956 11163
rect 10008 11160 10014 11212
rect 12526 11200 12532 11212
rect 12487 11172 12532 11200
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4890 11132 4896 11144
rect 4663 11104 4896 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5626 11092 5632 11144
rect 5684 11132 5690 11144
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5684 11104 6009 11132
rect 5684 11092 5690 11104
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7926 11132 7932 11144
rect 6779 11104 7932 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8076 11104 8121 11132
rect 8076 11092 8082 11104
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 11572 11104 12572 11132
rect 11572 11092 11578 11104
rect 7098 11064 7104 11076
rect 7059 11036 7104 11064
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 12342 11024 12348 11076
rect 12400 11064 12406 11076
rect 12544 11064 12572 11104
rect 12728 11104 12817 11132
rect 12728 11064 12756 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12986 11064 12992 11076
rect 12400 11036 12480 11064
rect 12544 11036 12756 11064
rect 12820 11036 12992 11064
rect 12400 11024 12406 11036
rect 6178 10956 6184 11008
rect 6236 10996 6242 11008
rect 6730 10996 6736 11008
rect 6236 10968 6736 10996
rect 6236 10956 6242 10968
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 12452 10996 12480 11036
rect 12820 10996 12848 11036
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 12452 10968 12848 10996
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 5626 10792 5632 10804
rect 5587 10764 5632 10792
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 5868 10764 6469 10792
rect 5868 10752 5874 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 6457 10755 6515 10761
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8021 10795 8079 10801
rect 8021 10792 8033 10795
rect 7984 10764 8033 10792
rect 7984 10752 7990 10764
rect 8021 10761 8033 10764
rect 8067 10761 8079 10795
rect 8021 10755 8079 10761
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 9950 10792 9956 10804
rect 9815 10764 9956 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10468 10764 10609 10792
rect 10468 10752 10474 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11572 10764 11805 10792
rect 11572 10752 11578 10764
rect 11793 10761 11805 10764
rect 11839 10792 11851 10795
rect 12066 10792 12072 10804
rect 11839 10764 12072 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12710 10792 12716 10804
rect 12299 10764 12716 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 2590 10684 2596 10736
rect 2648 10724 2654 10736
rect 2961 10727 3019 10733
rect 2961 10724 2973 10727
rect 2648 10696 2973 10724
rect 2648 10684 2654 10696
rect 2961 10693 2973 10696
rect 3007 10693 3019 10727
rect 2961 10687 3019 10693
rect 4433 10727 4491 10733
rect 4433 10693 4445 10727
rect 4479 10724 4491 10727
rect 4479 10696 5212 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2866 10656 2872 10668
rect 2779 10628 2872 10656
rect 2866 10616 2872 10628
rect 2924 10656 2930 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 2924 10628 3617 10656
rect 2924 10616 2930 10628
rect 3605 10625 3617 10628
rect 3651 10656 3663 10659
rect 4062 10656 4068 10668
rect 3651 10628 4068 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1762 10588 1768 10600
rect 1443 10560 1768 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 3973 10591 4031 10597
rect 2547 10560 3188 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3160 10452 3188 10560
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4798 10588 4804 10600
rect 4019 10560 4804 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4798 10548 4804 10560
rect 4856 10588 4862 10600
rect 5092 10588 5120 10619
rect 4856 10560 5120 10588
rect 4856 10548 4862 10560
rect 3326 10520 3332 10532
rect 3239 10492 3332 10520
rect 3326 10480 3332 10492
rect 3384 10520 3390 10532
rect 4985 10523 5043 10529
rect 3384 10492 4568 10520
rect 3384 10480 3390 10492
rect 3418 10452 3424 10464
rect 3160 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4540 10461 4568 10492
rect 4985 10489 4997 10523
rect 5031 10520 5043 10523
rect 5184 10520 5212 10696
rect 5718 10684 5724 10736
rect 5776 10724 5782 10736
rect 6089 10727 6147 10733
rect 6089 10724 6101 10727
rect 5776 10696 6101 10724
rect 5776 10684 5782 10696
rect 6089 10693 6101 10696
rect 6135 10724 6147 10727
rect 6730 10724 6736 10736
rect 6135 10696 6736 10724
rect 6135 10693 6147 10696
rect 6089 10687 6147 10693
rect 6730 10684 6736 10696
rect 6788 10684 6794 10736
rect 8570 10656 8576 10668
rect 8531 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10656 8634 10668
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8628 10628 9045 10656
rect 8628 10616 8634 10628
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 10183 10628 11253 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 11241 10625 11253 10628
rect 11287 10656 11299 10659
rect 11532 10656 11560 10752
rect 11287 10628 11560 10656
rect 12437 10659 12495 10665
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12526 10656 12532 10668
rect 12483 10628 12532 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12526 10616 12532 10628
rect 12584 10656 12590 10668
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12584 10628 12909 10656
rect 12584 10616 12590 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10588 7987 10591
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 7975 10560 8401 10588
rect 7975 10557 7987 10560
rect 7929 10551 7987 10557
rect 8389 10557 8401 10560
rect 8435 10588 8447 10591
rect 9398 10588 9404 10600
rect 8435 10560 9404 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 6178 10520 6184 10532
rect 5031 10492 6184 10520
rect 5031 10489 5043 10492
rect 4985 10483 5043 10489
rect 6178 10480 6184 10492
rect 6236 10480 6242 10532
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 11057 10523 11115 10529
rect 11057 10520 11069 10523
rect 10560 10492 11069 10520
rect 10560 10480 10566 10492
rect 11057 10489 11069 10492
rect 11103 10489 11115 10523
rect 11057 10483 11115 10489
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10421 4583 10455
rect 4890 10452 4896 10464
rect 4851 10424 4896 10452
rect 4525 10415 4583 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7561 10455 7619 10461
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 8110 10452 8116 10464
rect 7607 10424 8116 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 8110 10412 8116 10424
rect 8168 10452 8174 10464
rect 8481 10455 8539 10461
rect 8481 10452 8493 10455
rect 8168 10424 8493 10452
rect 8168 10412 8174 10424
rect 8481 10421 8493 10424
rect 8527 10452 8539 10455
rect 9398 10452 9404 10464
rect 8527 10424 9404 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 10410 10452 10416 10464
rect 9916 10424 10416 10452
rect 9916 10412 9922 10424
rect 10410 10412 10416 10424
rect 10468 10452 10474 10464
rect 10965 10455 11023 10461
rect 10965 10452 10977 10455
rect 10468 10424 10977 10452
rect 10468 10412 10474 10424
rect 10965 10421 10977 10424
rect 11011 10421 11023 10455
rect 10965 10415 11023 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 3326 10248 3332 10260
rect 3287 10220 3332 10248
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 3476 10220 4445 10248
rect 3476 10208 3482 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4433 10211 4491 10217
rect 4801 10251 4859 10257
rect 4801 10217 4813 10251
rect 4847 10248 4859 10251
rect 5166 10248 5172 10260
rect 4847 10220 5172 10248
rect 4847 10217 4859 10220
rect 4801 10211 4859 10217
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 5902 10248 5908 10260
rect 5583 10220 5908 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6457 10251 6515 10257
rect 6457 10248 6469 10251
rect 6043 10220 6469 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6457 10217 6469 10220
rect 6503 10248 6515 10251
rect 6822 10248 6828 10260
rect 6503 10220 6828 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7834 10208 7840 10260
rect 7892 10248 7898 10260
rect 8021 10251 8079 10257
rect 8021 10248 8033 10251
rect 7892 10220 8033 10248
rect 7892 10208 7898 10220
rect 8021 10217 8033 10220
rect 8067 10248 8079 10251
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 8067 10220 9045 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 9033 10217 9045 10220
rect 9079 10217 9091 10251
rect 9033 10211 9091 10217
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9824 10220 9873 10248
rect 9824 10208 9830 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 11517 10251 11575 10257
rect 11517 10217 11529 10251
rect 11563 10248 11575 10251
rect 12342 10248 12348 10260
rect 11563 10220 12348 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 6549 10183 6607 10189
rect 6549 10180 6561 10183
rect 6236 10152 6561 10180
rect 6236 10140 6242 10152
rect 6549 10149 6561 10152
rect 6595 10149 6607 10183
rect 11977 10183 12035 10189
rect 11977 10180 11989 10183
rect 6549 10143 6607 10149
rect 11532 10152 11989 10180
rect 11532 10124 11560 10152
rect 11977 10149 11989 10152
rect 12023 10180 12035 10183
rect 13078 10180 13084 10192
rect 12023 10152 13084 10180
rect 12023 10149 12035 10152
rect 11977 10143 12035 10149
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 1670 10072 1676 10124
rect 1728 10112 1734 10124
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 1728 10084 2697 10112
rect 1728 10072 1734 10084
rect 2685 10081 2697 10084
rect 2731 10081 2743 10115
rect 2685 10075 2743 10081
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10112 7803 10115
rect 8018 10112 8024 10124
rect 7791 10084 8024 10112
rect 7791 10081 7803 10084
rect 7745 10075 7803 10081
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8386 10112 8392 10124
rect 8347 10084 8392 10112
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 11514 10072 11520 10124
rect 11572 10072 11578 10124
rect 11885 10115 11943 10121
rect 11885 10081 11897 10115
rect 11931 10112 11943 10115
rect 12342 10112 12348 10124
rect 11931 10084 12348 10112
rect 11931 10081 11943 10084
rect 11885 10075 11943 10081
rect 12342 10072 12348 10084
rect 12400 10112 12406 10124
rect 12434 10112 12440 10124
rect 12400 10084 12440 10112
rect 12400 10072 12406 10084
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 2038 10004 2044 10056
rect 2096 10044 2102 10056
rect 2777 10047 2835 10053
rect 2777 10044 2789 10047
rect 2096 10016 2789 10044
rect 2096 10004 2102 10016
rect 2777 10013 2789 10016
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 2866 10004 2872 10056
rect 2924 10044 2930 10056
rect 2924 10016 2969 10044
rect 2924 10004 2930 10016
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4212 10016 4905 10044
rect 4212 10004 4218 10016
rect 4893 10013 4905 10016
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 6730 10044 6736 10056
rect 6691 10016 6736 10044
rect 4985 10007 5043 10013
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 2884 9976 2912 10004
rect 2464 9948 2912 9976
rect 2464 9936 2470 9948
rect 4798 9936 4804 9988
rect 4856 9976 4862 9988
rect 5000 9976 5028 10007
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 8478 10044 8484 10056
rect 8439 10016 8484 10044
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 8628 10016 8673 10044
rect 8628 10004 8634 10016
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12124 10016 12169 10044
rect 12124 10004 12130 10016
rect 4856 9948 5028 9976
rect 4856 9936 4862 9948
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5868 9948 6101 9976
rect 5868 9936 5874 9948
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 7377 9979 7435 9985
rect 7377 9945 7389 9979
rect 7423 9976 7435 9979
rect 7834 9976 7840 9988
rect 7423 9948 7840 9976
rect 7423 9945 7435 9948
rect 7377 9939 7435 9945
rect 7834 9936 7840 9948
rect 7892 9936 7898 9988
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 1581 9911 1639 9917
rect 1581 9908 1593 9911
rect 1452 9880 1593 9908
rect 1452 9868 1458 9880
rect 1581 9877 1593 9880
rect 1627 9877 1639 9911
rect 1581 9871 1639 9877
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2130 9908 2136 9920
rect 2087 9880 2136 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 2314 9908 2320 9920
rect 2275 9880 2320 9908
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 10597 9911 10655 9917
rect 10597 9908 10609 9911
rect 10560 9880 10609 9908
rect 10560 9868 10566 9880
rect 10597 9877 10609 9880
rect 10643 9877 10655 9911
rect 10597 9871 10655 9877
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 1670 9704 1676 9716
rect 1631 9676 1676 9704
rect 1670 9664 1676 9676
rect 1728 9664 1734 9716
rect 2038 9704 2044 9716
rect 1999 9676 2044 9704
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 6178 9704 6184 9716
rect 6139 9676 6184 9704
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8665 9707 8723 9713
rect 8665 9704 8677 9707
rect 8444 9676 8677 9704
rect 8444 9664 8450 9676
rect 8665 9673 8677 9676
rect 8711 9704 8723 9707
rect 11241 9707 11299 9713
rect 8711 9676 8892 9704
rect 8711 9673 8723 9676
rect 8665 9667 8723 9673
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4249 9639 4307 9645
rect 4249 9636 4261 9639
rect 4120 9608 4261 9636
rect 4120 9596 4126 9608
rect 4249 9605 4261 9608
rect 4295 9605 4307 9639
rect 4249 9599 4307 9605
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5353 9639 5411 9645
rect 5353 9636 5365 9639
rect 5132 9608 5365 9636
rect 5132 9596 5138 9608
rect 5353 9605 5365 9608
rect 5399 9605 5411 9639
rect 6454 9636 6460 9648
rect 6415 9608 6460 9636
rect 5353 9599 5411 9605
rect 6454 9596 6460 9608
rect 6512 9596 6518 9648
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 7101 9639 7159 9645
rect 7101 9636 7113 9639
rect 6972 9608 7113 9636
rect 6972 9596 6978 9608
rect 7101 9605 7113 9608
rect 7147 9605 7159 9639
rect 7101 9599 7159 9605
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2188 9540 2881 9568
rect 2188 9528 2194 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 2884 9500 2912 9531
rect 3418 9500 3424 9512
rect 2884 9472 3424 9500
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9500 4951 9503
rect 5166 9500 5172 9512
rect 4939 9472 5172 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5316 9472 5549 9500
rect 5316 9460 5322 9472
rect 5537 9469 5549 9472
rect 5583 9500 5595 9503
rect 6472 9500 6500 9596
rect 6638 9500 6644 9512
rect 5583 9472 6500 9500
rect 6599 9472 6644 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 7116 9500 7144 9599
rect 7834 9568 7840 9580
rect 7795 9540 7840 9568
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8864 9577 8892 9676
rect 11241 9673 11253 9707
rect 11287 9704 11299 9707
rect 12066 9704 12072 9716
rect 11287 9676 12072 9704
rect 11287 9673 11299 9676
rect 11241 9667 11299 9673
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 11609 9639 11667 9645
rect 11609 9605 11621 9639
rect 11655 9636 11667 9639
rect 12342 9636 12348 9648
rect 11655 9608 12348 9636
rect 11655 9605 11667 9608
rect 11609 9599 11667 9605
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 7374 9500 7380 9512
rect 7116 9472 7380 9500
rect 7374 9460 7380 9472
rect 7432 9500 7438 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7432 9472 7757 9500
rect 7432 9460 7438 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 8570 9460 8576 9512
rect 8628 9500 8634 9512
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 8628 9472 9321 9500
rect 8628 9460 8634 9472
rect 9309 9469 9321 9472
rect 9355 9469 9367 9503
rect 10042 9500 10048 9512
rect 9955 9472 10048 9500
rect 9309 9463 9367 9469
rect 10042 9460 10048 9472
rect 10100 9500 10106 9512
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 10100 9472 10333 9500
rect 10100 9460 10106 9472
rect 10321 9469 10333 9472
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 3114 9435 3172 9441
rect 3114 9432 3126 9435
rect 2792 9404 3126 9432
rect 2792 9376 2820 9404
rect 3114 9401 3126 9404
rect 3160 9401 3172 9435
rect 3114 9395 3172 9401
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7653 9435 7711 9441
rect 7653 9432 7665 9435
rect 7064 9404 7665 9432
rect 7064 9392 7070 9404
rect 7653 9401 7665 9404
rect 7699 9401 7711 9435
rect 7653 9395 7711 9401
rect 8389 9435 8447 9441
rect 8389 9401 8401 9435
rect 8435 9432 8447 9435
rect 8478 9432 8484 9444
rect 8435 9404 8484 9432
rect 8435 9401 8447 9404
rect 8389 9395 8447 9401
rect 8478 9392 8484 9404
rect 8536 9432 8542 9444
rect 9398 9432 9404 9444
rect 8536 9404 9404 9432
rect 8536 9392 8542 9404
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 1820 9336 2329 9364
rect 1820 9324 1826 9336
rect 2317 9333 2329 9336
rect 2363 9364 2375 9367
rect 2406 9364 2412 9376
rect 2363 9336 2412 9364
rect 2363 9333 2375 9336
rect 2317 9327 2375 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2832 9336 2877 9364
rect 2832 9324 2838 9336
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 4212 9336 5181 9364
rect 4212 9324 4218 9336
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 5169 9327 5227 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 9858 9364 9864 9376
rect 9819 9336 9864 9364
rect 9858 9324 9864 9336
rect 9916 9364 9922 9376
rect 10962 9364 10968 9376
rect 9916 9336 10968 9364
rect 9916 9324 9922 9336
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11572 9336 11897 9364
rect 11572 9324 11578 9336
rect 11885 9333 11897 9336
rect 11931 9364 11943 9367
rect 12066 9364 12072 9376
rect 11931 9336 12072 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2556 9132 2881 9160
rect 2556 9120 2562 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 2869 9123 2927 9129
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 4341 9163 4399 9169
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 4890 9160 4896 9172
rect 4387 9132 4896 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5258 9160 5264 9172
rect 5219 9132 5264 9160
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 6730 9160 6736 9172
rect 5592 9132 6736 9160
rect 5592 9120 5598 9132
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 7156 9132 7849 9160
rect 7156 9120 7162 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 7837 9123 7895 9129
rect 2130 9092 2136 9104
rect 1504 9064 2136 9092
rect 1504 9033 1532 9064
rect 2130 9052 2136 9064
rect 2188 9052 2194 9104
rect 5718 9052 5724 9104
rect 5776 9052 5782 9104
rect 7006 9052 7012 9104
rect 7064 9092 7070 9104
rect 7285 9095 7343 9101
rect 7285 9092 7297 9095
rect 7064 9064 7297 9092
rect 7064 9052 7070 9064
rect 7285 9061 7297 9064
rect 7331 9061 7343 9095
rect 7285 9055 7343 9061
rect 1762 9033 1768 9036
rect 1489 9027 1547 9033
rect 1489 8993 1501 9027
rect 1535 8993 1547 9027
rect 1756 9024 1768 9033
rect 1723 8996 1768 9024
rect 1489 8987 1547 8993
rect 1756 8987 1768 8996
rect 1762 8984 1768 8987
rect 1820 8984 1826 9036
rect 3418 8984 3424 9036
rect 3476 9024 3482 9036
rect 5166 9024 5172 9036
rect 3476 8996 5172 9024
rect 3476 8984 3482 8996
rect 5166 8984 5172 8996
rect 5224 9024 5230 9036
rect 5353 9027 5411 9033
rect 5353 9024 5365 9027
rect 5224 8996 5365 9024
rect 5224 8984 5230 8996
rect 5353 8993 5365 8996
rect 5399 8993 5411 9027
rect 5353 8987 5411 8993
rect 5620 9027 5678 9033
rect 5620 8993 5632 9027
rect 5666 9024 5678 9027
rect 5736 9024 5764 9052
rect 6178 9024 6184 9036
rect 5666 8996 6184 9024
rect 5666 8993 5678 8996
rect 5620 8987 5678 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 9024 8263 9027
rect 8754 9024 8760 9036
rect 8251 8996 8760 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 8754 8984 8760 8996
rect 8812 9024 8818 9036
rect 9306 9024 9312 9036
rect 8812 8996 9312 9024
rect 8812 8984 8818 8996
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 4798 8956 4804 8968
rect 2832 8928 4804 8956
rect 2832 8916 2838 8928
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 7340 8928 8309 8956
rect 7340 8916 7346 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8956 8539 8959
rect 8570 8956 8576 8968
rect 8527 8928 8576 8956
rect 8527 8925 8539 8928
rect 8481 8919 8539 8925
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8888 7803 8891
rect 8496 8888 8524 8919
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 7791 8860 8524 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 10226 8820 10232 8832
rect 9539 8792 10232 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2096 8588 2697 8616
rect 2096 8576 2102 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 4948 8588 5641 8616
rect 4948 8576 4954 8588
rect 5629 8585 5641 8588
rect 5675 8585 5687 8619
rect 6178 8616 6184 8628
rect 6139 8588 6184 8616
rect 5629 8579 5687 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 6730 8616 6736 8628
rect 6687 8588 6736 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 8754 8616 8760 8628
rect 8715 8588 8760 8616
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8904 8588 9229 8616
rect 8904 8576 8910 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9217 8579 9275 8585
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 3160 8452 3249 8480
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 3050 8412 3056 8424
rect 2639 8384 3056 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 2225 8347 2283 8353
rect 2225 8313 2237 8347
rect 2271 8344 2283 8347
rect 2774 8344 2780 8356
rect 2271 8316 2780 8344
rect 2271 8313 2283 8316
rect 2225 8307 2283 8313
rect 2774 8304 2780 8316
rect 2832 8344 2838 8356
rect 3160 8344 3188 8452
rect 3237 8449 3249 8452
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 3476 8452 4261 8480
rect 3476 8440 3482 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 6748 8480 6776 8576
rect 9232 8480 9260 8579
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 6748 8452 6960 8480
rect 9232 8452 9873 8480
rect 4249 8443 4307 8449
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 6932 8412 6960 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10226 8480 10232 8492
rect 10091 8452 10232 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 7081 8415 7139 8421
rect 7081 8412 7093 8415
rect 6932 8384 7093 8412
rect 7081 8381 7093 8384
rect 7127 8381 7139 8415
rect 7081 8375 7139 8381
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9490 8412 9496 8424
rect 8812 8384 9496 8412
rect 8812 8372 8818 8384
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9876 8412 9904 8443
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10134 8412 10140 8424
rect 9876 8384 10140 8412
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 2832 8316 3188 8344
rect 4157 8347 4215 8353
rect 2832 8304 2838 8316
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4516 8347 4574 8353
rect 4516 8344 4528 8347
rect 4203 8316 4528 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4516 8313 4528 8316
rect 4562 8344 4574 8347
rect 4798 8344 4804 8356
rect 4562 8316 4804 8344
rect 4562 8313 4574 8316
rect 4516 8307 4574 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 9769 8347 9827 8353
rect 9769 8344 9781 8347
rect 9600 8316 9781 8344
rect 3145 8279 3203 8285
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 3694 8276 3700 8288
rect 3191 8248 3700 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 7834 8276 7840 8288
rect 7248 8248 7840 8276
rect 7248 8236 7254 8248
rect 7834 8236 7840 8248
rect 7892 8276 7898 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7892 8248 8217 8276
rect 7892 8236 7898 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 9398 8276 9404 8288
rect 9359 8248 9404 8276
rect 8205 8239 8263 8245
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 9600 8276 9628 8316
rect 9769 8313 9781 8316
rect 9815 8313 9827 8347
rect 9769 8307 9827 8313
rect 9548 8248 9628 8276
rect 10505 8279 10563 8285
rect 9548 8236 9554 8248
rect 10505 8245 10517 8279
rect 10551 8276 10563 8279
rect 10686 8276 10692 8288
rect 10551 8248 10692 8276
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 1728 8044 2421 8072
rect 1728 8032 1734 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 3694 8032 3700 8084
rect 3752 8072 3758 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3752 8044 4077 8072
rect 3752 8032 3758 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4522 8032 4528 8084
rect 4580 8032 4586 8084
rect 5166 8072 5172 8084
rect 5127 8044 5172 8072
rect 5166 8032 5172 8044
rect 5224 8072 5230 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5224 8044 5457 8072
rect 5224 8032 5230 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6638 8072 6644 8084
rect 6595 8044 6644 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 7009 8075 7067 8081
rect 7009 8041 7021 8075
rect 7055 8072 7067 8075
rect 7282 8072 7288 8084
rect 7055 8044 7288 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 8481 8075 8539 8081
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 8570 8072 8576 8084
rect 8527 8044 8576 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 13081 8075 13139 8081
rect 13081 8072 13093 8075
rect 10827 8044 13093 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 13081 8041 13093 8044
rect 13127 8041 13139 8075
rect 13081 8035 13139 8041
rect 2041 8007 2099 8013
rect 2041 7973 2053 8007
rect 2087 8004 2099 8007
rect 2590 8004 2596 8016
rect 2087 7976 2596 8004
rect 2087 7973 2099 7976
rect 2041 7967 2099 7973
rect 2590 7964 2596 7976
rect 2648 7964 2654 8016
rect 2777 8007 2835 8013
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 2958 8004 2964 8016
rect 2823 7976 2964 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 2958 7964 2964 7976
rect 3016 8004 3022 8016
rect 4540 8004 4568 8032
rect 8294 8004 8300 8016
rect 3016 7976 4568 8004
rect 7024 7976 8300 8004
rect 3016 7964 3022 7976
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1762 7936 1768 7948
rect 1719 7908 1768 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 3326 7936 3332 7948
rect 2915 7908 3332 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4396 7908 4445 7936
rect 4396 7896 4402 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 7024 7936 7052 7976
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 4571 7908 7052 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 2774 7760 2780 7812
rect 2832 7800 2838 7812
rect 2976 7800 3004 7831
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4540 7868 4568 7899
rect 7190 7896 7196 7948
rect 7248 7936 7254 7948
rect 7357 7939 7415 7945
rect 7357 7936 7369 7939
rect 7248 7908 7369 7936
rect 7248 7896 7254 7908
rect 7357 7905 7369 7908
rect 7403 7905 7415 7939
rect 7357 7899 7415 7905
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9916 7908 10057 7936
rect 9916 7896 9922 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 4120 7840 4568 7868
rect 4709 7871 4767 7877
rect 4120 7828 4126 7840
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 4798 7868 4804 7880
rect 4755 7840 4804 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 6822 7868 6828 7880
rect 6227 7840 6828 7868
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 6822 7828 6828 7840
rect 6880 7868 6886 7880
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 6880 7840 7113 7868
rect 6880 7828 6886 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 2832 7772 3004 7800
rect 2832 7760 2838 7772
rect 7116 7732 7144 7831
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9824 7840 10149 7868
rect 9824 7828 9830 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10284 7840 10333 7868
rect 10284 7828 10290 7840
rect 10321 7837 10333 7840
rect 10367 7868 10379 7871
rect 10796 7868 10824 8035
rect 11974 7945 11980 7948
rect 11968 7899 11980 7945
rect 12032 7936 12038 7948
rect 12032 7908 12068 7936
rect 11974 7896 11980 7899
rect 12032 7896 12038 7908
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 10367 7840 10824 7868
rect 11532 7840 11713 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 9401 7803 9459 7809
rect 9401 7800 9413 7803
rect 8352 7772 9413 7800
rect 8352 7760 8358 7772
rect 9401 7769 9413 7772
rect 9447 7800 9459 7803
rect 9490 7800 9496 7812
rect 9447 7772 9496 7800
rect 9447 7769 9459 7772
rect 9401 7763 9459 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 11532 7744 11560 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 7834 7732 7840 7744
rect 7116 7704 7840 7732
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 9125 7735 9183 7741
rect 9125 7701 9137 7735
rect 9171 7732 9183 7735
rect 9306 7732 9312 7744
rect 9171 7704 9312 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 9674 7732 9680 7744
rect 9635 7704 9680 7732
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 11514 7732 11520 7744
rect 11475 7704 11520 7732
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 1857 7531 1915 7537
rect 1857 7528 1869 7531
rect 1452 7500 1869 7528
rect 1452 7488 1458 7500
rect 1857 7497 1869 7500
rect 1903 7497 1915 7531
rect 4062 7528 4068 7540
rect 4023 7500 4068 7528
rect 1857 7491 1915 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 5169 7531 5227 7537
rect 5169 7528 5181 7531
rect 5132 7500 5181 7528
rect 5132 7488 5138 7500
rect 5169 7497 5181 7500
rect 5215 7497 5227 7531
rect 5169 7491 5227 7497
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6822 7528 6828 7540
rect 6687 7500 6828 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7466 7528 7472 7540
rect 7427 7500 7472 7528
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 9582 7528 9588 7540
rect 9048 7500 9588 7528
rect 1765 7463 1823 7469
rect 1765 7429 1777 7463
rect 1811 7460 1823 7463
rect 2498 7460 2504 7472
rect 1811 7432 2504 7460
rect 1811 7429 1823 7432
rect 1765 7423 1823 7429
rect 2314 7392 2320 7404
rect 2275 7364 2320 7392
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2424 7401 2452 7432
rect 2498 7420 2504 7432
rect 2556 7420 2562 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4614 7460 4620 7472
rect 4304 7432 4620 7460
rect 4304 7420 4310 7432
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 7929 7395 7987 7401
rect 2455 7364 2489 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 7975 7364 8953 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8941 7361 8953 7364
rect 8987 7392 8999 7395
rect 9048 7392 9076 7500
rect 9582 7488 9588 7500
rect 9640 7528 9646 7540
rect 11241 7531 11299 7537
rect 11241 7528 11253 7531
rect 9640 7500 11253 7528
rect 9640 7488 9646 7500
rect 11241 7497 11253 7500
rect 11287 7497 11299 7531
rect 11241 7491 11299 7497
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 11974 7528 11980 7540
rect 11931 7500 11980 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 11974 7488 11980 7500
rect 12032 7528 12038 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 12032 7500 12173 7528
rect 12032 7488 12038 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 13262 7528 13268 7540
rect 12483 7500 13268 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 9214 7420 9220 7472
rect 9272 7460 9278 7472
rect 9309 7463 9367 7469
rect 9309 7460 9321 7463
rect 9272 7432 9321 7460
rect 9272 7420 9278 7432
rect 9309 7429 9321 7432
rect 9355 7460 9367 7463
rect 9858 7460 9864 7472
rect 9355 7432 9864 7460
rect 9355 7429 9367 7432
rect 9309 7423 9367 7429
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 8987 7364 9076 7392
rect 12176 7392 12204 7491
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 12952 7432 13308 7460
rect 12952 7420 12958 7432
rect 13280 7404 13308 7432
rect 12802 7392 12808 7404
rect 12176 7364 12808 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 12802 7352 12808 7364
rect 12860 7392 12866 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12860 7364 13001 7392
rect 12860 7352 12866 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13262 7352 13268 7404
rect 13320 7352 13326 7404
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2590 7324 2596 7336
rect 2271 7296 2596 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 3326 7324 3332 7336
rect 3287 7296 3332 7324
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 4798 7324 4804 7336
rect 3835 7296 4804 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 5074 7324 5080 7336
rect 4939 7296 5080 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 7466 7324 7472 7336
rect 6871 7296 7472 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 8202 7324 8208 7336
rect 8163 7296 8208 7324
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7324 8815 7327
rect 9122 7324 9128 7336
rect 8803 7296 9128 7324
rect 8803 7293 8815 7296
rect 8757 7287 8815 7293
rect 9122 7284 9128 7296
rect 9180 7324 9186 7336
rect 9674 7324 9680 7336
rect 9180 7296 9680 7324
rect 9180 7284 9186 7296
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7324 9919 7327
rect 10686 7324 10692 7336
rect 9907 7296 10692 7324
rect 9907 7293 9919 7296
rect 9861 7287 9919 7293
rect 9876 7256 9904 7287
rect 10686 7284 10692 7296
rect 10744 7324 10750 7336
rect 11514 7324 11520 7336
rect 10744 7296 11520 7324
rect 10744 7284 10750 7296
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 8036 7228 9904 7256
rect 10128 7259 10186 7265
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4396 7160 4445 7188
rect 4396 7148 4402 7160
rect 4433 7157 4445 7160
rect 4479 7157 4491 7191
rect 4433 7151 4491 7157
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4580 7160 4721 7188
rect 4580 7148 4586 7160
rect 4709 7157 4721 7160
rect 4755 7188 4767 7191
rect 5166 7188 5172 7200
rect 4755 7160 5172 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7009 7191 7067 7197
rect 7009 7188 7021 7191
rect 6972 7160 7021 7188
rect 6972 7148 6978 7160
rect 7009 7157 7021 7160
rect 7055 7157 7067 7191
rect 7009 7151 7067 7157
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 8036 7197 8064 7228
rect 10128 7225 10140 7259
rect 10174 7256 10186 7259
rect 10226 7256 10232 7268
rect 10174 7228 10232 7256
rect 10174 7225 10186 7228
rect 10128 7219 10186 7225
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 12894 7256 12900 7268
rect 12855 7228 12900 7256
rect 12894 7216 12900 7228
rect 12952 7256 12958 7268
rect 13449 7259 13507 7265
rect 13449 7256 13461 7259
rect 12952 7228 13461 7256
rect 12952 7216 12958 7228
rect 13449 7225 13461 7228
rect 13495 7225 13507 7259
rect 13449 7219 13507 7225
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7892 7160 8033 7188
rect 7892 7148 7898 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8478 7188 8484 7200
rect 8343 7160 8484 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 8665 7191 8723 7197
rect 8665 7157 8677 7191
rect 8711 7188 8723 7191
rect 9214 7188 9220 7200
rect 8711 7160 9220 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9674 7188 9680 7200
rect 9635 7160 9680 7188
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12676 7160 12817 7188
rect 12676 7148 12682 7160
rect 12805 7157 12817 7160
rect 12851 7188 12863 7191
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 12851 7160 13829 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 13817 7151 13875 7157
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 1949 6987 2007 6993
rect 1949 6953 1961 6987
rect 1995 6984 2007 6987
rect 2222 6984 2228 6996
rect 1995 6956 2228 6984
rect 1995 6953 2007 6956
rect 1949 6947 2007 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 2685 6987 2743 6993
rect 2685 6953 2697 6987
rect 2731 6984 2743 6987
rect 2774 6984 2780 6996
rect 2731 6956 2780 6984
rect 2731 6953 2743 6956
rect 2685 6947 2743 6953
rect 2774 6944 2780 6956
rect 2832 6944 2838 6996
rect 7190 6984 7196 6996
rect 7151 6956 7196 6984
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 7561 6987 7619 6993
rect 7561 6953 7573 6987
rect 7607 6984 7619 6987
rect 8202 6984 8208 6996
rect 7607 6956 8208 6984
rect 7607 6953 7619 6956
rect 7561 6947 7619 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 9122 6984 9128 6996
rect 9083 6956 9128 6984
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9861 6987 9919 6993
rect 9861 6984 9873 6987
rect 9272 6956 9873 6984
rect 9272 6944 9278 6956
rect 9861 6953 9873 6956
rect 9907 6953 9919 6987
rect 9861 6947 9919 6953
rect 10229 6987 10287 6993
rect 10229 6953 10241 6987
rect 10275 6984 10287 6987
rect 10502 6984 10508 6996
rect 10275 6956 10508 6984
rect 10275 6953 10287 6956
rect 10229 6947 10287 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 12802 6984 12808 6996
rect 12763 6956 12808 6984
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2130 6848 2136 6860
rect 2087 6820 2136 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2130 6808 2136 6820
rect 2188 6848 2194 6860
rect 2498 6848 2504 6860
rect 2188 6820 2504 6848
rect 2188 6808 2194 6820
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 4706 6808 4712 6860
rect 4764 6848 4770 6860
rect 5166 6848 5172 6860
rect 4764 6820 5172 6848
rect 4764 6808 4770 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 6144 6820 6285 6848
rect 6144 6808 6150 6820
rect 6273 6817 6285 6820
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6848 7987 6851
rect 8386 6848 8392 6860
rect 7975 6820 8392 6848
rect 7975 6817 7987 6820
rect 7929 6811 7987 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 11698 6857 11704 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 10008 6820 10333 6848
rect 10008 6808 10014 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 10965 6851 11023 6857
rect 10965 6817 10977 6851
rect 11011 6848 11023 6851
rect 11681 6851 11704 6857
rect 11681 6848 11693 6851
rect 11011 6820 11693 6848
rect 11011 6817 11023 6820
rect 10965 6811 11023 6817
rect 11681 6817 11693 6820
rect 11756 6848 11762 6860
rect 11756 6820 11829 6848
rect 11681 6811 11704 6817
rect 11698 6808 11704 6811
rect 11756 6808 11762 6820
rect 8478 6780 8484 6792
rect 8439 6752 8484 6780
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 8662 6780 8668 6792
rect 8623 6752 8668 6780
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 9490 6712 9496 6724
rect 9403 6684 9496 6712
rect 9490 6672 9496 6684
rect 9548 6712 9554 6724
rect 10226 6712 10232 6724
rect 9548 6684 10232 6712
rect 9548 6672 9554 6684
rect 10226 6672 10232 6684
rect 10284 6712 10290 6724
rect 10428 6712 10456 6743
rect 10284 6684 10456 6712
rect 10284 6672 10290 6684
rect 934 6604 940 6656
rect 992 6644 998 6656
rect 2225 6647 2283 6653
rect 2225 6644 2237 6647
rect 992 6616 2237 6644
rect 992 6604 998 6616
rect 2225 6613 2237 6616
rect 2271 6613 2283 6647
rect 2225 6607 2283 6613
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 5442 6644 5448 6656
rect 5399 6616 5448 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 6457 6647 6515 6653
rect 6457 6644 6469 6647
rect 6236 6616 6469 6644
rect 6236 6604 6242 6616
rect 6457 6613 6469 6616
rect 6503 6613 6515 6647
rect 6457 6607 6515 6613
rect 8021 6647 8079 6653
rect 8021 6613 8033 6647
rect 8067 6644 8079 6647
rect 8570 6644 8576 6656
rect 8067 6616 8576 6644
rect 8067 6613 8079 6616
rect 8021 6607 8079 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 11238 6644 11244 6656
rect 11199 6616 11244 6644
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11440 6644 11468 6743
rect 11606 6644 11612 6656
rect 11440 6616 11612 6644
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 3326 6440 3332 6452
rect 1811 6412 3332 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 2041 6375 2099 6381
rect 2041 6372 2053 6375
rect 1452 6344 2053 6372
rect 1452 6332 1458 6344
rect 2041 6341 2053 6344
rect 2087 6341 2099 6375
rect 2041 6335 2099 6341
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 2148 6236 2176 6412
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 5166 6440 5172 6452
rect 5127 6412 5172 6440
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6144 6412 6561 6440
rect 6144 6400 6150 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 7558 6440 7564 6452
rect 7519 6412 7564 6440
rect 6549 6403 6607 6409
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8444 6412 9045 6440
rect 8444 6400 8450 6412
rect 9033 6409 9045 6412
rect 9079 6409 9091 6443
rect 9033 6403 9091 6409
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 9950 6440 9956 6452
rect 9732 6412 9956 6440
rect 9732 6400 9738 6412
rect 9950 6400 9956 6412
rect 10008 6440 10014 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 10008 6412 10057 6440
rect 10008 6400 10014 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10502 6440 10508 6452
rect 10463 6412 10508 6440
rect 10045 6403 10103 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10778 6440 10784 6452
rect 10739 6412 10784 6440
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11756 6412 11805 6440
rect 11756 6400 11762 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 3602 6372 3608 6384
rect 3563 6344 3608 6372
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 4982 6332 4988 6384
rect 5040 6372 5046 6384
rect 5813 6375 5871 6381
rect 5813 6372 5825 6375
rect 5040 6344 5825 6372
rect 5040 6332 5046 6344
rect 5813 6341 5825 6344
rect 5859 6341 5871 6375
rect 5813 6335 5871 6341
rect 5994 6332 6000 6384
rect 6052 6372 6058 6384
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 6052 6344 6193 6372
rect 6052 6332 6058 6344
rect 6181 6341 6193 6344
rect 6227 6341 6239 6375
rect 6181 6335 6239 6341
rect 1903 6208 2176 6236
rect 2961 6239 3019 6245
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3620 6236 3648 6332
rect 3007 6208 3648 6236
rect 4433 6239 4491 6245
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4479 6208 4537 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4525 6205 4537 6208
rect 4571 6236 4583 6239
rect 4706 6236 4712 6248
rect 4571 6208 4712 6236
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 5629 6239 5687 6245
rect 5629 6205 5641 6239
rect 5675 6236 5687 6239
rect 6012 6236 6040 6332
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 9398 6304 9404 6316
rect 8619 6276 9404 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 9398 6264 9404 6276
rect 9456 6304 9462 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9456 6276 9505 6304
rect 9456 6264 9462 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 9640 6276 9685 6304
rect 9640 6264 9646 6276
rect 11054 6264 11060 6316
rect 11112 6264 11118 6316
rect 11425 6307 11483 6313
rect 11425 6273 11437 6307
rect 11471 6304 11483 6307
rect 11716 6304 11744 6400
rect 11471 6276 11744 6304
rect 11471 6273 11483 6276
rect 11425 6267 11483 6273
rect 5675 6208 6040 6236
rect 7009 6239 7067 6245
rect 5675 6205 5687 6208
rect 5629 6199 5687 6205
rect 7009 6205 7021 6239
rect 7055 6236 7067 6239
rect 7558 6236 7564 6248
rect 7055 6208 7564 6236
rect 7055 6205 7067 6208
rect 7009 6199 7067 6205
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 11072 6236 11100 6264
rect 11716 6236 11744 6276
rect 13170 6236 13176 6248
rect 11072 6208 11192 6236
rect 11716 6208 13176 6236
rect 11164 6168 11192 6208
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 11974 6168 11980 6180
rect 11164 6140 11980 6168
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 2498 6100 2504 6112
rect 2459 6072 2504 6100
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 3142 6100 3148 6112
rect 3103 6072 3148 6100
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 5810 6100 5816 6112
rect 4755 6072 5816 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 7190 6100 7196 6112
rect 7151 6072 7196 6100
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 8113 6103 8171 6109
rect 8113 6069 8125 6103
rect 8159 6100 8171 6103
rect 8662 6100 8668 6112
rect 8159 6072 8668 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 8941 6103 8999 6109
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 9398 6100 9404 6112
rect 8987 6072 9404 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11296 6072 11341 6100
rect 11296 6060 11302 6072
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 11572 6072 12173 6100
rect 11572 6060 11578 6072
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 12161 6063 12219 6069
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12492 6072 12537 6100
rect 12492 6060 12498 6072
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7834 5896 7840 5908
rect 7607 5868 7840 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 7929 5899 7987 5905
rect 7929 5865 7941 5899
rect 7975 5896 7987 5899
rect 8478 5896 8484 5908
rect 7975 5868 8484 5896
rect 7975 5865 7987 5868
rect 7929 5859 7987 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 9490 5896 9496 5908
rect 9451 5868 9496 5896
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 10686 5896 10692 5908
rect 10647 5868 10692 5896
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 8846 5788 8852 5840
rect 8904 5828 8910 5840
rect 9125 5831 9183 5837
rect 9125 5828 9137 5831
rect 8904 5800 9137 5828
rect 8904 5788 8910 5800
rect 9125 5797 9137 5800
rect 9171 5828 9183 5831
rect 9582 5828 9588 5840
rect 9171 5800 9588 5828
rect 9171 5797 9183 5800
rect 9125 5791 9183 5797
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 2774 5760 2780 5772
rect 2363 5732 2780 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4338 5760 4344 5772
rect 4111 5732 4344 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5960 5732 6009 5760
rect 5960 5720 5966 5732
rect 5997 5729 6009 5732
rect 6043 5729 6055 5763
rect 8386 5760 8392 5772
rect 8347 5732 8392 5760
rect 5997 5723 6055 5729
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 11885 5763 11943 5769
rect 10275 5732 10916 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 10888 5704 10916 5732
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 11974 5760 11980 5772
rect 11931 5732 11980 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 5552 5664 6193 5692
rect 4246 5624 4252 5636
rect 4207 5596 4252 5624
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 5552 5568 5580 5664
rect 6181 5661 6193 5664
rect 6227 5661 6239 5695
rect 6181 5655 6239 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8352 5664 8493 5692
rect 8352 5652 8358 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8662 5692 8668 5704
rect 8623 5664 8668 5692
rect 8481 5655 8539 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9398 5692 9404 5704
rect 8996 5664 9404 5692
rect 8996 5652 9002 5664
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 10778 5692 10784 5704
rect 10739 5664 10784 5692
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 12989 5695 13047 5701
rect 10928 5664 10973 5692
rect 10928 5652 10934 5664
rect 12989 5661 13001 5695
rect 13035 5692 13047 5695
rect 13078 5692 13084 5704
rect 13035 5664 13084 5692
rect 13035 5661 13047 5664
rect 12989 5655 13047 5661
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 5629 5627 5687 5633
rect 5629 5593 5641 5627
rect 5675 5624 5687 5627
rect 7006 5624 7012 5636
rect 5675 5596 7012 5624
rect 5675 5593 5687 5596
rect 5629 5587 5687 5593
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 11054 5624 11060 5636
rect 10980 5596 11060 5624
rect 2222 5516 2228 5568
rect 2280 5556 2286 5568
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 2280 5528 2513 5556
rect 2280 5516 2286 5528
rect 2501 5525 2513 5528
rect 2547 5525 2559 5559
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 2501 5519 2559 5525
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 6917 5559 6975 5565
rect 6917 5556 6929 5559
rect 6880 5528 6929 5556
rect 6880 5516 6886 5528
rect 6917 5525 6929 5528
rect 6963 5525 6975 5559
rect 6917 5519 6975 5525
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8202 5556 8208 5568
rect 8067 5528 8208 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 10980 5556 11008 5596
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 11146 5584 11152 5636
rect 11204 5624 11210 5636
rect 11425 5627 11483 5633
rect 11425 5624 11437 5627
rect 11204 5596 11437 5624
rect 11204 5584 11210 5596
rect 11425 5593 11437 5596
rect 11471 5624 11483 5627
rect 12342 5624 12348 5636
rect 11471 5596 12348 5624
rect 11471 5593 11483 5596
rect 11425 5587 11483 5593
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 12529 5627 12587 5633
rect 12529 5593 12541 5627
rect 12575 5624 12587 5627
rect 13170 5624 13176 5636
rect 12575 5596 13176 5624
rect 12575 5593 12587 5596
rect 12529 5587 12587 5593
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 10367 5528 11008 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 12069 5559 12127 5565
rect 12069 5556 12081 5559
rect 11572 5528 12081 5556
rect 11572 5516 11578 5528
rect 12069 5525 12081 5528
rect 12115 5525 12127 5559
rect 12069 5519 12127 5525
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12768 5528 12817 5556
rect 12768 5516 12774 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 12805 5519 12863 5525
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 2869 5355 2927 5361
rect 2869 5352 2881 5355
rect 2832 5324 2881 5352
rect 2832 5312 2838 5324
rect 2869 5321 2881 5324
rect 2915 5321 2927 5355
rect 4798 5352 4804 5364
rect 4759 5324 4804 5352
rect 2869 5315 2927 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 6086 5352 6092 5364
rect 6047 5324 6092 5352
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 11241 5355 11299 5361
rect 11241 5352 11253 5355
rect 10836 5324 11253 5352
rect 10836 5312 10842 5324
rect 11241 5321 11253 5324
rect 11287 5321 11299 5355
rect 11974 5352 11980 5364
rect 11935 5324 11980 5352
rect 11241 5315 11299 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12618 5352 12624 5364
rect 12483 5324 12624 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 10686 5244 10692 5296
rect 10744 5284 10750 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 10744 5256 11621 5284
rect 10744 5244 10750 5256
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 11609 5247 11667 5253
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13170 5216 13176 5228
rect 13127 5188 13176 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 13446 5176 13452 5228
rect 13504 5216 13510 5228
rect 13722 5216 13728 5228
rect 13504 5188 13728 5216
rect 13504 5176 13510 5188
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5148 2099 5151
rect 2130 5148 2136 5160
rect 2087 5120 2136 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5148 3479 5151
rect 3510 5148 3516 5160
rect 3467 5120 3516 5148
rect 3467 5117 3479 5120
rect 3421 5111 3479 5117
rect 3510 5108 3516 5120
rect 3568 5148 3574 5160
rect 4522 5148 4528 5160
rect 3568 5120 4528 5148
rect 3568 5108 3574 5120
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6822 5148 6828 5160
rect 6052 5120 6828 5148
rect 6052 5108 6058 5120
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 10042 5148 10048 5160
rect 9355 5120 10048 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 10042 5108 10048 5120
rect 10100 5148 10106 5160
rect 11606 5148 11612 5160
rect 10100 5120 11612 5148
rect 10100 5108 10106 5120
rect 11606 5108 11612 5120
rect 11664 5108 11670 5160
rect 3329 5083 3387 5089
rect 3329 5049 3341 5083
rect 3375 5080 3387 5083
rect 3688 5083 3746 5089
rect 3688 5080 3700 5083
rect 3375 5052 3700 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 3688 5049 3700 5052
rect 3734 5080 3746 5083
rect 3970 5080 3976 5092
rect 3734 5052 3976 5080
rect 3734 5049 3746 5052
rect 3688 5043 3746 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 5718 5080 5724 5092
rect 5679 5052 5724 5080
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 6641 5083 6699 5089
rect 6641 5049 6653 5083
rect 6687 5080 6699 5083
rect 7070 5083 7128 5089
rect 7070 5080 7082 5083
rect 6687 5052 7082 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 7070 5049 7082 5052
rect 7116 5080 7128 5083
rect 8018 5080 8024 5092
rect 7116 5052 8024 5080
rect 7116 5049 7128 5052
rect 7070 5043 7128 5049
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 9582 5089 9588 5092
rect 8849 5083 8907 5089
rect 8849 5080 8861 5083
rect 8720 5052 8861 5080
rect 8720 5040 8726 5052
rect 8849 5049 8861 5052
rect 8895 5080 8907 5083
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 8895 5052 9229 5080
rect 8895 5049 8907 5052
rect 8849 5043 8907 5049
rect 9217 5049 9229 5052
rect 9263 5080 9275 5083
rect 9576 5080 9588 5089
rect 9263 5052 9588 5080
rect 9263 5049 9275 5052
rect 9217 5043 9275 5049
rect 9576 5043 9588 5052
rect 9582 5040 9588 5043
rect 9640 5040 9646 5092
rect 12710 5040 12716 5092
rect 12768 5080 12774 5092
rect 12897 5083 12955 5089
rect 12897 5080 12909 5083
rect 12768 5052 12909 5080
rect 12768 5040 12774 5052
rect 12897 5049 12909 5052
rect 12943 5049 12955 5083
rect 12897 5043 12955 5049
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 7432 4984 8217 5012
rect 7432 4972 7438 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 10686 5012 10692 5024
rect 10647 4984 10692 5012
rect 8205 4975 8263 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 12802 5012 12808 5024
rect 12763 4984 12808 5012
rect 12802 4972 12808 4984
rect 12860 5012 12866 5024
rect 13449 5015 13507 5021
rect 13449 5012 13461 5015
rect 12860 4984 13461 5012
rect 12860 4972 12866 4984
rect 13449 4981 13461 4984
rect 13495 4981 13507 5015
rect 13449 4975 13507 4981
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 2409 4811 2467 4817
rect 2409 4808 2421 4811
rect 2188 4780 2421 4808
rect 2188 4768 2194 4780
rect 2409 4777 2421 4780
rect 2455 4777 2467 4811
rect 2409 4771 2467 4777
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 3510 4808 3516 4820
rect 3292 4780 3516 4808
rect 3292 4768 3298 4780
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 4801 4811 4859 4817
rect 4801 4808 4813 4811
rect 4580 4780 4813 4808
rect 4580 4768 4586 4780
rect 4801 4777 4813 4780
rect 4847 4777 4859 4811
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 4801 4771 4859 4777
rect 4816 4740 4844 4771
rect 7006 4768 7012 4780
rect 7064 4808 7070 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7064 4780 7849 4808
rect 7064 4768 7070 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 8260 4780 9321 4808
rect 8260 4768 8266 4780
rect 9309 4777 9321 4780
rect 9355 4808 9367 4811
rect 9674 4808 9680 4820
rect 9355 4780 9680 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10652 4780 10701 4808
rect 10652 4768 10658 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 10689 4771 10747 4777
rect 11238 4768 11244 4820
rect 11296 4808 11302 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11296 4780 11805 4808
rect 11296 4768 11302 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 5994 4740 6000 4752
rect 4816 4712 6000 4740
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 4816 4672 4844 4712
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 12253 4743 12311 4749
rect 12253 4740 12265 4743
rect 11256 4712 12265 4740
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 2832 4644 2877 4672
rect 4816 4644 4997 4672
rect 2832 4632 2838 4644
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 5241 4675 5299 4681
rect 5241 4672 5253 4675
rect 5132 4644 5253 4672
rect 5132 4632 5138 4644
rect 5241 4641 5253 4644
rect 5287 4672 5299 4675
rect 5534 4672 5540 4684
rect 5287 4644 5540 4672
rect 5287 4641 5299 4644
rect 5241 4635 5299 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 6380 4644 8156 4672
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2866 4604 2872 4616
rect 2363 4576 2872 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3970 4604 3976 4616
rect 3099 4576 3976 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 6380 4548 6408 4644
rect 8128 4613 8156 4644
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9306 4672 9312 4684
rect 8720 4644 9312 4672
rect 8720 4632 8726 4644
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 10318 4632 10324 4684
rect 10376 4672 10382 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 10376 4644 10609 4672
rect 10376 4632 10382 4644
rect 10597 4641 10609 4644
rect 10643 4672 10655 4675
rect 10778 4672 10784 4684
rect 10643 4644 10784 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11256 4681 11284 4712
rect 12253 4709 12265 4712
rect 12299 4709 12311 4743
rect 12253 4703 12311 4709
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 11112 4644 11253 4672
rect 11112 4632 11118 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12805 4675 12863 4681
rect 12805 4672 12817 4675
rect 12207 4644 12817 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12805 4641 12817 4644
rect 12851 4641 12863 4675
rect 12805 4635 12863 4641
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8478 4604 8484 4616
rect 8159 4576 8484 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 6362 4536 6368 4548
rect 6275 4508 6368 4536
rect 6362 4496 6368 4508
rect 6420 4496 6426 4548
rect 7466 4536 7472 4548
rect 7427 4508 7472 4536
rect 7466 4496 7472 4508
rect 7524 4496 7530 4548
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 7282 4468 7288 4480
rect 7243 4440 7288 4468
rect 7282 4428 7288 4440
rect 7340 4468 7346 4480
rect 7944 4468 7972 4567
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 12176 4604 12204 4635
rect 12894 4632 12900 4684
rect 12952 4672 12958 4684
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 12952 4644 13369 4672
rect 12952 4632 12958 4644
rect 13357 4641 13369 4644
rect 13403 4672 13415 4675
rect 13446 4672 13452 4684
rect 13403 4644 13452 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 11020 4576 12204 4604
rect 11020 4564 11026 4576
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12492 4576 12537 4604
rect 12492 4564 12498 4576
rect 8386 4496 8392 4548
rect 8444 4536 8450 4548
rect 8849 4539 8907 4545
rect 8849 4536 8861 4539
rect 8444 4508 8861 4536
rect 8444 4496 8450 4508
rect 8849 4505 8861 4508
rect 8895 4505 8907 4539
rect 8849 4499 8907 4505
rect 10229 4539 10287 4545
rect 10229 4505 10241 4539
rect 10275 4536 10287 4539
rect 12894 4536 12900 4548
rect 10275 4508 12900 4536
rect 10275 4505 10287 4508
rect 10229 4499 10287 4505
rect 12894 4496 12900 4508
rect 12952 4536 12958 4548
rect 13173 4539 13231 4545
rect 13173 4536 13185 4539
rect 12952 4508 13185 4536
rect 12952 4496 12958 4508
rect 13173 4505 13185 4508
rect 13219 4505 13231 4539
rect 13173 4499 13231 4505
rect 7340 4440 7972 4468
rect 7340 4428 7346 4440
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 8352 4440 8493 4468
rect 8352 4428 8358 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 8481 4431 8539 4437
rect 9953 4471 10011 4477
rect 9953 4437 9965 4471
rect 9999 4468 10011 4471
rect 10042 4468 10048 4480
rect 9999 4440 10048 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 11701 4471 11759 4477
rect 11701 4437 11713 4471
rect 11747 4468 11759 4471
rect 11974 4468 11980 4480
rect 11747 4440 11980 4468
rect 11747 4437 11759 4440
rect 11701 4431 11759 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 13538 4468 13544 4480
rect 13499 4440 13544 4468
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2501 4267 2559 4273
rect 2501 4233 2513 4267
rect 2547 4264 2559 4267
rect 3970 4264 3976 4276
rect 2547 4236 3976 4264
rect 2547 4233 2559 4236
rect 2501 4227 2559 4233
rect 3970 4224 3976 4236
rect 4028 4264 4034 4276
rect 4433 4267 4491 4273
rect 4433 4264 4445 4267
rect 4028 4236 4445 4264
rect 4028 4224 4034 4236
rect 4433 4233 4445 4236
rect 4479 4233 4491 4267
rect 4433 4227 4491 4233
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 10413 4267 10471 4273
rect 10413 4264 10425 4267
rect 9824 4236 10425 4264
rect 9824 4224 9830 4236
rect 10413 4233 10425 4236
rect 10459 4264 10471 4267
rect 10594 4264 10600 4276
rect 10459 4236 10600 4264
rect 10459 4233 10471 4236
rect 10413 4227 10471 4233
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 10778 4264 10784 4276
rect 10739 4236 10784 4264
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 11882 4224 11888 4276
rect 11940 4264 11946 4276
rect 12069 4267 12127 4273
rect 12069 4264 12081 4267
rect 11940 4236 12081 4264
rect 11940 4224 11946 4236
rect 12069 4233 12081 4236
rect 12115 4264 12127 4267
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 12115 4236 12173 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 12437 4267 12495 4273
rect 12437 4264 12449 4267
rect 12400 4236 12449 4264
rect 12400 4224 12406 4236
rect 12437 4233 12449 4236
rect 12483 4233 12495 4267
rect 13446 4264 13452 4276
rect 13407 4236 13452 4264
rect 12437 4227 12495 4233
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 8018 4156 8024 4208
rect 8076 4196 8082 4208
rect 10686 4196 10692 4208
rect 8076 4168 8248 4196
rect 8076 4156 8082 4168
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6052 4100 6837 4128
rect 6052 4088 6058 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 8220 4128 8248 4168
rect 9876 4168 10692 4196
rect 9876 4137 9904 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8220 4100 9137 4128
rect 6825 4091 6883 4097
rect 9125 4097 9137 4100
rect 9171 4128 9183 4131
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9171 4100 9873 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 12066 4128 12072 4140
rect 9861 4091 9919 4097
rect 11900 4100 12072 4128
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1670 4060 1676 4072
rect 1443 4032 1676 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1670 4020 1676 4032
rect 1728 4020 1734 4072
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4060 3111 4063
rect 3142 4060 3148 4072
rect 3099 4032 3148 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3326 4069 3332 4072
rect 3320 4060 3332 4069
rect 3252 4032 3332 4060
rect 2961 3995 3019 4001
rect 2961 3961 2973 3995
rect 3007 3992 3019 3995
rect 3252 3992 3280 4032
rect 3320 4023 3332 4032
rect 3326 4020 3332 4023
rect 3384 4020 3390 4072
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4060 5595 4063
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 5583 4032 6193 4060
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 6181 4029 6193 4032
rect 6227 4060 6239 4063
rect 6270 4060 6276 4072
rect 6227 4032 6276 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 7092 4063 7150 4069
rect 7092 4060 7104 4063
rect 7024 4032 7104 4060
rect 5074 3992 5080 4004
rect 3007 3964 3280 3992
rect 4987 3964 5080 3992
rect 3007 3961 3019 3964
rect 2961 3955 3019 3961
rect 5074 3952 5080 3964
rect 5132 3992 5138 4004
rect 5445 3995 5503 4001
rect 5445 3992 5457 3995
rect 5132 3964 5457 3992
rect 5132 3952 5138 3964
rect 5445 3961 5457 3964
rect 5491 3992 5503 3995
rect 6641 3995 6699 4001
rect 5491 3964 6592 3992
rect 5491 3961 5503 3964
rect 5445 3955 5503 3961
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6564 3924 6592 3964
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 6730 3992 6736 4004
rect 6687 3964 6736 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 6730 3952 6736 3964
rect 6788 3992 6794 4004
rect 7024 3992 7052 4032
rect 7092 4029 7104 4032
rect 7138 4060 7150 4063
rect 7374 4060 7380 4072
rect 7138 4032 7380 4060
rect 7138 4029 7150 4032
rect 7092 4023 7150 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8536 4032 8769 4060
rect 8536 4020 8542 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 9490 4060 9496 4072
rect 8757 4023 8815 4029
rect 9140 4032 9496 4060
rect 9140 4004 9168 4032
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 9674 4060 9680 4072
rect 9635 4032 9680 4060
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10873 4063 10931 4069
rect 10873 4060 10885 4063
rect 10836 4032 10885 4060
rect 10836 4020 10842 4032
rect 10873 4029 10885 4032
rect 10919 4060 10931 4063
rect 11425 4063 11483 4069
rect 11425 4060 11437 4063
rect 10919 4032 11437 4060
rect 10919 4029 10931 4032
rect 10873 4023 10931 4029
rect 11425 4029 11437 4032
rect 11471 4060 11483 4063
rect 11900 4060 11928 4100
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12894 4128 12900 4140
rect 12855 4100 12900 4128
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13446 4128 13452 4140
rect 13127 4100 13452 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 11471 4032 11928 4060
rect 11471 4029 11483 4032
rect 11425 4023 11483 4029
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12434 4060 12440 4072
rect 12032 4032 12440 4060
rect 12032 4020 12038 4032
rect 12434 4020 12440 4032
rect 12492 4060 12498 4072
rect 13096 4060 13124 4091
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 12492 4032 13124 4060
rect 12492 4020 12498 4032
rect 6788 3964 7052 3992
rect 6788 3952 6794 3964
rect 9122 3952 9128 4004
rect 9180 3952 9186 4004
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 6564 3896 8217 3924
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 9306 3924 9312 3936
rect 9267 3896 9312 3924
rect 8205 3887 8263 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9548 3896 9781 3924
rect 9548 3884 9554 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 11054 3924 11060 3936
rect 11015 3896 11060 3924
rect 9769 3887 9827 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 11974 3924 11980 3936
rect 11931 3896 11980 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 12069 3927 12127 3933
rect 12069 3893 12081 3927
rect 12115 3924 12127 3927
rect 12342 3924 12348 3936
rect 12115 3896 12348 3924
rect 12115 3893 12127 3896
rect 12069 3887 12127 3893
rect 12342 3884 12348 3896
rect 12400 3924 12406 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 12400 3896 12817 3924
rect 12400 3884 12406 3896
rect 12805 3893 12817 3896
rect 12851 3893 12863 3927
rect 12805 3887 12863 3893
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 2409 3723 2467 3729
rect 2409 3720 2421 3723
rect 1995 3692 2421 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 2409 3689 2421 3692
rect 2455 3720 2467 3723
rect 2682 3720 2688 3732
rect 2455 3692 2688 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3292 3692 3433 3720
rect 3292 3680 3298 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 4525 3723 4583 3729
rect 4525 3689 4537 3723
rect 4571 3720 4583 3723
rect 5445 3723 5503 3729
rect 5445 3720 5457 3723
rect 4571 3692 5457 3720
rect 4571 3689 4583 3692
rect 4525 3683 4583 3689
rect 5445 3689 5457 3692
rect 5491 3720 5503 3723
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 5491 3692 6561 3720
rect 5491 3689 5503 3692
rect 5445 3683 5503 3689
rect 6549 3689 6561 3692
rect 6595 3689 6607 3723
rect 6549 3683 6607 3689
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 7009 3723 7067 3729
rect 7009 3720 7021 3723
rect 6880 3692 7021 3720
rect 6880 3680 6886 3692
rect 7009 3689 7021 3692
rect 7055 3720 7067 3723
rect 7190 3720 7196 3732
rect 7055 3692 7196 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7926 3720 7932 3732
rect 7887 3692 7932 3720
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 9309 3723 9367 3729
rect 9309 3720 9321 3723
rect 8628 3692 9321 3720
rect 8628 3680 8634 3692
rect 9309 3689 9321 3692
rect 9355 3720 9367 3723
rect 9490 3720 9496 3732
rect 9355 3692 9496 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 9858 3720 9864 3732
rect 9819 3692 9864 3720
rect 9858 3680 9864 3692
rect 9916 3720 9922 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 9916 3692 10425 3720
rect 9916 3680 9922 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13170 3720 13176 3732
rect 13035 3692 13176 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 4893 3655 4951 3661
rect 4893 3621 4905 3655
rect 4939 3652 4951 3655
rect 5074 3652 5080 3664
rect 4939 3624 5080 3652
rect 4939 3621 4951 3624
rect 4893 3615 4951 3621
rect 5074 3612 5080 3624
rect 5132 3652 5138 3664
rect 5994 3652 6000 3664
rect 5132 3624 5488 3652
rect 5955 3624 6000 3652
rect 5132 3612 5138 3624
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3584 2375 3587
rect 2777 3587 2835 3593
rect 2777 3584 2789 3587
rect 2363 3556 2789 3584
rect 2363 3553 2375 3556
rect 2317 3547 2375 3553
rect 2777 3553 2789 3556
rect 2823 3584 2835 3587
rect 3418 3584 3424 3596
rect 2823 3556 3424 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 4764 3556 5365 3584
rect 4764 3544 4770 3556
rect 5353 3553 5365 3556
rect 5399 3553 5411 3587
rect 5353 3547 5411 3553
rect 5460 3528 5488 3624
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 6457 3655 6515 3661
rect 6457 3621 6469 3655
rect 6503 3652 6515 3655
rect 6730 3652 6736 3664
rect 6503 3624 6736 3652
rect 6503 3621 6515 3624
rect 6457 3615 6515 3621
rect 6730 3612 6736 3624
rect 6788 3652 6794 3664
rect 7653 3655 7711 3661
rect 6788 3624 7144 3652
rect 6788 3612 6794 3624
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 6963 3556 7052 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3516 1455 3519
rect 2682 3516 2688 3528
rect 1443 3488 2688 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3516 2872 3528
rect 2827 3488 2872 3516
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3326 3516 3332 3528
rect 3099 3488 3332 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 5442 3516 5448 3528
rect 5355 3488 5448 3516
rect 5442 3476 5448 3488
rect 5500 3516 5506 3528
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 5500 3488 5549 3516
rect 5500 3476 5506 3488
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 7024 3460 7052 3556
rect 7116 3525 7144 3624
rect 7653 3621 7665 3655
rect 7699 3652 7711 3655
rect 7834 3652 7840 3664
rect 7699 3624 7840 3652
rect 7699 3621 7711 3624
rect 7653 3615 7711 3621
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 8846 3652 8852 3664
rect 8807 3624 8852 3652
rect 8846 3612 8852 3624
rect 8904 3612 8910 3664
rect 11517 3655 11575 3661
rect 11517 3621 11529 3655
rect 11563 3652 11575 3655
rect 11876 3655 11934 3661
rect 11876 3652 11888 3655
rect 11563 3624 11888 3652
rect 11563 3621 11575 3624
rect 11517 3615 11575 3621
rect 11876 3621 11888 3624
rect 11922 3652 11934 3655
rect 11974 3652 11980 3664
rect 11922 3624 11980 3652
rect 11922 3621 11934 3624
rect 11876 3615 11934 3621
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 8386 3584 8392 3596
rect 8159 3556 8392 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 8386 3544 8392 3556
rect 8444 3584 8450 3596
rect 8754 3584 8760 3596
rect 8444 3556 8760 3584
rect 8444 3544 8450 3556
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 10505 3519 10563 3525
rect 10505 3516 10517 3519
rect 10468 3488 10517 3516
rect 10468 3476 10474 3488
rect 10505 3485 10517 3488
rect 10551 3485 10563 3519
rect 10686 3516 10692 3528
rect 10647 3488 10692 3516
rect 10505 3479 10563 3485
rect 10686 3476 10692 3488
rect 10744 3516 10750 3528
rect 10870 3516 10876 3528
rect 10744 3488 10876 3516
rect 10744 3476 10750 3488
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10928 3488 11069 3516
rect 10928 3476 10934 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11606 3516 11612 3528
rect 11567 3488 11612 3516
rect 11057 3479 11115 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 4985 3451 5043 3457
rect 4985 3417 4997 3451
rect 5031 3448 5043 3451
rect 5350 3448 5356 3460
rect 5031 3420 5356 3448
rect 5031 3417 5043 3420
rect 4985 3411 5043 3417
rect 5350 3408 5356 3420
rect 5408 3408 5414 3460
rect 7006 3448 7012 3460
rect 6919 3420 7012 3448
rect 7006 3408 7012 3420
rect 7064 3448 7070 3460
rect 7558 3448 7564 3460
rect 7064 3420 7564 3448
rect 7064 3408 7070 3420
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 10045 3451 10103 3457
rect 10045 3417 10057 3451
rect 10091 3448 10103 3451
rect 10962 3448 10968 3460
rect 10091 3420 10968 3448
rect 10091 3417 10103 3420
rect 10045 3411 10103 3417
rect 10962 3408 10968 3420
rect 11020 3408 11026 3460
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 5074 3380 5080 3392
rect 4212 3352 5080 3380
rect 4212 3340 4218 3352
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 8294 3380 8300 3392
rect 8255 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 2866 3176 2872 3188
rect 1719 3148 2872 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 2866 3136 2872 3148
rect 2924 3176 2930 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 2924 3148 4905 3176
rect 2924 3136 2930 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 6822 3176 6828 3188
rect 6687 3148 6828 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 8202 3176 8208 3188
rect 7239 3148 8208 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8386 3176 8392 3188
rect 8343 3148 8392 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 8754 3176 8760 3188
rect 8711 3148 8760 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10137 3179 10195 3185
rect 10137 3176 10149 3179
rect 9732 3148 10149 3176
rect 9732 3136 9738 3148
rect 10137 3145 10149 3148
rect 10183 3145 10195 3179
rect 10137 3139 10195 3145
rect 10410 3136 10416 3188
rect 10468 3176 10474 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 10468 3148 10701 3176
rect 10468 3136 10474 3148
rect 10689 3145 10701 3148
rect 10735 3145 10747 3179
rect 10689 3139 10747 3145
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11330 3176 11336 3188
rect 11195 3148 11336 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 11330 3136 11336 3148
rect 11388 3176 11394 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11388 3148 11805 3176
rect 11388 3136 11394 3148
rect 11793 3145 11805 3148
rect 11839 3145 11851 3179
rect 11793 3139 11851 3145
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 12710 3176 12716 3188
rect 12483 3148 12716 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 4433 3111 4491 3117
rect 4433 3077 4445 3111
rect 4479 3108 4491 3111
rect 4706 3108 4712 3120
rect 4479 3080 4712 3108
rect 4479 3077 4491 3080
rect 4433 3071 4491 3077
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 6840 3108 6868 3136
rect 8113 3111 8171 3117
rect 8113 3108 8125 3111
rect 6840 3080 8125 3108
rect 8113 3077 8125 3080
rect 8159 3077 8171 3111
rect 8113 3071 8171 3077
rect 10226 3068 10232 3120
rect 10284 3108 10290 3120
rect 10962 3108 10968 3120
rect 10284 3080 10968 3108
rect 10284 3068 10290 3080
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 11425 3111 11483 3117
rect 11425 3108 11437 3111
rect 11112 3080 11437 3108
rect 11112 3068 11118 3080
rect 11425 3077 11437 3080
rect 11471 3077 11483 3111
rect 11808 3108 11836 3139
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 11808 3080 12940 3108
rect 11425 3071 11483 3077
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 4890 3040 4896 3052
rect 4847 3012 4896 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 4890 3000 4896 3012
rect 4948 3040 4954 3052
rect 5442 3040 5448 3052
rect 4948 3012 5304 3040
rect 5403 3012 5448 3040
rect 4948 3000 4954 3012
rect 5276 2984 5304 3012
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 12912 3049 12940 3080
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 6880 3012 7849 3040
rect 6880 3000 6886 3012
rect 7837 3009 7849 3012
rect 7883 3040 7895 3043
rect 12897 3043 12955 3049
rect 7883 3012 8892 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8864 2984 8892 3012
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13446 3040 13452 3052
rect 13127 3012 13452 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 1728 2944 2145 2972
rect 1728 2932 1734 2944
rect 2133 2941 2145 2944
rect 2179 2972 2191 2975
rect 3234 2972 3240 2984
rect 2179 2944 3240 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 5258 2972 5264 2984
rect 5171 2944 5264 2972
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7926 2972 7932 2984
rect 7607 2944 7932 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2972 8171 2975
rect 8202 2972 8208 2984
rect 8159 2944 8208 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 1946 2904 1952 2916
rect 1907 2876 1952 2904
rect 1946 2864 1952 2876
rect 2004 2904 2010 2916
rect 2378 2907 2436 2913
rect 2378 2904 2390 2907
rect 2004 2876 2390 2904
rect 2004 2864 2010 2876
rect 2378 2873 2390 2876
rect 2424 2873 2436 2907
rect 2378 2867 2436 2873
rect 4430 2864 4436 2916
rect 4488 2904 4494 2916
rect 5353 2907 5411 2913
rect 5353 2904 5365 2907
rect 4488 2876 5365 2904
rect 4488 2864 4494 2876
rect 5353 2873 5365 2876
rect 5399 2904 5411 2907
rect 5905 2907 5963 2913
rect 5905 2904 5917 2907
rect 5399 2876 5917 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 5905 2873 5917 2876
rect 5951 2904 5963 2907
rect 6086 2904 6092 2916
rect 5951 2876 6092 2904
rect 5951 2873 5963 2876
rect 5905 2867 5963 2873
rect 6086 2864 6092 2876
rect 6144 2864 6150 2916
rect 7653 2907 7711 2913
rect 7653 2873 7665 2907
rect 7699 2904 7711 2907
rect 7834 2904 7840 2916
rect 7699 2876 7840 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 7834 2864 7840 2876
rect 7892 2864 7898 2916
rect 8772 2904 8800 2935
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 9013 2975 9071 2981
rect 9013 2972 9025 2975
rect 8904 2944 9025 2972
rect 8904 2932 8910 2944
rect 9013 2941 9025 2944
rect 9059 2941 9071 2975
rect 11238 2972 11244 2984
rect 11199 2944 11244 2972
rect 9013 2935 9071 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 13814 2972 13820 2984
rect 13775 2944 13820 2972
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 9582 2904 9588 2916
rect 8772 2876 9588 2904
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 12253 2907 12311 2913
rect 12253 2873 12265 2907
rect 12299 2904 12311 2907
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 12299 2876 12817 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 12805 2873 12817 2876
rect 12851 2904 12863 2907
rect 13722 2904 13728 2916
rect 12851 2876 13728 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 3510 2836 3516 2848
rect 3471 2808 3516 2836
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 13446 2836 13452 2848
rect 13407 2808 13452 2836
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 1670 2632 1676 2644
rect 1631 2604 1676 2632
rect 1670 2592 1676 2604
rect 1728 2592 1734 2644
rect 2406 2632 2412 2644
rect 2367 2604 2412 2632
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 3326 2632 3332 2644
rect 2823 2604 3332 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 4893 2635 4951 2641
rect 4893 2632 4905 2635
rect 3476 2604 4905 2632
rect 3476 2592 3482 2604
rect 4893 2601 4905 2604
rect 4939 2601 4951 2635
rect 4893 2595 4951 2601
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5224 2604 5365 2632
rect 5224 2592 5230 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6822 2632 6828 2644
rect 6411 2604 6828 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 10778 2632 10784 2644
rect 8619 2604 10784 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 2424 2496 2452 2592
rect 4338 2564 4344 2576
rect 4299 2536 4344 2564
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 4801 2567 4859 2573
rect 4801 2533 4813 2567
rect 4847 2564 4859 2567
rect 5184 2564 5212 2592
rect 4847 2536 5212 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 6086 2524 6092 2576
rect 6144 2564 6150 2576
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 6144 2536 6653 2564
rect 6144 2524 6150 2536
rect 6641 2533 6653 2536
rect 6687 2564 6699 2567
rect 7653 2567 7711 2573
rect 6687 2536 6960 2564
rect 6687 2533 6699 2536
rect 6641 2527 6699 2533
rect 1811 2468 2452 2496
rect 2869 2499 2927 2505
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 4356 2496 4384 2524
rect 6932 2505 6960 2536
rect 7653 2533 7665 2567
rect 7699 2564 7711 2567
rect 8588 2564 8616 2595
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 11974 2632 11980 2644
rect 11471 2604 11980 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12621 2635 12679 2641
rect 12621 2601 12633 2635
rect 12667 2632 12679 2635
rect 12802 2632 12808 2644
rect 12667 2604 12808 2632
rect 12667 2601 12679 2604
rect 12621 2595 12679 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 13078 2632 13084 2644
rect 13035 2604 13084 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 7699 2536 8616 2564
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 9122 2524 9128 2576
rect 9180 2564 9186 2576
rect 9217 2567 9275 2573
rect 9217 2564 9229 2567
rect 9180 2536 9229 2564
rect 9180 2524 9186 2536
rect 9217 2533 9229 2536
rect 9263 2564 9275 2567
rect 9585 2567 9643 2573
rect 9585 2564 9597 2567
rect 9263 2536 9597 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 9585 2533 9597 2536
rect 9631 2564 9643 2567
rect 10290 2567 10348 2573
rect 10290 2564 10302 2567
rect 9631 2536 10302 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 10290 2533 10302 2536
rect 10336 2564 10348 2567
rect 10686 2564 10692 2576
rect 10336 2536 10692 2564
rect 10336 2533 10348 2536
rect 10290 2527 10348 2533
rect 10686 2524 10692 2536
rect 10744 2524 10750 2576
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 13004 2564 13032 2595
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 13872 2604 14013 2632
rect 13872 2592 13878 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 14001 2595 14059 2601
rect 13630 2564 13636 2576
rect 12115 2536 13032 2564
rect 13096 2536 13636 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 5261 2499 5319 2505
rect 5261 2496 5273 2499
rect 4356 2468 5273 2496
rect 2869 2459 2927 2465
rect 5261 2465 5273 2468
rect 5307 2465 5319 2499
rect 5261 2459 5319 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 2884 2428 2912 2459
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 8478 2496 8484 2508
rect 7984 2468 8484 2496
rect 7984 2456 7990 2468
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 13096 2505 13124 2536
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 10045 2499 10103 2505
rect 10045 2496 10057 2499
rect 9732 2468 10057 2496
rect 9732 2456 9738 2468
rect 10045 2465 10057 2468
rect 10091 2465 10103 2499
rect 10045 2459 10103 2465
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 12483 2468 13093 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 13081 2465 13093 2468
rect 13127 2465 13139 2499
rect 13081 2459 13139 2465
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 2884 2400 3525 2428
rect 3513 2397 3525 2400
rect 3559 2428 3571 2431
rect 4614 2428 4620 2440
rect 3559 2400 4620 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5500 2400 5917 2428
rect 5500 2388 5506 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 8754 2428 8760 2440
rect 8715 2400 8760 2428
rect 5905 2391 5963 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 13446 2428 13452 2440
rect 13311 2400 13452 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13446 2388 13452 2400
rect 13504 2428 13510 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13504 2400 13645 2428
rect 13504 2388 13510 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 1949 2363 2007 2369
rect 1949 2329 1961 2363
rect 1995 2360 2007 2363
rect 2958 2360 2964 2372
rect 1995 2332 2964 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 2958 2320 2964 2332
rect 3016 2320 3022 2372
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 3326 2292 3332 2304
rect 3099 2264 3332 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 3326 2252 3332 2264
rect 3384 2252 3390 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 5810 552 5816 604
rect 5868 592 5874 604
rect 6914 592 6920 604
rect 5868 564 6920 592
rect 5868 552 5874 564
rect 6914 552 6920 564
rect 6972 552 6978 604
rect 7374 552 7380 604
rect 7432 592 7438 604
rect 8018 592 8024 604
rect 7432 564 8024 592
rect 7432 552 7438 564
rect 8018 552 8024 564
rect 8076 552 8082 604
rect 10318 552 10324 604
rect 10376 592 10382 604
rect 10594 592 10600 604
rect 10376 564 10600 592
rect 10376 552 10382 564
rect 10594 552 10600 564
rect 10652 552 10658 604
rect 12158 552 12164 604
rect 12216 592 12222 604
rect 12342 592 12348 604
rect 12216 564 12348 592
rect 12216 552 12222 564
rect 12342 552 12348 564
rect 12400 552 12406 604
rect 12986 552 12992 604
rect 13044 592 13050 604
rect 13262 592 13268 604
rect 13044 564 13268 592
rect 13044 552 13050 564
rect 13262 552 13268 564
rect 13320 552 13326 604
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 11612 36184 11664 36236
rect 11428 36116 11480 36168
rect 12440 35980 12492 36032
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 204 35776 256 35828
rect 1308 35776 1360 35828
rect 6920 35776 6972 35828
rect 8484 35819 8536 35828
rect 8484 35785 8493 35819
rect 8493 35785 8527 35819
rect 8527 35785 8536 35819
rect 8484 35776 8536 35785
rect 11612 35819 11664 35828
rect 11612 35785 11621 35819
rect 11621 35785 11655 35819
rect 11655 35785 11664 35819
rect 11612 35776 11664 35785
rect 11980 35776 12032 35828
rect 10048 35572 10100 35624
rect 11428 35504 11480 35556
rect 8024 35436 8076 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 1768 35232 1820 35284
rect 3976 35232 4028 35284
rect 5448 35232 5500 35284
rect 7380 35232 7432 35284
rect 9864 35164 9916 35216
rect 2412 35096 2464 35148
rect 4068 35139 4120 35148
rect 4068 35105 4077 35139
rect 4077 35105 4111 35139
rect 4111 35105 4120 35139
rect 4068 35096 4120 35105
rect 5172 35139 5224 35148
rect 5172 35105 5181 35139
rect 5181 35105 5215 35139
rect 5215 35105 5224 35139
rect 5172 35096 5224 35105
rect 6736 35096 6788 35148
rect 7472 35139 7524 35148
rect 7472 35105 7481 35139
rect 7481 35105 7515 35139
rect 7515 35105 7524 35139
rect 7472 35096 7524 35105
rect 11428 35096 11480 35148
rect 4160 34960 4212 35012
rect 5724 34935 5776 34944
rect 5724 34901 5733 34935
rect 5733 34901 5767 34935
rect 5767 34901 5776 34935
rect 5724 34892 5776 34901
rect 8116 34935 8168 34944
rect 8116 34901 8125 34935
rect 8125 34901 8159 34935
rect 8159 34901 8168 34935
rect 8116 34892 8168 34901
rect 11152 34892 11204 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 572 34688 624 34740
rect 2044 34731 2096 34740
rect 2044 34697 2053 34731
rect 2053 34697 2087 34731
rect 2087 34697 2096 34731
rect 2044 34688 2096 34697
rect 2596 34688 2648 34740
rect 6184 34688 6236 34740
rect 6644 34688 6696 34740
rect 7472 34688 7524 34740
rect 8300 34688 8352 34740
rect 9864 34688 9916 34740
rect 10324 34731 10376 34740
rect 10324 34697 10333 34731
rect 10333 34697 10367 34731
rect 10367 34697 10376 34731
rect 13636 34731 13688 34740
rect 10324 34688 10376 34697
rect 1400 34620 1452 34672
rect 2412 34595 2464 34604
rect 2412 34561 2421 34595
rect 2421 34561 2455 34595
rect 2455 34561 2464 34595
rect 2412 34552 2464 34561
rect 2596 34552 2648 34604
rect 3332 34552 3384 34604
rect 4160 34552 4212 34604
rect 2044 34484 2096 34536
rect 3240 34484 3292 34536
rect 4896 34620 4948 34672
rect 13636 34697 13645 34731
rect 13645 34697 13679 34731
rect 13679 34697 13688 34731
rect 13636 34688 13688 34697
rect 11152 34595 11204 34604
rect 11152 34561 11161 34595
rect 11161 34561 11195 34595
rect 11195 34561 11204 34595
rect 11152 34552 11204 34561
rect 5724 34484 5776 34536
rect 6736 34484 6788 34536
rect 7196 34484 7248 34536
rect 7932 34484 7984 34536
rect 9956 34527 10008 34536
rect 9956 34493 9965 34527
rect 9965 34493 9999 34527
rect 9999 34493 10008 34527
rect 9956 34484 10008 34493
rect 13452 34527 13504 34536
rect 13452 34493 13461 34527
rect 13461 34493 13495 34527
rect 13495 34493 13504 34527
rect 13452 34484 13504 34493
rect 4344 34416 4396 34468
rect 5172 34459 5224 34468
rect 5172 34425 5181 34459
rect 5181 34425 5215 34459
rect 5215 34425 5224 34459
rect 5172 34416 5224 34425
rect 8116 34416 8168 34468
rect 8576 34416 8628 34468
rect 4068 34348 4120 34400
rect 5264 34348 5316 34400
rect 10508 34391 10560 34400
rect 10508 34357 10517 34391
rect 10517 34357 10551 34391
rect 10551 34357 10560 34391
rect 10508 34348 10560 34357
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 1400 34144 1452 34196
rect 2136 34144 2188 34196
rect 4160 34144 4212 34196
rect 4988 34144 5040 34196
rect 6920 34187 6972 34196
rect 6920 34153 6929 34187
rect 6929 34153 6963 34187
rect 6963 34153 6972 34187
rect 6920 34144 6972 34153
rect 7748 34144 7800 34196
rect 9864 34187 9916 34196
rect 9864 34153 9873 34187
rect 9873 34153 9907 34187
rect 9907 34153 9916 34187
rect 9864 34144 9916 34153
rect 11980 34144 12032 34196
rect 1952 34008 2004 34060
rect 3332 34008 3384 34060
rect 4068 34051 4120 34060
rect 4068 34017 4077 34051
rect 4077 34017 4111 34051
rect 4111 34017 4120 34051
rect 4068 34008 4120 34017
rect 5448 34008 5500 34060
rect 6644 34008 6696 34060
rect 7564 34008 7616 34060
rect 11152 34008 11204 34060
rect 6828 33804 6880 33856
rect 7932 33804 7984 33856
rect 8300 33804 8352 33856
rect 11428 33804 11480 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 940 33600 992 33652
rect 1952 33643 2004 33652
rect 1952 33609 1961 33643
rect 1961 33609 1995 33643
rect 1995 33609 2004 33643
rect 1952 33600 2004 33609
rect 2964 33643 3016 33652
rect 2964 33609 2973 33643
rect 2973 33609 3007 33643
rect 3007 33609 3016 33643
rect 2964 33600 3016 33609
rect 11152 33643 11204 33652
rect 11152 33609 11161 33643
rect 11161 33609 11195 33643
rect 11195 33609 11204 33643
rect 11152 33600 11204 33609
rect 6828 33507 6880 33516
rect 6828 33473 6837 33507
rect 6837 33473 6871 33507
rect 6871 33473 6880 33507
rect 6828 33464 6880 33473
rect 10508 33464 10560 33516
rect 10784 33507 10836 33516
rect 10784 33473 10793 33507
rect 10793 33473 10827 33507
rect 10827 33473 10836 33507
rect 10784 33464 10836 33473
rect 11980 33464 12032 33516
rect 2780 33439 2832 33448
rect 2780 33405 2789 33439
rect 2789 33405 2823 33439
rect 2823 33405 2832 33439
rect 2780 33396 2832 33405
rect 7380 33328 7432 33380
rect 9864 33328 9916 33380
rect 2412 33303 2464 33312
rect 2412 33269 2421 33303
rect 2421 33269 2455 33303
rect 2455 33269 2464 33303
rect 2412 33260 2464 33269
rect 3332 33303 3384 33312
rect 3332 33269 3341 33303
rect 3341 33269 3375 33303
rect 3375 33269 3384 33303
rect 3332 33260 3384 33269
rect 4068 33260 4120 33312
rect 4712 33260 4764 33312
rect 5448 33260 5500 33312
rect 6644 33303 6696 33312
rect 6644 33269 6653 33303
rect 6653 33269 6687 33303
rect 6687 33269 6696 33303
rect 6644 33260 6696 33269
rect 7288 33260 7340 33312
rect 8208 33303 8260 33312
rect 8208 33269 8217 33303
rect 8217 33269 8251 33303
rect 8251 33269 8260 33303
rect 8208 33260 8260 33269
rect 10140 33303 10192 33312
rect 10140 33269 10149 33303
rect 10149 33269 10183 33303
rect 10183 33269 10192 33303
rect 10140 33260 10192 33269
rect 11428 33260 11480 33312
rect 12256 33260 12308 33312
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 2780 33099 2832 33108
rect 2780 33065 2789 33099
rect 2789 33065 2823 33099
rect 2823 33065 2832 33099
rect 2780 33056 2832 33065
rect 6828 33099 6880 33108
rect 6828 33065 6837 33099
rect 6837 33065 6871 33099
rect 6871 33065 6880 33099
rect 6828 33056 6880 33065
rect 7564 33056 7616 33108
rect 10784 33056 10836 33108
rect 1492 32988 1544 33040
rect 12256 33031 12308 33040
rect 12256 32997 12265 33031
rect 12265 32997 12299 33031
rect 12299 32997 12308 33031
rect 12256 32988 12308 32997
rect 1768 32920 1820 32972
rect 5816 32920 5868 32972
rect 8392 32963 8444 32972
rect 8392 32929 8401 32963
rect 8401 32929 8435 32963
rect 8435 32929 8444 32963
rect 8392 32920 8444 32929
rect 10508 32920 10560 32972
rect 13544 32920 13596 32972
rect 7380 32852 7432 32904
rect 8484 32895 8536 32904
rect 8484 32861 8493 32895
rect 8493 32861 8527 32895
rect 8527 32861 8536 32895
rect 8484 32852 8536 32861
rect 8576 32895 8628 32904
rect 8576 32861 8585 32895
rect 8585 32861 8619 32895
rect 8619 32861 8628 32895
rect 8576 32852 8628 32861
rect 10140 32852 10192 32904
rect 11152 32852 11204 32904
rect 12256 32852 12308 32904
rect 12072 32784 12124 32836
rect 7012 32716 7064 32768
rect 7932 32716 7984 32768
rect 9404 32716 9456 32768
rect 10324 32759 10376 32768
rect 10324 32725 10333 32759
rect 10333 32725 10367 32759
rect 10367 32725 10376 32759
rect 10324 32716 10376 32725
rect 11980 32716 12032 32768
rect 13084 32716 13136 32768
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 6828 32512 6880 32564
rect 8484 32512 8536 32564
rect 9680 32512 9732 32564
rect 10508 32555 10560 32564
rect 5816 32444 5868 32496
rect 8668 32487 8720 32496
rect 8668 32453 8677 32487
rect 8677 32453 8711 32487
rect 8711 32453 8720 32487
rect 8668 32444 8720 32453
rect 7380 32376 7432 32428
rect 7840 32376 7892 32428
rect 3976 32351 4028 32360
rect 3976 32317 3985 32351
rect 3985 32317 4019 32351
rect 4019 32317 4028 32351
rect 3976 32308 4028 32317
rect 6920 32308 6972 32360
rect 9404 32419 9456 32428
rect 9404 32385 9413 32419
rect 9413 32385 9447 32419
rect 9447 32385 9456 32419
rect 9404 32376 9456 32385
rect 9496 32376 9548 32428
rect 10508 32521 10517 32555
rect 10517 32521 10551 32555
rect 10551 32521 10560 32555
rect 10508 32512 10560 32521
rect 13544 32555 13596 32564
rect 13544 32521 13553 32555
rect 13553 32521 13587 32555
rect 13587 32521 13596 32555
rect 13544 32512 13596 32521
rect 10784 32444 10836 32496
rect 13084 32419 13136 32428
rect 13084 32385 13093 32419
rect 13093 32385 13127 32419
rect 13127 32385 13136 32419
rect 13084 32376 13136 32385
rect 9312 32308 9364 32360
rect 4896 32240 4948 32292
rect 7380 32240 7432 32292
rect 8484 32240 8536 32292
rect 8760 32240 8812 32292
rect 1768 32172 1820 32224
rect 5356 32215 5408 32224
rect 5356 32181 5365 32215
rect 5365 32181 5399 32215
rect 5399 32181 5408 32215
rect 5356 32172 5408 32181
rect 6828 32215 6880 32224
rect 6828 32181 6837 32215
rect 6837 32181 6871 32215
rect 6871 32181 6880 32215
rect 6828 32172 6880 32181
rect 7840 32215 7892 32224
rect 7840 32181 7849 32215
rect 7849 32181 7883 32215
rect 7883 32181 7892 32215
rect 7840 32172 7892 32181
rect 8944 32172 8996 32224
rect 10048 32172 10100 32224
rect 11336 32172 11388 32224
rect 12072 32240 12124 32292
rect 12532 32240 12584 32292
rect 12440 32215 12492 32224
rect 12440 32181 12449 32215
rect 12449 32181 12483 32215
rect 12483 32181 12492 32215
rect 12440 32172 12492 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 5908 31968 5960 32020
rect 8392 31968 8444 32020
rect 10784 32011 10836 32020
rect 10784 31977 10793 32011
rect 10793 31977 10827 32011
rect 10827 31977 10836 32011
rect 10784 31968 10836 31977
rect 11152 32011 11204 32020
rect 11152 31977 11161 32011
rect 11161 31977 11195 32011
rect 11195 31977 11204 32011
rect 11152 31968 11204 31977
rect 1676 31943 1728 31952
rect 1676 31909 1685 31943
rect 1685 31909 1719 31943
rect 1719 31909 1728 31943
rect 1676 31900 1728 31909
rect 5080 31900 5132 31952
rect 5356 31900 5408 31952
rect 5448 31900 5500 31952
rect 6828 31900 6880 31952
rect 8944 31943 8996 31952
rect 8944 31909 8953 31943
rect 8953 31909 8987 31943
rect 8987 31909 8996 31943
rect 8944 31900 8996 31909
rect 10140 31900 10192 31952
rect 3976 31832 4028 31884
rect 6920 31875 6972 31884
rect 6920 31841 6929 31875
rect 6929 31841 6963 31875
rect 6963 31841 6972 31875
rect 6920 31832 6972 31841
rect 7012 31832 7064 31884
rect 10048 31875 10100 31884
rect 10048 31841 10057 31875
rect 10057 31841 10091 31875
rect 10091 31841 10100 31875
rect 10048 31832 10100 31841
rect 10876 31832 10928 31884
rect 11428 31875 11480 31884
rect 11428 31841 11437 31875
rect 11437 31841 11471 31875
rect 11471 31841 11480 31875
rect 11428 31832 11480 31841
rect 12256 31832 12308 31884
rect 1676 31764 1728 31816
rect 7380 31807 7432 31816
rect 7380 31773 7389 31807
rect 7389 31773 7423 31807
rect 7423 31773 7432 31807
rect 7380 31764 7432 31773
rect 10140 31807 10192 31816
rect 7840 31696 7892 31748
rect 10140 31773 10149 31807
rect 10149 31773 10183 31807
rect 10183 31773 10192 31807
rect 10140 31764 10192 31773
rect 8208 31696 8260 31748
rect 9496 31696 9548 31748
rect 14004 31696 14056 31748
rect 14924 31696 14976 31748
rect 8668 31628 8720 31680
rect 12808 31671 12860 31680
rect 12808 31637 12817 31671
rect 12817 31637 12851 31671
rect 12851 31637 12860 31671
rect 12808 31628 12860 31637
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 4252 31424 4304 31476
rect 5080 31467 5132 31476
rect 5080 31433 5089 31467
rect 5089 31433 5123 31467
rect 5123 31433 5132 31467
rect 5080 31424 5132 31433
rect 6828 31424 6880 31476
rect 7012 31467 7064 31476
rect 7012 31433 7021 31467
rect 7021 31433 7055 31467
rect 7055 31433 7064 31467
rect 7012 31424 7064 31433
rect 7472 31467 7524 31476
rect 7472 31433 7481 31467
rect 7481 31433 7515 31467
rect 7515 31433 7524 31467
rect 7472 31424 7524 31433
rect 8208 31424 8260 31476
rect 8392 31424 8444 31476
rect 1676 31399 1728 31408
rect 1676 31365 1685 31399
rect 1685 31365 1719 31399
rect 1719 31365 1728 31399
rect 1676 31356 1728 31365
rect 7656 31288 7708 31340
rect 8116 31331 8168 31340
rect 8116 31297 8125 31331
rect 8125 31297 8159 31331
rect 8159 31297 8168 31331
rect 8116 31288 8168 31297
rect 10048 31424 10100 31476
rect 11152 31424 11204 31476
rect 12164 31424 12216 31476
rect 12256 31424 12308 31476
rect 10324 31288 10376 31340
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 10968 31331 11020 31340
rect 10968 31297 10977 31331
rect 10977 31297 11011 31331
rect 11011 31297 11020 31331
rect 10968 31288 11020 31297
rect 7932 31263 7984 31272
rect 7932 31229 7941 31263
rect 7941 31229 7975 31263
rect 7975 31229 7984 31263
rect 7932 31220 7984 31229
rect 9772 31220 9824 31272
rect 10048 31220 10100 31272
rect 6644 31152 6696 31204
rect 5448 31127 5500 31136
rect 5448 31093 5457 31127
rect 5457 31093 5491 31127
rect 5491 31093 5500 31127
rect 5448 31084 5500 31093
rect 7564 31127 7616 31136
rect 7564 31093 7573 31127
rect 7573 31093 7607 31127
rect 7607 31093 7616 31127
rect 7564 31084 7616 31093
rect 8576 31084 8628 31136
rect 9496 31084 9548 31136
rect 9772 31084 9824 31136
rect 10140 31084 10192 31136
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 10784 31127 10836 31136
rect 10784 31093 10793 31127
rect 10793 31093 10827 31127
rect 10827 31093 10836 31127
rect 10784 31084 10836 31093
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 8484 30923 8536 30932
rect 8484 30889 8493 30923
rect 8493 30889 8527 30923
rect 8527 30889 8536 30923
rect 8484 30880 8536 30889
rect 10140 30880 10192 30932
rect 10508 30880 10560 30932
rect 10876 30880 10928 30932
rect 7656 30855 7708 30864
rect 7656 30821 7665 30855
rect 7665 30821 7699 30855
rect 7699 30821 7708 30855
rect 7656 30812 7708 30821
rect 10968 30812 11020 30864
rect 11796 30855 11848 30864
rect 11796 30821 11805 30855
rect 11805 30821 11839 30855
rect 11839 30821 11848 30855
rect 11796 30812 11848 30821
rect 11888 30812 11940 30864
rect 12440 30812 12492 30864
rect 4528 30787 4580 30796
rect 4528 30753 4537 30787
rect 4537 30753 4571 30787
rect 4571 30753 4580 30787
rect 4528 30744 4580 30753
rect 7104 30744 7156 30796
rect 8208 30744 8260 30796
rect 9864 30744 9916 30796
rect 11980 30744 12032 30796
rect 4620 30719 4672 30728
rect 4620 30685 4629 30719
rect 4629 30685 4663 30719
rect 4663 30685 4672 30719
rect 4620 30676 4672 30685
rect 4896 30676 4948 30728
rect 7012 30719 7064 30728
rect 7012 30685 7021 30719
rect 7021 30685 7055 30719
rect 7055 30685 7064 30719
rect 7012 30676 7064 30685
rect 8576 30719 8628 30728
rect 8576 30685 8585 30719
rect 8585 30685 8619 30719
rect 8619 30685 8628 30719
rect 8576 30676 8628 30685
rect 10232 30719 10284 30728
rect 10232 30685 10241 30719
rect 10241 30685 10275 30719
rect 10275 30685 10284 30719
rect 10232 30676 10284 30685
rect 11152 30676 11204 30728
rect 6644 30608 6696 30660
rect 9680 30651 9732 30660
rect 9680 30617 9689 30651
rect 9689 30617 9723 30651
rect 9723 30617 9732 30651
rect 9680 30608 9732 30617
rect 10784 30608 10836 30660
rect 4160 30583 4212 30592
rect 4160 30549 4169 30583
rect 4169 30549 4203 30583
rect 4203 30549 4212 30583
rect 4160 30540 4212 30549
rect 6000 30583 6052 30592
rect 6000 30549 6009 30583
rect 6009 30549 6043 30583
rect 6043 30549 6052 30583
rect 6000 30540 6052 30549
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 2228 30311 2280 30320
rect 2228 30277 2237 30311
rect 2237 30277 2271 30311
rect 2271 30277 2280 30311
rect 2228 30268 2280 30277
rect 1584 30243 1636 30252
rect 1584 30209 1593 30243
rect 1593 30209 1627 30243
rect 1627 30209 1636 30243
rect 1584 30200 1636 30209
rect 7012 30336 7064 30388
rect 5448 30268 5500 30320
rect 9496 30336 9548 30388
rect 10232 30336 10284 30388
rect 10784 30379 10836 30388
rect 10784 30345 10793 30379
rect 10793 30345 10827 30379
rect 10827 30345 10836 30379
rect 10784 30336 10836 30345
rect 11152 30336 11204 30388
rect 11796 30379 11848 30388
rect 11796 30345 11805 30379
rect 11805 30345 11839 30379
rect 11839 30345 11848 30379
rect 11796 30336 11848 30345
rect 11980 30336 12032 30388
rect 6184 30200 6236 30252
rect 6000 30132 6052 30184
rect 6644 30132 6696 30184
rect 8668 30268 8720 30320
rect 8300 30132 8352 30184
rect 4804 30064 4856 30116
rect 8576 30064 8628 30116
rect 9680 30064 9732 30116
rect 9864 30064 9916 30116
rect 4896 30039 4948 30048
rect 4896 30005 4905 30039
rect 4905 30005 4939 30039
rect 4939 30005 4948 30039
rect 4896 29996 4948 30005
rect 7104 30039 7156 30048
rect 7104 30005 7113 30039
rect 7113 30005 7147 30039
rect 7147 30005 7156 30039
rect 7104 29996 7156 30005
rect 7564 30039 7616 30048
rect 7564 30005 7573 30039
rect 7573 30005 7607 30039
rect 7607 30005 7616 30039
rect 7564 29996 7616 30005
rect 8208 29996 8260 30048
rect 10140 29996 10192 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 4620 29792 4672 29844
rect 7104 29835 7156 29844
rect 7104 29801 7113 29835
rect 7113 29801 7147 29835
rect 7147 29801 7156 29835
rect 7104 29792 7156 29801
rect 7288 29792 7340 29844
rect 7656 29792 7708 29844
rect 8300 29792 8352 29844
rect 10232 29792 10284 29844
rect 2780 29767 2832 29776
rect 2780 29733 2789 29767
rect 2789 29733 2823 29767
rect 2823 29733 2832 29767
rect 2780 29724 2832 29733
rect 4068 29724 4120 29776
rect 7012 29724 7064 29776
rect 9864 29724 9916 29776
rect 2964 29656 3016 29708
rect 4160 29656 4212 29708
rect 5724 29656 5776 29708
rect 6000 29699 6052 29708
rect 6000 29665 6009 29699
rect 6009 29665 6043 29699
rect 6043 29665 6052 29699
rect 6000 29656 6052 29665
rect 6276 29656 6328 29708
rect 8484 29656 8536 29708
rect 9496 29656 9548 29708
rect 10784 29656 10836 29708
rect 2872 29631 2924 29640
rect 2872 29597 2881 29631
rect 2881 29597 2915 29631
rect 2915 29597 2924 29631
rect 2872 29588 2924 29597
rect 3056 29631 3108 29640
rect 3056 29597 3065 29631
rect 3065 29597 3099 29631
rect 3099 29597 3108 29631
rect 3056 29588 3108 29597
rect 4252 29588 4304 29640
rect 4620 29588 4672 29640
rect 4804 29588 4856 29640
rect 5356 29588 5408 29640
rect 7656 29631 7708 29640
rect 7656 29597 7665 29631
rect 7665 29597 7699 29631
rect 7699 29597 7708 29631
rect 7656 29588 7708 29597
rect 7840 29631 7892 29640
rect 7840 29597 7849 29631
rect 7849 29597 7883 29631
rect 7883 29597 7892 29631
rect 7840 29588 7892 29597
rect 1400 29452 1452 29504
rect 3516 29495 3568 29504
rect 3516 29461 3525 29495
rect 3525 29461 3559 29495
rect 3559 29461 3568 29495
rect 3516 29452 3568 29461
rect 5172 29495 5224 29504
rect 5172 29461 5181 29495
rect 5181 29461 5215 29495
rect 5215 29461 5224 29495
rect 5172 29452 5224 29461
rect 7196 29495 7248 29504
rect 7196 29461 7205 29495
rect 7205 29461 7239 29495
rect 7239 29461 7248 29495
rect 7196 29452 7248 29461
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 2872 29248 2924 29300
rect 4160 29248 4212 29300
rect 4528 29248 4580 29300
rect 7656 29248 7708 29300
rect 8668 29248 8720 29300
rect 3056 29180 3108 29232
rect 4252 29180 4304 29232
rect 5264 29180 5316 29232
rect 6276 29223 6328 29232
rect 6276 29189 6285 29223
rect 6285 29189 6319 29223
rect 6319 29189 6328 29223
rect 6276 29180 6328 29189
rect 9220 29180 9272 29232
rect 9588 29180 9640 29232
rect 4896 29112 4948 29164
rect 5356 29155 5408 29164
rect 5356 29121 5365 29155
rect 5365 29121 5399 29155
rect 5399 29121 5408 29155
rect 5356 29112 5408 29121
rect 5540 29112 5592 29164
rect 1400 29087 1452 29096
rect 1400 29053 1409 29087
rect 1409 29053 1443 29087
rect 1443 29053 1452 29087
rect 1400 29044 1452 29053
rect 3608 29087 3660 29096
rect 3608 29053 3617 29087
rect 3617 29053 3651 29087
rect 3651 29053 3660 29087
rect 3608 29044 3660 29053
rect 4804 29044 4856 29096
rect 5172 29087 5224 29096
rect 5172 29053 5181 29087
rect 5181 29053 5215 29087
rect 5215 29053 5224 29087
rect 5172 29044 5224 29053
rect 1492 28976 1544 29028
rect 6092 29044 6144 29096
rect 6000 28976 6052 29028
rect 7196 29112 7248 29164
rect 7472 29155 7524 29164
rect 7472 29121 7481 29155
rect 7481 29121 7515 29155
rect 7515 29121 7524 29155
rect 7472 29112 7524 29121
rect 9864 29112 9916 29164
rect 9312 29044 9364 29096
rect 9588 29044 9640 29096
rect 10416 29044 10468 29096
rect 7748 28976 7800 29028
rect 9864 28976 9916 29028
rect 3424 28908 3476 28960
rect 6828 28951 6880 28960
rect 6828 28917 6837 28951
rect 6837 28917 6871 28951
rect 6871 28917 6880 28951
rect 6828 28908 6880 28917
rect 9680 28951 9732 28960
rect 9680 28917 9689 28951
rect 9689 28917 9723 28951
rect 9723 28917 9732 28951
rect 9680 28908 9732 28917
rect 10784 28951 10836 28960
rect 10784 28917 10793 28951
rect 10793 28917 10827 28951
rect 10827 28917 10836 28951
rect 10784 28908 10836 28917
rect 11428 28908 11480 28960
rect 12900 28908 12952 28960
rect 14004 28908 14056 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 2780 28747 2832 28756
rect 2780 28713 2789 28747
rect 2789 28713 2823 28747
rect 2823 28713 2832 28747
rect 2780 28704 2832 28713
rect 4620 28704 4672 28756
rect 5172 28704 5224 28756
rect 5908 28704 5960 28756
rect 7196 28704 7248 28756
rect 7472 28704 7524 28756
rect 7840 28704 7892 28756
rect 9864 28747 9916 28756
rect 9864 28713 9873 28747
rect 9873 28713 9907 28747
rect 9907 28713 9916 28747
rect 9864 28704 9916 28713
rect 2872 28636 2924 28688
rect 5448 28636 5500 28688
rect 6828 28636 6880 28688
rect 7288 28679 7340 28688
rect 7288 28645 7297 28679
rect 7297 28645 7331 28679
rect 7331 28645 7340 28679
rect 7288 28636 7340 28645
rect 11060 28636 11112 28688
rect 1584 28568 1636 28620
rect 8852 28568 8904 28620
rect 10600 28611 10652 28620
rect 10600 28577 10609 28611
rect 10609 28577 10643 28611
rect 10643 28577 10652 28611
rect 10600 28568 10652 28577
rect 5816 28500 5868 28552
rect 3148 28432 3200 28484
rect 8576 28432 8628 28484
rect 11336 28568 11388 28620
rect 3424 28364 3476 28416
rect 5172 28407 5224 28416
rect 5172 28373 5181 28407
rect 5181 28373 5215 28407
rect 5215 28373 5224 28407
rect 5172 28364 5224 28373
rect 5356 28364 5408 28416
rect 5632 28364 5684 28416
rect 8300 28407 8352 28416
rect 8300 28373 8309 28407
rect 8309 28373 8343 28407
rect 8343 28373 8352 28407
rect 8300 28364 8352 28373
rect 8852 28407 8904 28416
rect 8852 28373 8861 28407
rect 8861 28373 8895 28407
rect 8895 28373 8904 28407
rect 8852 28364 8904 28373
rect 11980 28364 12032 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 5448 28203 5500 28212
rect 5448 28169 5457 28203
rect 5457 28169 5491 28203
rect 5491 28169 5500 28203
rect 5448 28160 5500 28169
rect 5816 28203 5868 28212
rect 5816 28169 5825 28203
rect 5825 28169 5859 28203
rect 5859 28169 5868 28203
rect 5816 28160 5868 28169
rect 5908 28160 5960 28212
rect 7564 28160 7616 28212
rect 7840 28160 7892 28212
rect 9864 28160 9916 28212
rect 11060 28160 11112 28212
rect 11428 28160 11480 28212
rect 2412 28067 2464 28076
rect 1584 27956 1636 28008
rect 2412 28033 2421 28067
rect 2421 28033 2455 28067
rect 2455 28033 2464 28067
rect 2412 28024 2464 28033
rect 8484 28024 8536 28076
rect 8576 27999 8628 28008
rect 8576 27965 8585 27999
rect 8585 27965 8619 27999
rect 8619 27965 8628 27999
rect 8576 27956 8628 27965
rect 2688 27820 2740 27872
rect 7012 27863 7064 27872
rect 7012 27829 7021 27863
rect 7021 27829 7055 27863
rect 7055 27829 7064 27863
rect 7012 27820 7064 27829
rect 7380 27863 7432 27872
rect 7380 27829 7389 27863
rect 7389 27829 7423 27863
rect 7423 27829 7432 27863
rect 7380 27820 7432 27829
rect 8116 27863 8168 27872
rect 8116 27829 8125 27863
rect 8125 27829 8159 27863
rect 8159 27829 8168 27863
rect 8116 27820 8168 27829
rect 10600 27863 10652 27872
rect 10600 27829 10609 27863
rect 10609 27829 10643 27863
rect 10643 27829 10652 27863
rect 10600 27820 10652 27829
rect 10968 27820 11020 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 3424 27616 3476 27668
rect 1676 27591 1728 27600
rect 1676 27557 1685 27591
rect 1685 27557 1719 27591
rect 1719 27557 1728 27591
rect 1676 27548 1728 27557
rect 6184 27548 6236 27600
rect 7380 27616 7432 27668
rect 8484 27659 8536 27668
rect 8484 27625 8493 27659
rect 8493 27625 8527 27659
rect 8527 27625 8536 27659
rect 8484 27616 8536 27625
rect 9680 27659 9732 27668
rect 9680 27625 9689 27659
rect 9689 27625 9723 27659
rect 9723 27625 9732 27659
rect 9680 27616 9732 27625
rect 11428 27616 11480 27668
rect 11980 27591 12032 27600
rect 11980 27557 12014 27591
rect 12014 27557 12032 27591
rect 11980 27548 12032 27557
rect 1400 27523 1452 27532
rect 1400 27489 1409 27523
rect 1409 27489 1443 27523
rect 1443 27489 1452 27523
rect 1400 27480 1452 27489
rect 3516 27480 3568 27532
rect 5540 27480 5592 27532
rect 4528 27455 4580 27464
rect 4528 27421 4537 27455
rect 4537 27421 4571 27455
rect 4571 27421 4580 27455
rect 4528 27412 4580 27421
rect 5172 27412 5224 27464
rect 5448 27412 5500 27464
rect 6736 27523 6788 27532
rect 6736 27489 6745 27523
rect 6745 27489 6779 27523
rect 6779 27489 6788 27523
rect 6736 27480 6788 27489
rect 7932 27480 7984 27532
rect 8484 27412 8536 27464
rect 8760 27412 8812 27464
rect 6644 27344 6696 27396
rect 8760 27276 8812 27328
rect 11428 27523 11480 27532
rect 11428 27489 11437 27523
rect 11437 27489 11471 27523
rect 11471 27489 11480 27523
rect 11428 27480 11480 27489
rect 9496 27412 9548 27464
rect 9680 27412 9732 27464
rect 9404 27319 9456 27328
rect 9404 27285 9413 27319
rect 9413 27285 9447 27319
rect 9447 27285 9456 27319
rect 10232 27455 10284 27464
rect 10232 27421 10241 27455
rect 10241 27421 10275 27455
rect 10275 27421 10284 27455
rect 10232 27412 10284 27421
rect 9404 27276 9456 27285
rect 11152 27276 11204 27328
rect 13084 27319 13136 27328
rect 13084 27285 13093 27319
rect 13093 27285 13127 27319
rect 13127 27285 13136 27319
rect 13084 27276 13136 27285
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 1400 27072 1452 27124
rect 3516 27115 3568 27124
rect 3516 27081 3525 27115
rect 3525 27081 3559 27115
rect 3559 27081 3568 27115
rect 3516 27072 3568 27081
rect 4528 27072 4580 27124
rect 6736 27072 6788 27124
rect 7196 27072 7248 27124
rect 8576 27072 8628 27124
rect 10416 27115 10468 27124
rect 3976 26936 4028 26988
rect 8300 27004 8352 27056
rect 7472 26936 7524 26988
rect 10416 27081 10425 27115
rect 10425 27081 10459 27115
rect 10459 27081 10468 27115
rect 10416 27072 10468 27081
rect 11428 27072 11480 27124
rect 9496 26979 9548 26988
rect 9496 26945 9505 26979
rect 9505 26945 9539 26979
rect 9539 26945 9548 26979
rect 9496 26936 9548 26945
rect 11060 26936 11112 26988
rect 11980 27004 12032 27056
rect 12532 26936 12584 26988
rect 13360 26936 13412 26988
rect 10416 26868 10468 26920
rect 12808 26868 12860 26920
rect 13728 26868 13780 26920
rect 4068 26800 4120 26852
rect 4988 26800 5040 26852
rect 7288 26843 7340 26852
rect 7288 26809 7297 26843
rect 7297 26809 7331 26843
rect 7331 26809 7340 26843
rect 7288 26800 7340 26809
rect 4620 26732 4672 26784
rect 5448 26732 5500 26784
rect 6828 26775 6880 26784
rect 6828 26741 6837 26775
rect 6837 26741 6871 26775
rect 6871 26741 6880 26775
rect 6828 26732 6880 26741
rect 7932 26775 7984 26784
rect 7932 26741 7941 26775
rect 7941 26741 7975 26775
rect 7975 26741 7984 26775
rect 7932 26732 7984 26741
rect 8392 26775 8444 26784
rect 8392 26741 8401 26775
rect 8401 26741 8435 26775
rect 8435 26741 8444 26775
rect 8392 26732 8444 26741
rect 9588 26732 9640 26784
rect 9864 26732 9916 26784
rect 10784 26732 10836 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 4528 26528 4580 26580
rect 5816 26528 5868 26580
rect 6184 26528 6236 26580
rect 7472 26528 7524 26580
rect 8760 26528 8812 26580
rect 9312 26528 9364 26580
rect 9496 26528 9548 26580
rect 10232 26528 10284 26580
rect 11336 26528 11388 26580
rect 8208 26392 8260 26444
rect 9680 26392 9732 26444
rect 8300 26324 8352 26376
rect 9588 26324 9640 26376
rect 9956 26324 10008 26376
rect 10140 26324 10192 26376
rect 11060 26367 11112 26376
rect 11060 26333 11069 26367
rect 11069 26333 11103 26367
rect 11103 26333 11112 26367
rect 11060 26324 11112 26333
rect 4068 26188 4120 26240
rect 4528 26188 4580 26240
rect 6736 26188 6788 26240
rect 9496 26188 9548 26240
rect 10968 26188 11020 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 3976 26027 4028 26036
rect 3976 25993 3985 26027
rect 3985 25993 4019 26027
rect 4019 25993 4028 26027
rect 3976 25984 4028 25993
rect 5448 26027 5500 26036
rect 5448 25993 5457 26027
rect 5457 25993 5491 26027
rect 5491 25993 5500 26027
rect 5448 25984 5500 25993
rect 7104 25984 7156 26036
rect 8024 26027 8076 26036
rect 8024 25993 8033 26027
rect 8033 25993 8067 26027
rect 8067 25993 8076 26027
rect 8024 25984 8076 25993
rect 8208 25984 8260 26036
rect 9404 25984 9456 26036
rect 11060 25984 11112 26036
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 10876 25916 10928 25968
rect 7472 25891 7524 25900
rect 4068 25823 4120 25832
rect 4068 25789 4077 25823
rect 4077 25789 4111 25823
rect 4111 25789 4120 25823
rect 4068 25780 4120 25789
rect 7472 25857 7481 25891
rect 7481 25857 7515 25891
rect 7515 25857 7524 25891
rect 7472 25848 7524 25857
rect 5448 25780 5500 25832
rect 6920 25780 6972 25832
rect 8208 25780 8260 25832
rect 10784 25848 10836 25900
rect 11336 25848 11388 25900
rect 9496 25780 9548 25832
rect 10508 25823 10560 25832
rect 10508 25789 10517 25823
rect 10517 25789 10551 25823
rect 10551 25789 10560 25823
rect 10508 25780 10560 25789
rect 10968 25823 11020 25832
rect 10968 25789 10977 25823
rect 10977 25789 11011 25823
rect 11011 25789 11020 25823
rect 10968 25780 11020 25789
rect 7288 25755 7340 25764
rect 7288 25721 7297 25755
rect 7297 25721 7331 25755
rect 7331 25721 7340 25755
rect 7288 25712 7340 25721
rect 9404 25712 9456 25764
rect 2228 25687 2280 25696
rect 2228 25653 2237 25687
rect 2237 25653 2271 25687
rect 2271 25653 2280 25687
rect 2228 25644 2280 25653
rect 6920 25644 6972 25696
rect 9312 25644 9364 25696
rect 9680 25644 9732 25696
rect 9956 25644 10008 25696
rect 10600 25687 10652 25696
rect 10600 25653 10609 25687
rect 10609 25653 10643 25687
rect 10643 25653 10652 25687
rect 10600 25644 10652 25653
rect 12716 25644 12768 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 5448 25483 5500 25492
rect 5448 25449 5457 25483
rect 5457 25449 5491 25483
rect 5491 25449 5500 25483
rect 5448 25440 5500 25449
rect 6644 25440 6696 25492
rect 8668 25440 8720 25492
rect 9220 25483 9272 25492
rect 9220 25449 9229 25483
rect 9229 25449 9263 25483
rect 9263 25449 9272 25483
rect 9220 25440 9272 25449
rect 9588 25440 9640 25492
rect 10140 25440 10192 25492
rect 7472 25372 7524 25424
rect 10508 25372 10560 25424
rect 11152 25372 11204 25424
rect 4068 25347 4120 25356
rect 4068 25313 4077 25347
rect 4077 25313 4111 25347
rect 4111 25313 4120 25347
rect 4068 25304 4120 25313
rect 4160 25304 4212 25356
rect 7012 25304 7064 25356
rect 12716 25347 12768 25356
rect 12716 25313 12725 25347
rect 12725 25313 12759 25347
rect 12759 25313 12768 25347
rect 12716 25304 12768 25313
rect 13176 25304 13228 25356
rect 13912 25304 13964 25356
rect 8208 25236 8260 25288
rect 8392 25236 8444 25288
rect 10048 25168 10100 25220
rect 10508 25168 10560 25220
rect 10968 25279 11020 25288
rect 10968 25245 10977 25279
rect 10977 25245 11011 25279
rect 11011 25245 11020 25279
rect 10968 25236 11020 25245
rect 11336 25168 11388 25220
rect 13084 25168 13136 25220
rect 6736 25100 6788 25152
rect 8392 25100 8444 25152
rect 9312 25100 9364 25152
rect 10416 25143 10468 25152
rect 10416 25109 10425 25143
rect 10425 25109 10459 25143
rect 10459 25109 10468 25143
rect 10416 25100 10468 25109
rect 12348 25143 12400 25152
rect 12348 25109 12357 25143
rect 12357 25109 12391 25143
rect 12391 25109 12400 25143
rect 12348 25100 12400 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 4068 24896 4120 24948
rect 5172 24939 5224 24948
rect 5172 24905 5181 24939
rect 5181 24905 5215 24939
rect 5215 24905 5224 24939
rect 5172 24896 5224 24905
rect 6184 24939 6236 24948
rect 6184 24905 6193 24939
rect 6193 24905 6227 24939
rect 6227 24905 6236 24939
rect 6184 24896 6236 24905
rect 7012 24896 7064 24948
rect 9312 24896 9364 24948
rect 10048 24896 10100 24948
rect 12716 24896 12768 24948
rect 12072 24828 12124 24880
rect 5632 24803 5684 24812
rect 5632 24769 5641 24803
rect 5641 24769 5675 24803
rect 5675 24769 5684 24803
rect 5632 24760 5684 24769
rect 6920 24760 6972 24812
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 8300 24803 8352 24812
rect 8300 24769 8309 24803
rect 8309 24769 8343 24803
rect 8343 24769 8352 24803
rect 8300 24760 8352 24769
rect 8392 24760 8444 24812
rect 9588 24760 9640 24812
rect 11336 24803 11388 24812
rect 11336 24769 11345 24803
rect 11345 24769 11379 24803
rect 11379 24769 11388 24803
rect 11336 24760 11388 24769
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 8944 24735 8996 24744
rect 8944 24701 8953 24735
rect 8953 24701 8987 24735
rect 8987 24701 8996 24735
rect 8944 24692 8996 24701
rect 6920 24624 6972 24676
rect 10416 24624 10468 24676
rect 11336 24624 11388 24676
rect 12256 24624 12308 24676
rect 13176 24624 13228 24676
rect 4160 24599 4212 24608
rect 4160 24565 4169 24599
rect 4169 24565 4203 24599
rect 4203 24565 4212 24599
rect 4160 24556 4212 24565
rect 9312 24556 9364 24608
rect 10324 24556 10376 24608
rect 10692 24599 10744 24608
rect 10692 24565 10701 24599
rect 10701 24565 10735 24599
rect 10735 24565 10744 24599
rect 10692 24556 10744 24565
rect 12716 24556 12768 24608
rect 13728 24556 13780 24608
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 5632 24352 5684 24404
rect 6920 24352 6972 24404
rect 8208 24352 8260 24404
rect 9588 24352 9640 24404
rect 10416 24352 10468 24404
rect 10600 24352 10652 24404
rect 11428 24395 11480 24404
rect 11428 24361 11437 24395
rect 11437 24361 11471 24395
rect 11471 24361 11480 24395
rect 11428 24352 11480 24361
rect 6184 24284 6236 24336
rect 7472 24284 7524 24336
rect 4252 24216 4304 24268
rect 6644 24216 6696 24268
rect 10692 24216 10744 24268
rect 11060 24216 11112 24268
rect 5632 24191 5684 24200
rect 5632 24157 5641 24191
rect 5641 24157 5675 24191
rect 5675 24157 5684 24191
rect 5632 24148 5684 24157
rect 10784 24148 10836 24200
rect 10876 24148 10928 24200
rect 11152 24148 11204 24200
rect 7012 24123 7064 24132
rect 7012 24089 7021 24123
rect 7021 24089 7055 24123
rect 7055 24089 7064 24123
rect 7012 24080 7064 24089
rect 4528 24012 4580 24064
rect 8208 24012 8260 24064
rect 9312 24012 9364 24064
rect 10048 24055 10100 24064
rect 10048 24021 10057 24055
rect 10057 24021 10091 24055
rect 10091 24021 10100 24055
rect 10048 24012 10100 24021
rect 10140 24012 10192 24064
rect 12992 24055 13044 24064
rect 12992 24021 13001 24055
rect 13001 24021 13035 24055
rect 13035 24021 13044 24055
rect 12992 24012 13044 24021
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 6184 23808 6236 23860
rect 8668 23851 8720 23860
rect 8668 23817 8677 23851
rect 8677 23817 8711 23851
rect 8711 23817 8720 23851
rect 8668 23808 8720 23817
rect 10784 23851 10836 23860
rect 10784 23817 10793 23851
rect 10793 23817 10827 23851
rect 10827 23817 10836 23851
rect 10784 23808 10836 23817
rect 11060 23851 11112 23860
rect 11060 23817 11069 23851
rect 11069 23817 11103 23851
rect 11103 23817 11112 23851
rect 11060 23808 11112 23817
rect 11428 23808 11480 23860
rect 12992 23715 13044 23724
rect 8760 23647 8812 23656
rect 8760 23613 8769 23647
rect 8769 23613 8803 23647
rect 8803 23613 8812 23647
rect 8760 23604 8812 23613
rect 9312 23604 9364 23656
rect 10784 23604 10836 23656
rect 12164 23647 12216 23656
rect 12164 23613 12173 23647
rect 12173 23613 12207 23647
rect 12207 23613 12216 23647
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 12164 23604 12216 23613
rect 12348 23604 12400 23656
rect 12624 23604 12676 23656
rect 12716 23604 12768 23656
rect 5632 23468 5684 23520
rect 6736 23468 6788 23520
rect 9496 23468 9548 23520
rect 10232 23468 10284 23520
rect 12440 23511 12492 23520
rect 12440 23477 12449 23511
rect 12449 23477 12483 23511
rect 12483 23477 12492 23511
rect 12440 23468 12492 23477
rect 12624 23468 12676 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 4436 23264 4488 23316
rect 4896 23264 4948 23316
rect 9312 23307 9364 23316
rect 9312 23273 9321 23307
rect 9321 23273 9355 23307
rect 9355 23273 9364 23307
rect 9312 23264 9364 23273
rect 9864 23264 9916 23316
rect 10048 23264 10100 23316
rect 10876 23264 10928 23316
rect 11152 23264 11204 23316
rect 12072 23264 12124 23316
rect 12348 23264 12400 23316
rect 10600 23196 10652 23248
rect 9772 23128 9824 23180
rect 10048 23128 10100 23180
rect 11336 23196 11388 23248
rect 12072 23171 12124 23180
rect 12072 23137 12081 23171
rect 12081 23137 12115 23171
rect 12115 23137 12124 23171
rect 12072 23128 12124 23137
rect 12164 23128 12216 23180
rect 5356 23060 5408 23112
rect 10600 23060 10652 23112
rect 10508 23035 10560 23044
rect 10508 23001 10517 23035
rect 10517 23001 10551 23035
rect 10551 23001 10560 23035
rect 10508 22992 10560 23001
rect 2504 22924 2556 22976
rect 2780 22924 2832 22976
rect 4804 22967 4856 22976
rect 4804 22933 4813 22967
rect 4813 22933 4847 22967
rect 4847 22933 4856 22967
rect 4804 22924 4856 22933
rect 5816 22967 5868 22976
rect 5816 22933 5825 22967
rect 5825 22933 5859 22967
rect 5859 22933 5868 22967
rect 5816 22924 5868 22933
rect 7656 22967 7708 22976
rect 7656 22933 7665 22967
rect 7665 22933 7699 22967
rect 7699 22933 7708 22967
rect 7656 22924 7708 22933
rect 8760 22924 8812 22976
rect 9312 22924 9364 22976
rect 12348 22924 12400 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 4896 22763 4948 22772
rect 4896 22729 4905 22763
rect 4905 22729 4939 22763
rect 4939 22729 4948 22763
rect 4896 22720 4948 22729
rect 5356 22720 5408 22772
rect 7196 22720 7248 22772
rect 7380 22720 7432 22772
rect 8300 22720 8352 22772
rect 4620 22652 4672 22704
rect 7932 22652 7984 22704
rect 2504 22627 2556 22636
rect 2504 22593 2513 22627
rect 2513 22593 2547 22627
rect 2547 22593 2556 22627
rect 2504 22584 2556 22593
rect 4252 22584 4304 22636
rect 5816 22584 5868 22636
rect 6920 22584 6972 22636
rect 7656 22584 7708 22636
rect 8300 22584 8352 22636
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 9404 22720 9456 22772
rect 10600 22763 10652 22772
rect 10600 22729 10609 22763
rect 10609 22729 10643 22763
rect 10643 22729 10652 22763
rect 10600 22720 10652 22729
rect 10876 22763 10928 22772
rect 10876 22729 10885 22763
rect 10885 22729 10919 22763
rect 10919 22729 10928 22763
rect 10876 22720 10928 22729
rect 11336 22763 11388 22772
rect 11336 22729 11345 22763
rect 11345 22729 11379 22763
rect 11379 22729 11388 22763
rect 11336 22720 11388 22729
rect 11428 22720 11480 22772
rect 12164 22763 12216 22772
rect 12164 22729 12173 22763
rect 12173 22729 12207 22763
rect 12207 22729 12216 22763
rect 12164 22720 12216 22729
rect 9864 22627 9916 22636
rect 9864 22593 9873 22627
rect 9873 22593 9907 22627
rect 9907 22593 9916 22627
rect 9864 22584 9916 22593
rect 10324 22516 10376 22568
rect 11428 22516 11480 22568
rect 4068 22448 4120 22500
rect 2964 22380 3016 22432
rect 4160 22380 4212 22432
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 5908 22380 5960 22432
rect 7932 22423 7984 22432
rect 7932 22389 7941 22423
rect 7941 22389 7975 22423
rect 7975 22389 7984 22423
rect 7932 22380 7984 22389
rect 9496 22380 9548 22432
rect 12072 22380 12124 22432
rect 12624 22423 12676 22432
rect 12624 22389 12633 22423
rect 12633 22389 12667 22423
rect 12667 22389 12676 22423
rect 12624 22380 12676 22389
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 8300 22176 8352 22228
rect 9680 22219 9732 22228
rect 9680 22185 9689 22219
rect 9689 22185 9723 22219
rect 9723 22185 9732 22219
rect 9680 22176 9732 22185
rect 9772 22176 9824 22228
rect 10048 22176 10100 22228
rect 4160 22108 4212 22160
rect 8208 22108 8260 22160
rect 3240 22040 3292 22092
rect 2964 22015 3016 22024
rect 2964 21981 2973 22015
rect 2973 21981 3007 22015
rect 3007 21981 3016 22015
rect 2964 21972 3016 21981
rect 6276 22040 6328 22092
rect 6736 22040 6788 22092
rect 7380 22083 7432 22092
rect 7380 22049 7414 22083
rect 7414 22049 7432 22083
rect 7380 22040 7432 22049
rect 9956 22108 10008 22160
rect 12900 22176 12952 22228
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 12348 22083 12400 22092
rect 12348 22049 12382 22083
rect 12382 22049 12400 22083
rect 12348 22040 12400 22049
rect 3332 21904 3384 21956
rect 2136 21836 2188 21888
rect 2780 21836 2832 21888
rect 5632 21972 5684 22024
rect 8300 21972 8352 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 11520 21972 11572 22024
rect 5448 21879 5500 21888
rect 5448 21845 5457 21879
rect 5457 21845 5491 21879
rect 5491 21845 5500 21879
rect 5448 21836 5500 21845
rect 5908 21836 5960 21888
rect 6736 21836 6788 21888
rect 8668 21836 8720 21888
rect 9496 21836 9548 21888
rect 10600 21836 10652 21888
rect 13452 21879 13504 21888
rect 13452 21845 13461 21879
rect 13461 21845 13495 21879
rect 13495 21845 13504 21879
rect 13452 21836 13504 21845
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 5172 21632 5224 21684
rect 6276 21675 6328 21684
rect 6276 21641 6285 21675
rect 6285 21641 6319 21675
rect 6319 21641 6328 21675
rect 6276 21632 6328 21641
rect 7656 21632 7708 21684
rect 9956 21632 10008 21684
rect 10232 21632 10284 21684
rect 12348 21632 12400 21684
rect 12624 21675 12676 21684
rect 12624 21641 12633 21675
rect 12633 21641 12667 21675
rect 12667 21641 12676 21675
rect 12624 21632 12676 21641
rect 13636 21675 13688 21684
rect 13636 21641 13645 21675
rect 13645 21641 13679 21675
rect 13679 21641 13688 21675
rect 13636 21632 13688 21641
rect 3240 21564 3292 21616
rect 2872 21428 2924 21480
rect 4528 21539 4580 21548
rect 4528 21505 4537 21539
rect 4537 21505 4571 21539
rect 4571 21505 4580 21539
rect 4528 21496 4580 21505
rect 5448 21496 5500 21548
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 4252 21428 4304 21480
rect 8208 21428 8260 21480
rect 12164 21428 12216 21480
rect 13452 21471 13504 21480
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 2412 21335 2464 21344
rect 2412 21301 2421 21335
rect 2421 21301 2455 21335
rect 2455 21301 2464 21335
rect 2412 21292 2464 21301
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 4160 21292 4212 21344
rect 4988 21292 5040 21344
rect 5356 21292 5408 21344
rect 7932 21292 7984 21344
rect 8116 21292 8168 21344
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 11520 21292 11572 21344
rect 12624 21292 12676 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 2964 21131 3016 21140
rect 2964 21097 2973 21131
rect 2973 21097 3007 21131
rect 3007 21097 3016 21131
rect 2964 21088 3016 21097
rect 3240 21131 3292 21140
rect 3240 21097 3249 21131
rect 3249 21097 3283 21131
rect 3283 21097 3292 21131
rect 3240 21088 3292 21097
rect 3332 21088 3384 21140
rect 4436 21131 4488 21140
rect 4436 21097 4445 21131
rect 4445 21097 4479 21131
rect 4479 21097 4488 21131
rect 4436 21088 4488 21097
rect 2320 21020 2372 21072
rect 3976 21020 4028 21072
rect 4804 21088 4856 21140
rect 6920 21088 6972 21140
rect 8208 21088 8260 21140
rect 10048 21088 10100 21140
rect 6000 21020 6052 21072
rect 2136 20995 2188 21004
rect 2136 20961 2145 20995
rect 2145 20961 2179 20995
rect 2179 20961 2188 20995
rect 2136 20952 2188 20961
rect 5632 20952 5684 21004
rect 10968 20952 11020 21004
rect 4068 20884 4120 20936
rect 4528 20884 4580 20936
rect 9312 20884 9364 20936
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 4160 20816 4212 20868
rect 11152 20748 11204 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 2136 20587 2188 20596
rect 2136 20553 2145 20587
rect 2145 20553 2179 20587
rect 2179 20553 2188 20587
rect 2136 20544 2188 20553
rect 3976 20544 4028 20596
rect 4160 20544 4212 20596
rect 5632 20544 5684 20596
rect 4068 20476 4120 20528
rect 4252 20408 4304 20460
rect 11060 20544 11112 20596
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 9312 20451 9364 20460
rect 9312 20417 9321 20451
rect 9321 20417 9355 20451
rect 9355 20417 9364 20451
rect 9312 20408 9364 20417
rect 5264 20272 5316 20324
rect 5816 20272 5868 20324
rect 7104 20315 7156 20324
rect 7104 20281 7116 20315
rect 7116 20281 7156 20315
rect 7104 20272 7156 20281
rect 11152 20272 11204 20324
rect 4528 20204 4580 20256
rect 4988 20247 5040 20256
rect 4988 20213 4997 20247
rect 4997 20213 5031 20247
rect 5031 20213 5040 20247
rect 4988 20204 5040 20213
rect 6000 20204 6052 20256
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 10692 20247 10744 20256
rect 10692 20213 10701 20247
rect 10701 20213 10735 20247
rect 10735 20213 10744 20247
rect 10692 20204 10744 20213
rect 11520 20204 11572 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 4436 20000 4488 20052
rect 6736 20000 6788 20052
rect 6828 20000 6880 20052
rect 9312 20000 9364 20052
rect 10324 20043 10376 20052
rect 10324 20009 10333 20043
rect 10333 20009 10367 20043
rect 10367 20009 10376 20043
rect 10324 20000 10376 20009
rect 11060 20000 11112 20052
rect 6000 19932 6052 19984
rect 6276 19907 6328 19916
rect 6276 19873 6285 19907
rect 6285 19873 6319 19907
rect 6319 19873 6328 19907
rect 6276 19864 6328 19873
rect 6368 19907 6420 19916
rect 6368 19873 6377 19907
rect 6377 19873 6411 19907
rect 6411 19873 6420 19907
rect 6368 19864 6420 19873
rect 10968 19932 11020 19984
rect 10232 19864 10284 19916
rect 11520 19864 11572 19916
rect 8208 19796 8260 19848
rect 12440 19796 12492 19848
rect 2596 19703 2648 19712
rect 2596 19669 2605 19703
rect 2605 19669 2639 19703
rect 2639 19669 2648 19703
rect 2596 19660 2648 19669
rect 4436 19660 4488 19712
rect 8668 19703 8720 19712
rect 8668 19669 8677 19703
rect 8677 19669 8711 19703
rect 8711 19669 8720 19703
rect 8668 19660 8720 19669
rect 9680 19660 9732 19712
rect 9864 19703 9916 19712
rect 9864 19669 9873 19703
rect 9873 19669 9907 19703
rect 9907 19669 9916 19703
rect 9864 19660 9916 19669
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 13544 19660 13596 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 6000 19456 6052 19508
rect 9864 19388 9916 19440
rect 2596 19363 2648 19372
rect 2596 19329 2605 19363
rect 2605 19329 2639 19363
rect 2639 19329 2648 19363
rect 2596 19320 2648 19329
rect 3516 19184 3568 19236
rect 6368 19252 6420 19304
rect 9496 19252 9548 19304
rect 10692 19320 10744 19372
rect 11152 19320 11204 19372
rect 12532 19320 12584 19372
rect 9864 19252 9916 19304
rect 11060 19252 11112 19304
rect 12624 19252 12676 19304
rect 6276 19184 6328 19236
rect 7840 19184 7892 19236
rect 3976 19159 4028 19168
rect 3976 19125 3985 19159
rect 3985 19125 4019 19159
rect 4019 19125 4028 19159
rect 3976 19116 4028 19125
rect 6000 19159 6052 19168
rect 6000 19125 6009 19159
rect 6009 19125 6043 19159
rect 6043 19125 6052 19159
rect 6000 19116 6052 19125
rect 12072 19184 12124 19236
rect 6828 19116 6880 19168
rect 8392 19116 8444 19168
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 9404 19159 9456 19168
rect 9404 19125 9413 19159
rect 9413 19125 9447 19159
rect 9447 19125 9456 19159
rect 9404 19116 9456 19125
rect 9680 19116 9732 19168
rect 10048 19116 10100 19168
rect 10324 19116 10376 19168
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 11060 19116 11112 19168
rect 12348 19116 12400 19168
rect 12716 19116 12768 19168
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 2596 18955 2648 18964
rect 2596 18921 2605 18955
rect 2605 18921 2639 18955
rect 2639 18921 2648 18955
rect 2596 18912 2648 18921
rect 6184 18912 6236 18964
rect 7104 18955 7156 18964
rect 7104 18921 7113 18955
rect 7113 18921 7147 18955
rect 7147 18921 7156 18955
rect 7104 18912 7156 18921
rect 7656 18912 7708 18964
rect 11152 18955 11204 18964
rect 11152 18921 11161 18955
rect 11161 18921 11195 18955
rect 11195 18921 11204 18955
rect 11152 18912 11204 18921
rect 12072 18912 12124 18964
rect 12716 18912 12768 18964
rect 13452 18912 13504 18964
rect 1676 18887 1728 18896
rect 1676 18853 1685 18887
rect 1685 18853 1719 18887
rect 1719 18853 1728 18887
rect 1676 18844 1728 18853
rect 6000 18844 6052 18896
rect 6552 18844 6604 18896
rect 9496 18887 9548 18896
rect 9496 18853 9505 18887
rect 9505 18853 9539 18887
rect 9539 18853 9548 18887
rect 9496 18844 9548 18853
rect 10140 18844 10192 18896
rect 11336 18844 11388 18896
rect 6736 18776 6788 18828
rect 8024 18776 8076 18828
rect 8484 18776 8536 18828
rect 1676 18708 1728 18760
rect 6000 18708 6052 18760
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 9864 18776 9916 18828
rect 11060 18776 11112 18828
rect 8576 18708 8628 18717
rect 8668 18640 8720 18692
rect 5540 18572 5592 18624
rect 5816 18615 5868 18624
rect 5816 18581 5825 18615
rect 5825 18581 5859 18615
rect 5859 18581 5868 18615
rect 5816 18572 5868 18581
rect 7564 18615 7616 18624
rect 7564 18581 7573 18615
rect 7573 18581 7607 18615
rect 7607 18581 7616 18615
rect 7564 18572 7616 18581
rect 9496 18572 9548 18624
rect 10232 18708 10284 18760
rect 11152 18708 11204 18760
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 10324 18572 10376 18624
rect 10692 18615 10744 18624
rect 10692 18581 10701 18615
rect 10701 18581 10735 18615
rect 10735 18581 10744 18615
rect 10692 18572 10744 18581
rect 12624 18572 12676 18624
rect 12992 18572 13044 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 3516 18368 3568 18420
rect 4068 18368 4120 18420
rect 5356 18368 5408 18420
rect 6184 18411 6236 18420
rect 6184 18377 6193 18411
rect 6193 18377 6227 18411
rect 6227 18377 6236 18411
rect 6184 18368 6236 18377
rect 8576 18411 8628 18420
rect 8576 18377 8585 18411
rect 8585 18377 8619 18411
rect 8619 18377 8628 18411
rect 8576 18368 8628 18377
rect 10324 18368 10376 18420
rect 10968 18368 11020 18420
rect 11520 18368 11572 18420
rect 1676 18343 1728 18352
rect 1676 18309 1685 18343
rect 1685 18309 1719 18343
rect 1719 18309 1728 18343
rect 1676 18300 1728 18309
rect 7104 18343 7156 18352
rect 7104 18309 7113 18343
rect 7113 18309 7147 18343
rect 7147 18309 7156 18343
rect 7104 18300 7156 18309
rect 12072 18300 12124 18352
rect 12900 18300 12952 18352
rect 6000 18232 6052 18284
rect 7564 18275 7616 18284
rect 7564 18241 7573 18275
rect 7573 18241 7607 18275
rect 7607 18241 7616 18275
rect 7564 18232 7616 18241
rect 7656 18275 7708 18284
rect 7656 18241 7665 18275
rect 7665 18241 7699 18275
rect 7699 18241 7708 18275
rect 7656 18232 7708 18241
rect 8760 18232 8812 18284
rect 10876 18275 10928 18284
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 12440 18232 12492 18284
rect 13084 18275 13136 18284
rect 2596 18164 2648 18216
rect 5356 18164 5408 18216
rect 8668 18164 8720 18216
rect 9404 18164 9456 18216
rect 9496 18164 9548 18216
rect 10600 18164 10652 18216
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 4344 18096 4396 18148
rect 5540 18139 5592 18148
rect 5540 18105 5549 18139
rect 5549 18105 5583 18139
rect 5583 18105 5592 18139
rect 5540 18096 5592 18105
rect 11152 18096 11204 18148
rect 5448 18028 5500 18080
rect 6736 18028 6788 18080
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 8484 18028 8536 18080
rect 8668 18028 8720 18080
rect 10140 18071 10192 18080
rect 10140 18037 10149 18071
rect 10149 18037 10183 18071
rect 10183 18037 10192 18071
rect 10140 18028 10192 18037
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 11060 18028 11112 18080
rect 12348 18028 12400 18080
rect 12900 18071 12952 18080
rect 12900 18037 12909 18071
rect 12909 18037 12943 18071
rect 12943 18037 12952 18071
rect 12900 18028 12952 18037
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 3424 17824 3476 17876
rect 5172 17824 5224 17876
rect 7656 17824 7708 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 9864 17824 9916 17876
rect 10876 17824 10928 17876
rect 12348 17824 12400 17876
rect 3976 17756 4028 17808
rect 9496 17799 9548 17808
rect 9496 17765 9505 17799
rect 9505 17765 9539 17799
rect 9539 17765 9548 17799
rect 9496 17756 9548 17765
rect 10232 17756 10284 17808
rect 12072 17799 12124 17808
rect 12072 17765 12081 17799
rect 12081 17765 12115 17799
rect 12115 17765 12124 17799
rect 12072 17756 12124 17765
rect 12256 17756 12308 17808
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 3332 17620 3384 17672
rect 7380 17688 7432 17740
rect 9312 17688 9364 17740
rect 9772 17688 9824 17740
rect 6828 17663 6880 17672
rect 2596 17552 2648 17604
rect 3424 17552 3476 17604
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 12992 17620 13044 17672
rect 11152 17552 11204 17604
rect 13084 17552 13136 17604
rect 1860 17484 1912 17536
rect 3516 17527 3568 17536
rect 3516 17493 3525 17527
rect 3525 17493 3559 17527
rect 3559 17493 3568 17527
rect 3516 17484 3568 17493
rect 6000 17484 6052 17536
rect 7472 17484 7524 17536
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 8760 17484 8812 17493
rect 11060 17527 11112 17536
rect 11060 17493 11069 17527
rect 11069 17493 11103 17527
rect 11103 17493 11112 17527
rect 12716 17527 12768 17536
rect 11060 17484 11112 17493
rect 12716 17493 12725 17527
rect 12725 17493 12759 17527
rect 12759 17493 12768 17527
rect 12716 17484 12768 17493
rect 12808 17484 12860 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 2780 17280 2832 17332
rect 4896 17323 4948 17332
rect 4896 17289 4905 17323
rect 4905 17289 4939 17323
rect 4939 17289 4948 17323
rect 4896 17280 4948 17289
rect 7472 17280 7524 17332
rect 9496 17280 9548 17332
rect 9864 17280 9916 17332
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 11152 17280 11204 17332
rect 12256 17323 12308 17332
rect 12256 17289 12265 17323
rect 12265 17289 12299 17323
rect 12299 17289 12308 17323
rect 12256 17280 12308 17289
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 3332 17255 3384 17264
rect 3332 17221 3341 17255
rect 3341 17221 3375 17255
rect 3375 17221 3384 17255
rect 3332 17212 3384 17221
rect 1584 17187 1636 17196
rect 1584 17153 1593 17187
rect 1593 17153 1627 17187
rect 1627 17153 1636 17187
rect 1584 17144 1636 17153
rect 3516 17144 3568 17196
rect 6092 17212 6144 17264
rect 6736 17212 6788 17264
rect 12808 17212 12860 17264
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 4344 17144 4396 17196
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 10968 17144 11020 17196
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 4896 17076 4948 17128
rect 10416 17076 10468 17128
rect 10784 17076 10836 17128
rect 11060 17076 11112 17128
rect 12808 17119 12860 17128
rect 12808 17085 12817 17119
rect 12817 17085 12851 17119
rect 12851 17085 12860 17119
rect 12808 17076 12860 17085
rect 4160 17008 4212 17060
rect 4528 17008 4580 17060
rect 9496 17008 9548 17060
rect 9772 17008 9824 17060
rect 4252 16940 4304 16992
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 6092 16940 6144 16992
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 8852 16940 8904 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 1400 16736 1452 16788
rect 2872 16736 2924 16788
rect 3424 16736 3476 16788
rect 4160 16779 4212 16788
rect 4160 16745 4169 16779
rect 4169 16745 4203 16779
rect 4203 16745 4212 16779
rect 4160 16736 4212 16745
rect 4528 16779 4580 16788
rect 4528 16745 4537 16779
rect 4537 16745 4571 16779
rect 4571 16745 4580 16779
rect 4528 16736 4580 16745
rect 4804 16736 4856 16788
rect 5540 16779 5592 16788
rect 5540 16745 5549 16779
rect 5549 16745 5583 16779
rect 5583 16745 5592 16779
rect 5540 16736 5592 16745
rect 3240 16600 3292 16652
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 2964 16532 3016 16584
rect 4068 16668 4120 16720
rect 6092 16736 6144 16788
rect 6828 16736 6880 16788
rect 8024 16736 8076 16788
rect 8484 16736 8536 16788
rect 9404 16736 9456 16788
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 12072 16736 12124 16788
rect 12716 16736 12768 16788
rect 6000 16711 6052 16720
rect 6000 16677 6034 16711
rect 6034 16677 6052 16711
rect 6000 16668 6052 16677
rect 6184 16668 6236 16720
rect 8852 16600 8904 16652
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 4344 16532 4396 16584
rect 4988 16532 5040 16584
rect 10048 16532 10100 16584
rect 11060 16600 11112 16652
rect 12072 16600 12124 16652
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 11888 16532 11940 16584
rect 6000 16396 6052 16448
rect 11152 16396 11204 16448
rect 12900 16396 12952 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 4528 16235 4580 16244
rect 4528 16201 4537 16235
rect 4537 16201 4571 16235
rect 4571 16201 4580 16235
rect 4528 16192 4580 16201
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 6552 16192 6604 16244
rect 6828 16192 6880 16244
rect 6920 16192 6972 16244
rect 8760 16192 8812 16244
rect 11060 16192 11112 16244
rect 12072 16235 12124 16244
rect 12072 16201 12081 16235
rect 12081 16201 12115 16235
rect 12115 16201 12124 16235
rect 12072 16192 12124 16201
rect 4804 16124 4856 16176
rect 10968 16124 11020 16176
rect 2964 16056 3016 16108
rect 5540 16056 5592 16108
rect 6000 16056 6052 16108
rect 7748 16031 7800 16040
rect 7748 15997 7757 16031
rect 7757 15997 7791 16031
rect 7791 15997 7800 16031
rect 7748 15988 7800 15997
rect 12072 16056 12124 16108
rect 8576 15988 8628 16040
rect 9680 15988 9732 16040
rect 11336 15988 11388 16040
rect 11888 15988 11940 16040
rect 5816 15920 5868 15972
rect 10600 15963 10652 15972
rect 10600 15929 10609 15963
rect 10609 15929 10643 15963
rect 10643 15929 10652 15963
rect 10600 15920 10652 15929
rect 2596 15852 2648 15904
rect 2872 15852 2924 15904
rect 3240 15895 3292 15904
rect 3240 15861 3249 15895
rect 3249 15861 3283 15895
rect 3283 15861 3292 15895
rect 3240 15852 3292 15861
rect 4068 15852 4120 15904
rect 5448 15852 5500 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 11336 15852 11388 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 6000 15648 6052 15700
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 8024 15691 8076 15700
rect 8024 15657 8033 15691
rect 8033 15657 8067 15691
rect 8067 15657 8076 15691
rect 8024 15648 8076 15657
rect 8576 15648 8628 15700
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 10692 15648 10744 15700
rect 12072 15648 12124 15700
rect 5908 15512 5960 15564
rect 7288 15512 7340 15564
rect 8392 15555 8444 15564
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 8484 15555 8536 15564
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 10416 15555 10468 15564
rect 8484 15512 8536 15521
rect 10416 15521 10425 15555
rect 10425 15521 10459 15555
rect 10459 15521 10468 15555
rect 10416 15512 10468 15521
rect 5172 15444 5224 15496
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6184 15444 6236 15496
rect 6368 15444 6420 15496
rect 8208 15444 8260 15496
rect 11152 15512 11204 15564
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 8484 15376 8536 15428
rect 9588 15376 9640 15428
rect 11060 15444 11112 15496
rect 11336 15444 11388 15496
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 5908 15104 5960 15156
rect 6368 15147 6420 15156
rect 6368 15113 6377 15147
rect 6377 15113 6411 15147
rect 6411 15113 6420 15147
rect 6368 15104 6420 15113
rect 8208 15104 8260 15156
rect 8300 15104 8352 15156
rect 8852 15147 8904 15156
rect 8852 15113 8861 15147
rect 8861 15113 8895 15147
rect 8895 15113 8904 15147
rect 8852 15104 8904 15113
rect 10324 15104 10376 15156
rect 9772 15036 9824 15088
rect 10692 15036 10744 15088
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 8300 14968 8352 15020
rect 8576 14968 8628 15020
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 1768 14900 1820 14952
rect 6092 14900 6144 14952
rect 8852 14900 8904 14952
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 9588 14832 9640 14884
rect 11336 14832 11388 14884
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 10048 14764 10100 14816
rect 10232 14807 10284 14816
rect 10232 14773 10241 14807
rect 10241 14773 10275 14807
rect 10275 14773 10284 14807
rect 10232 14764 10284 14773
rect 11152 14764 11204 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 2596 14560 2648 14612
rect 3424 14603 3476 14612
rect 3424 14569 3433 14603
rect 3433 14569 3467 14603
rect 3467 14569 3476 14603
rect 3424 14560 3476 14569
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 4712 14560 4764 14612
rect 5632 14560 5684 14612
rect 8300 14603 8352 14612
rect 8300 14569 8309 14603
rect 8309 14569 8343 14603
rect 8343 14569 8352 14603
rect 8300 14560 8352 14569
rect 5540 14492 5592 14544
rect 5816 14492 5868 14544
rect 7656 14492 7708 14544
rect 9312 14560 9364 14612
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 11060 14560 11112 14612
rect 13544 14535 13596 14544
rect 13544 14501 13553 14535
rect 13553 14501 13587 14535
rect 13587 14501 13596 14535
rect 13544 14492 13596 14501
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 2504 14356 2556 14408
rect 3240 14424 3292 14476
rect 4344 14424 4396 14476
rect 1952 14288 2004 14340
rect 4068 14356 4120 14408
rect 7196 14424 7248 14476
rect 8024 14424 8076 14476
rect 13268 14467 13320 14476
rect 13268 14433 13277 14467
rect 13277 14433 13311 14467
rect 13311 14433 13320 14467
rect 13268 14424 13320 14433
rect 4988 14356 5040 14408
rect 6092 14356 6144 14408
rect 7472 14356 7524 14408
rect 7012 14331 7064 14340
rect 7012 14297 7021 14331
rect 7021 14297 7055 14331
rect 7055 14297 7064 14331
rect 8576 14356 8628 14408
rect 10416 14356 10468 14408
rect 7012 14288 7064 14297
rect 10232 14288 10284 14340
rect 1768 14220 1820 14272
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 5540 14220 5592 14272
rect 7288 14220 7340 14272
rect 7748 14220 7800 14272
rect 8116 14220 8168 14272
rect 10048 14220 10100 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 1952 14016 2004 14068
rect 2504 14016 2556 14068
rect 3240 14059 3292 14068
rect 3240 14025 3249 14059
rect 3249 14025 3283 14059
rect 3283 14025 3292 14059
rect 3240 14016 3292 14025
rect 4712 14016 4764 14068
rect 4988 14016 5040 14068
rect 5816 14016 5868 14068
rect 6092 14059 6144 14068
rect 6092 14025 6101 14059
rect 6101 14025 6135 14059
rect 6135 14025 6144 14059
rect 6092 14016 6144 14025
rect 8024 14016 8076 14068
rect 3424 13948 3476 14000
rect 2228 13880 2280 13932
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 2596 13812 2648 13821
rect 2412 13676 2464 13728
rect 2596 13676 2648 13728
rect 3424 13812 3476 13864
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 3516 13744 3568 13796
rect 6092 13744 6144 13796
rect 7012 13812 7064 13864
rect 8576 13812 8628 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 8300 13719 8352 13728
rect 8300 13685 8309 13719
rect 8309 13685 8343 13719
rect 8343 13685 8352 13719
rect 8300 13676 8352 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 2320 13472 2372 13524
rect 2780 13472 2832 13524
rect 4068 13515 4120 13524
rect 4068 13481 4077 13515
rect 4077 13481 4111 13515
rect 4111 13481 4120 13515
rect 4068 13472 4120 13481
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 6092 13472 6144 13524
rect 7840 13472 7892 13524
rect 8116 13472 8168 13524
rect 4528 13447 4580 13456
rect 4528 13413 4537 13447
rect 4537 13413 4571 13447
rect 4571 13413 4580 13447
rect 4528 13404 4580 13413
rect 6460 13404 6512 13456
rect 7472 13404 7524 13456
rect 2596 13336 2648 13388
rect 2872 13379 2924 13388
rect 2872 13345 2881 13379
rect 2881 13345 2915 13379
rect 2915 13345 2924 13379
rect 2872 13336 2924 13345
rect 4712 13336 4764 13388
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 12072 13404 12124 13456
rect 7840 13336 7892 13388
rect 10048 13336 10100 13388
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 8760 13268 8812 13320
rect 9956 13268 10008 13320
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 11336 13268 11388 13320
rect 3516 13132 3568 13184
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 5816 13200 5868 13252
rect 7840 13243 7892 13252
rect 7840 13209 7849 13243
rect 7849 13209 7883 13243
rect 7883 13209 7892 13243
rect 7840 13200 7892 13209
rect 9312 13132 9364 13184
rect 9772 13132 9824 13184
rect 10508 13132 10560 13184
rect 10968 13175 11020 13184
rect 10968 13141 10977 13175
rect 10977 13141 11011 13175
rect 11011 13141 11020 13175
rect 10968 13132 11020 13141
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 2872 12928 2924 12980
rect 4528 12928 4580 12980
rect 7288 12928 7340 12980
rect 9680 12928 9732 12980
rect 10600 12928 10652 12980
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 7472 12860 7524 12912
rect 11336 12860 11388 12912
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 5172 12792 5224 12844
rect 7840 12792 7892 12844
rect 10968 12835 11020 12844
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 8300 12767 8352 12776
rect 8300 12733 8334 12767
rect 8334 12733 8352 12767
rect 2504 12699 2556 12708
rect 2504 12665 2516 12699
rect 2516 12665 2556 12699
rect 2504 12656 2556 12665
rect 4528 12656 4580 12708
rect 5080 12656 5132 12708
rect 5540 12656 5592 12708
rect 6460 12656 6512 12708
rect 8300 12724 8352 12733
rect 8116 12656 8168 12708
rect 8392 12656 8444 12708
rect 2964 12588 3016 12640
rect 3516 12588 3568 12640
rect 4712 12588 4764 12640
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 5448 12588 5500 12640
rect 9496 12656 9548 12708
rect 8668 12588 8720 12640
rect 8760 12588 8812 12640
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 12072 12588 12124 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 5172 12384 5224 12436
rect 5632 12384 5684 12436
rect 7104 12427 7156 12436
rect 7104 12393 7113 12427
rect 7113 12393 7147 12427
rect 7147 12393 7156 12427
rect 7104 12384 7156 12393
rect 7196 12384 7248 12436
rect 8668 12384 8720 12436
rect 9956 12427 10008 12436
rect 9956 12393 9965 12427
rect 9965 12393 9999 12427
rect 9999 12393 10008 12427
rect 9956 12384 10008 12393
rect 10968 12384 11020 12436
rect 11980 12384 12032 12436
rect 13084 12384 13136 12436
rect 1676 12359 1728 12368
rect 1676 12325 1685 12359
rect 1685 12325 1719 12359
rect 1719 12325 1728 12359
rect 1676 12316 1728 12325
rect 3240 12316 3292 12368
rect 5724 12316 5776 12368
rect 6184 12316 6236 12368
rect 8116 12316 8168 12368
rect 11428 12316 11480 12368
rect 11520 12316 11572 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 10416 12291 10468 12300
rect 2964 12180 3016 12232
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 7748 12180 7800 12232
rect 8208 12180 8260 12232
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 10048 12180 10100 12232
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 11060 12180 11112 12232
rect 11336 12180 11388 12232
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 9956 12112 10008 12164
rect 11428 12112 11480 12164
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 4988 12044 5040 12096
rect 5172 12044 5224 12096
rect 5448 12044 5500 12096
rect 11152 12087 11204 12096
rect 11152 12053 11161 12087
rect 11161 12053 11195 12087
rect 11195 12053 11204 12087
rect 11152 12044 11204 12053
rect 11796 12044 11848 12096
rect 12992 12087 13044 12096
rect 12992 12053 13001 12087
rect 13001 12053 13035 12087
rect 13035 12053 13044 12087
rect 12992 12044 13044 12053
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 2320 11840 2372 11892
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 7288 11840 7340 11892
rect 10048 11883 10100 11892
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 10508 11840 10560 11892
rect 11152 11840 11204 11892
rect 12624 11840 12676 11892
rect 13360 11840 13412 11892
rect 10692 11815 10744 11824
rect 10692 11781 10701 11815
rect 10701 11781 10735 11815
rect 10735 11781 10744 11815
rect 10692 11772 10744 11781
rect 12072 11772 12124 11824
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 3240 11704 3292 11756
rect 4804 11704 4856 11756
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 7840 11704 7892 11756
rect 8024 11704 8076 11756
rect 8392 11704 8444 11756
rect 11520 11704 11572 11756
rect 12992 11704 13044 11756
rect 5356 11636 5408 11688
rect 7104 11636 7156 11688
rect 8760 11636 8812 11688
rect 11060 11636 11112 11688
rect 11796 11636 11848 11688
rect 5448 11568 5500 11620
rect 11612 11568 11664 11620
rect 12532 11568 12584 11620
rect 13360 11568 13412 11620
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 7104 11500 7156 11552
rect 8208 11500 8260 11552
rect 8668 11500 8720 11552
rect 9772 11500 9824 11552
rect 11244 11500 11296 11552
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 12992 11500 13044 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 1768 11296 1820 11348
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 3608 11296 3660 11348
rect 5080 11296 5132 11348
rect 5172 11296 5224 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 5908 11339 5960 11348
rect 5908 11305 5917 11339
rect 5917 11305 5951 11339
rect 5951 11305 5960 11339
rect 5908 11296 5960 11305
rect 7196 11296 7248 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 11520 11296 11572 11348
rect 12808 11296 12860 11348
rect 7656 11228 7708 11280
rect 7932 11228 7984 11280
rect 8392 11228 8444 11280
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 7840 11203 7892 11212
rect 7840 11169 7849 11203
rect 7849 11169 7883 11203
rect 7883 11169 7892 11203
rect 7840 11160 7892 11169
rect 10416 11228 10468 11280
rect 11244 11228 11296 11280
rect 12624 11271 12676 11280
rect 12624 11237 12633 11271
rect 12633 11237 12667 11271
rect 12667 11237 12676 11271
rect 12624 11228 12676 11237
rect 9772 11160 9824 11212
rect 9956 11203 10008 11212
rect 9956 11169 9990 11203
rect 9990 11169 10008 11203
rect 9956 11160 10008 11169
rect 12532 11203 12584 11212
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12532 11160 12584 11169
rect 4896 11092 4948 11144
rect 5632 11092 5684 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 11520 11092 11572 11144
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 12348 11024 12400 11076
rect 6184 10956 6236 11008
rect 6736 10956 6788 11008
rect 12992 11024 13044 11076
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 5632 10795 5684 10804
rect 5632 10761 5641 10795
rect 5641 10761 5675 10795
rect 5675 10761 5684 10795
rect 5632 10752 5684 10761
rect 5816 10752 5868 10804
rect 7932 10752 7984 10804
rect 9956 10752 10008 10804
rect 10416 10752 10468 10804
rect 11520 10752 11572 10804
rect 12072 10752 12124 10804
rect 12716 10752 12768 10804
rect 2596 10684 2648 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 4068 10616 4120 10668
rect 1768 10548 1820 10600
rect 4804 10548 4856 10600
rect 3332 10523 3384 10532
rect 3332 10489 3341 10523
rect 3341 10489 3375 10523
rect 3375 10489 3384 10523
rect 3332 10480 3384 10489
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 5724 10684 5776 10736
rect 6736 10684 6788 10736
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 12532 10616 12584 10668
rect 9404 10548 9456 10600
rect 6184 10480 6236 10532
rect 10508 10480 10560 10532
rect 4896 10455 4948 10464
rect 4896 10421 4905 10455
rect 4905 10421 4939 10455
rect 4939 10421 4948 10455
rect 4896 10412 4948 10421
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 8116 10412 8168 10464
rect 9404 10412 9456 10464
rect 9864 10412 9916 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 3332 10251 3384 10260
rect 3332 10217 3341 10251
rect 3341 10217 3375 10251
rect 3375 10217 3384 10251
rect 3332 10208 3384 10217
rect 3424 10208 3476 10260
rect 5172 10208 5224 10260
rect 5908 10208 5960 10260
rect 6828 10208 6880 10260
rect 7840 10208 7892 10260
rect 9772 10208 9824 10260
rect 12348 10208 12400 10260
rect 6184 10140 6236 10192
rect 13084 10140 13136 10192
rect 1676 10072 1728 10124
rect 8024 10072 8076 10124
rect 8392 10115 8444 10124
rect 8392 10081 8401 10115
rect 8401 10081 8435 10115
rect 8435 10081 8444 10115
rect 8392 10072 8444 10081
rect 11520 10072 11572 10124
rect 12348 10072 12400 10124
rect 12440 10072 12492 10124
rect 2044 10004 2096 10056
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 4160 10004 4212 10056
rect 6736 10047 6788 10056
rect 2412 9936 2464 9988
rect 4804 9936 4856 9988
rect 6736 10013 6745 10047
rect 6745 10013 6779 10047
rect 6779 10013 6788 10047
rect 6736 10004 6788 10013
rect 8484 10047 8536 10056
rect 8484 10013 8493 10047
rect 8493 10013 8527 10047
rect 8527 10013 8536 10047
rect 8484 10004 8536 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 5816 9936 5868 9988
rect 7840 9936 7892 9988
rect 1400 9868 1452 9920
rect 2136 9868 2188 9920
rect 2320 9911 2372 9920
rect 2320 9877 2329 9911
rect 2329 9877 2363 9911
rect 2363 9877 2372 9911
rect 2320 9868 2372 9877
rect 10508 9868 10560 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 1676 9707 1728 9716
rect 1676 9673 1685 9707
rect 1685 9673 1719 9707
rect 1719 9673 1728 9707
rect 1676 9664 1728 9673
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 6184 9707 6236 9716
rect 6184 9673 6193 9707
rect 6193 9673 6227 9707
rect 6227 9673 6236 9707
rect 6184 9664 6236 9673
rect 8392 9664 8444 9716
rect 4068 9596 4120 9648
rect 5080 9596 5132 9648
rect 6460 9639 6512 9648
rect 6460 9605 6469 9639
rect 6469 9605 6503 9639
rect 6503 9605 6512 9639
rect 6460 9596 6512 9605
rect 6920 9596 6972 9648
rect 2136 9528 2188 9580
rect 3424 9460 3476 9512
rect 5172 9460 5224 9512
rect 5264 9460 5316 9512
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 12072 9664 12124 9716
rect 12348 9596 12400 9648
rect 7380 9460 7432 9512
rect 8576 9460 8628 9512
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 7012 9392 7064 9444
rect 8484 9392 8536 9444
rect 9404 9392 9456 9444
rect 1768 9324 1820 9376
rect 2412 9324 2464 9376
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 4160 9324 4212 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 10968 9324 11020 9376
rect 11520 9324 11572 9376
rect 12072 9324 12124 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 2504 9120 2556 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 4896 9120 4948 9172
rect 5264 9163 5316 9172
rect 5264 9129 5273 9163
rect 5273 9129 5307 9163
rect 5307 9129 5316 9163
rect 5264 9120 5316 9129
rect 5540 9120 5592 9172
rect 6736 9163 6788 9172
rect 6736 9129 6745 9163
rect 6745 9129 6779 9163
rect 6779 9129 6788 9163
rect 6736 9120 6788 9129
rect 7104 9120 7156 9172
rect 2136 9052 2188 9104
rect 5724 9052 5776 9104
rect 7012 9052 7064 9104
rect 1768 9027 1820 9036
rect 1768 8993 1802 9027
rect 1802 8993 1820 9027
rect 1768 8984 1820 8993
rect 3424 8984 3476 9036
rect 5172 8984 5224 9036
rect 6184 8984 6236 9036
rect 8760 8984 8812 9036
rect 9312 8984 9364 9036
rect 2780 8916 2832 8968
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 7288 8916 7340 8968
rect 8576 8916 8628 8968
rect 10232 8780 10284 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 2044 8576 2096 8628
rect 4896 8576 4948 8628
rect 6184 8619 6236 8628
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 6736 8576 6788 8628
rect 8760 8619 8812 8628
rect 8760 8585 8769 8619
rect 8769 8585 8803 8619
rect 8803 8585 8812 8619
rect 8760 8576 8812 8585
rect 8852 8576 8904 8628
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 2780 8304 2832 8356
rect 3424 8440 3476 8492
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 8760 8372 8812 8424
rect 9496 8372 9548 8424
rect 10232 8440 10284 8492
rect 10140 8372 10192 8424
rect 4804 8304 4856 8356
rect 3700 8279 3752 8288
rect 3700 8245 3709 8279
rect 3709 8245 3743 8279
rect 3743 8245 3752 8279
rect 3700 8236 3752 8245
rect 7196 8236 7248 8288
rect 7840 8236 7892 8288
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 9496 8236 9548 8288
rect 10692 8236 10744 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 1676 8032 1728 8084
rect 3700 8032 3752 8084
rect 4528 8032 4580 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 6644 8032 6696 8084
rect 7288 8032 7340 8084
rect 8576 8032 8628 8084
rect 2596 7964 2648 8016
rect 2964 7964 3016 8016
rect 1768 7896 1820 7948
rect 3332 7896 3384 7948
rect 4344 7896 4396 7948
rect 8300 7964 8352 8016
rect 2780 7760 2832 7812
rect 4068 7828 4120 7880
rect 7196 7896 7248 7948
rect 9864 7896 9916 7948
rect 4804 7828 4856 7880
rect 6828 7828 6880 7880
rect 9772 7828 9824 7880
rect 10232 7828 10284 7880
rect 11980 7939 12032 7948
rect 11980 7905 12014 7939
rect 12014 7905 12032 7939
rect 11980 7896 12032 7905
rect 8300 7760 8352 7812
rect 9496 7760 9548 7812
rect 7840 7692 7892 7744
rect 9312 7692 9364 7744
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 11520 7735 11572 7744
rect 11520 7701 11529 7735
rect 11529 7701 11563 7735
rect 11563 7701 11572 7735
rect 11520 7692 11572 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 1400 7488 1452 7540
rect 4068 7531 4120 7540
rect 4068 7497 4077 7531
rect 4077 7497 4111 7531
rect 4111 7497 4120 7531
rect 4068 7488 4120 7497
rect 5080 7488 5132 7540
rect 6828 7488 6880 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 2504 7420 2556 7472
rect 4252 7420 4304 7472
rect 4620 7420 4672 7472
rect 9588 7488 9640 7540
rect 11980 7488 12032 7540
rect 9220 7420 9272 7472
rect 9864 7420 9916 7472
rect 13268 7488 13320 7540
rect 12900 7420 12952 7472
rect 12808 7352 12860 7404
rect 13268 7352 13320 7404
rect 2596 7284 2648 7336
rect 3332 7327 3384 7336
rect 3332 7293 3341 7327
rect 3341 7293 3375 7327
rect 3375 7293 3384 7327
rect 3332 7284 3384 7293
rect 4804 7284 4856 7336
rect 5080 7284 5132 7336
rect 7472 7284 7524 7336
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 9128 7284 9180 7336
rect 9680 7284 9732 7336
rect 10692 7284 10744 7336
rect 11520 7284 11572 7336
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 4344 7148 4396 7200
rect 4528 7148 4580 7200
rect 5172 7148 5224 7200
rect 6920 7148 6972 7200
rect 7840 7148 7892 7200
rect 10232 7216 10284 7268
rect 12900 7259 12952 7268
rect 12900 7225 12909 7259
rect 12909 7225 12943 7259
rect 12943 7225 12952 7259
rect 12900 7216 12952 7225
rect 8484 7148 8536 7200
rect 9220 7148 9272 7200
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 12624 7148 12676 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 2228 6944 2280 6996
rect 2780 6944 2832 6996
rect 7196 6987 7248 6996
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 8208 6944 8260 6996
rect 9128 6987 9180 6996
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 9220 6944 9272 6996
rect 10508 6944 10560 6996
rect 12808 6987 12860 6996
rect 12808 6953 12817 6987
rect 12817 6953 12851 6987
rect 12851 6953 12860 6987
rect 12808 6944 12860 6953
rect 2136 6808 2188 6860
rect 2504 6808 2556 6860
rect 4712 6808 4764 6860
rect 5172 6851 5224 6860
rect 5172 6817 5181 6851
rect 5181 6817 5215 6851
rect 5215 6817 5224 6851
rect 5172 6808 5224 6817
rect 6092 6808 6144 6860
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 9956 6808 10008 6860
rect 11704 6851 11756 6860
rect 11704 6817 11727 6851
rect 11727 6817 11756 6851
rect 11704 6808 11756 6817
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 8668 6783 8720 6792
rect 8668 6749 8677 6783
rect 8677 6749 8711 6783
rect 8711 6749 8720 6783
rect 8668 6740 8720 6749
rect 9496 6715 9548 6724
rect 9496 6681 9505 6715
rect 9505 6681 9539 6715
rect 9539 6681 9548 6715
rect 9496 6672 9548 6681
rect 10232 6672 10284 6724
rect 940 6604 992 6656
rect 5448 6604 5500 6656
rect 6184 6604 6236 6656
rect 8576 6604 8628 6656
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 11612 6604 11664 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 1400 6332 1452 6384
rect 3332 6400 3384 6452
rect 5172 6443 5224 6452
rect 5172 6409 5181 6443
rect 5181 6409 5215 6443
rect 5215 6409 5224 6443
rect 5172 6400 5224 6409
rect 6092 6400 6144 6452
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 8392 6400 8444 6452
rect 9680 6400 9732 6452
rect 9956 6400 10008 6452
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 11704 6400 11756 6452
rect 3608 6375 3660 6384
rect 3608 6341 3617 6375
rect 3617 6341 3651 6375
rect 3651 6341 3660 6375
rect 3608 6332 3660 6341
rect 4988 6332 5040 6384
rect 6000 6332 6052 6384
rect 4712 6196 4764 6248
rect 9404 6264 9456 6316
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 11060 6264 11112 6316
rect 7564 6196 7616 6248
rect 13176 6196 13228 6248
rect 11980 6128 12032 6180
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 5816 6060 5868 6112
rect 7196 6103 7248 6112
rect 7196 6069 7205 6103
rect 7205 6069 7239 6103
rect 7239 6069 7248 6103
rect 7196 6060 7248 6069
rect 8668 6060 8720 6112
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11244 6103 11296 6112
rect 11244 6069 11253 6103
rect 11253 6069 11287 6103
rect 11287 6069 11296 6103
rect 11244 6060 11296 6069
rect 11520 6060 11572 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 7840 5856 7892 5908
rect 8484 5856 8536 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 10692 5899 10744 5908
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 8852 5788 8904 5840
rect 9588 5788 9640 5840
rect 2780 5720 2832 5772
rect 4344 5720 4396 5772
rect 5908 5720 5960 5772
rect 8392 5763 8444 5772
rect 8392 5729 8401 5763
rect 8401 5729 8435 5763
rect 8435 5729 8444 5763
rect 8392 5720 8444 5729
rect 11980 5720 12032 5772
rect 4252 5627 4304 5636
rect 4252 5593 4261 5627
rect 4261 5593 4295 5627
rect 4295 5593 4304 5627
rect 4252 5584 4304 5593
rect 8300 5652 8352 5704
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 8944 5652 8996 5704
rect 9404 5652 9456 5704
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 13084 5652 13136 5704
rect 7012 5584 7064 5636
rect 2228 5516 2280 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 6828 5516 6880 5568
rect 8208 5516 8260 5568
rect 11060 5584 11112 5636
rect 11152 5584 11204 5636
rect 12348 5584 12400 5636
rect 13176 5584 13228 5636
rect 11520 5516 11572 5568
rect 12716 5516 12768 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 2780 5312 2832 5364
rect 4804 5355 4856 5364
rect 4804 5321 4813 5355
rect 4813 5321 4847 5355
rect 4847 5321 4856 5355
rect 4804 5312 4856 5321
rect 6092 5355 6144 5364
rect 6092 5321 6101 5355
rect 6101 5321 6135 5355
rect 6135 5321 6144 5355
rect 6092 5312 6144 5321
rect 10784 5312 10836 5364
rect 11980 5355 12032 5364
rect 11980 5321 11989 5355
rect 11989 5321 12023 5355
rect 12023 5321 12032 5355
rect 11980 5312 12032 5321
rect 12624 5312 12676 5364
rect 10692 5244 10744 5296
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 13176 5176 13228 5228
rect 13452 5176 13504 5228
rect 13728 5176 13780 5228
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 3516 5108 3568 5160
rect 4528 5108 4580 5160
rect 6000 5108 6052 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 10048 5108 10100 5160
rect 11612 5108 11664 5160
rect 3976 5040 4028 5092
rect 5724 5083 5776 5092
rect 5724 5049 5733 5083
rect 5733 5049 5767 5083
rect 5767 5049 5776 5083
rect 5724 5040 5776 5049
rect 8024 5040 8076 5092
rect 8668 5040 8720 5092
rect 9588 5083 9640 5092
rect 9588 5049 9622 5083
rect 9622 5049 9640 5083
rect 9588 5040 9640 5049
rect 12716 5040 12768 5092
rect 7380 4972 7432 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 2136 4768 2188 4820
rect 3240 4768 3292 4820
rect 3516 4811 3568 4820
rect 3516 4777 3525 4811
rect 3525 4777 3559 4811
rect 3559 4777 3568 4811
rect 3516 4768 3568 4777
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 4528 4768 4580 4820
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 8208 4768 8260 4820
rect 9680 4768 9732 4820
rect 10600 4768 10652 4820
rect 11244 4768 11296 4820
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 6000 4700 6052 4752
rect 2780 4632 2832 4641
rect 5080 4632 5132 4684
rect 5540 4632 5592 4684
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 3976 4564 4028 4616
rect 8668 4632 8720 4684
rect 9312 4632 9364 4684
rect 10324 4632 10376 4684
rect 10784 4632 10836 4684
rect 11060 4632 11112 4684
rect 6368 4539 6420 4548
rect 6368 4505 6377 4539
rect 6377 4505 6411 4539
rect 6411 4505 6420 4539
rect 6368 4496 6420 4505
rect 7472 4539 7524 4548
rect 7472 4505 7481 4539
rect 7481 4505 7515 4539
rect 7515 4505 7524 4539
rect 7472 4496 7524 4505
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 8484 4564 8536 4616
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 10968 4564 11020 4616
rect 12900 4632 12952 4684
rect 13452 4632 13504 4684
rect 12440 4607 12492 4616
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 8392 4496 8444 4548
rect 12900 4496 12952 4548
rect 7288 4428 7340 4437
rect 8300 4428 8352 4480
rect 10048 4428 10100 4480
rect 11980 4428 12032 4480
rect 13544 4471 13596 4480
rect 13544 4437 13553 4471
rect 13553 4437 13587 4471
rect 13587 4437 13596 4471
rect 13544 4428 13596 4437
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 3976 4224 4028 4276
rect 9772 4224 9824 4276
rect 10600 4224 10652 4276
rect 10784 4267 10836 4276
rect 10784 4233 10793 4267
rect 10793 4233 10827 4267
rect 10827 4233 10836 4267
rect 10784 4224 10836 4233
rect 11888 4224 11940 4276
rect 12348 4224 12400 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 8024 4156 8076 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 6000 4088 6052 4140
rect 10692 4156 10744 4208
rect 1676 4020 1728 4072
rect 3148 4020 3200 4072
rect 3332 4063 3384 4072
rect 3332 4029 3366 4063
rect 3366 4029 3384 4063
rect 3332 4020 3384 4029
rect 6276 4020 6328 4072
rect 5080 3995 5132 4004
rect 5080 3961 5089 3995
rect 5089 3961 5123 3995
rect 5123 3961 5132 3995
rect 5080 3952 5132 3961
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 6736 3952 6788 4004
rect 7380 4020 7432 4072
rect 8484 4020 8536 4072
rect 9496 4020 9548 4072
rect 9680 4063 9732 4072
rect 9680 4029 9689 4063
rect 9689 4029 9723 4063
rect 9723 4029 9732 4063
rect 9680 4020 9732 4029
rect 10784 4020 10836 4072
rect 12072 4088 12124 4140
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 11980 4020 12032 4072
rect 12440 4020 12492 4072
rect 13452 4088 13504 4140
rect 9128 3952 9180 4004
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9496 3884 9548 3936
rect 11060 3927 11112 3936
rect 11060 3893 11069 3927
rect 11069 3893 11103 3927
rect 11103 3893 11112 3927
rect 11060 3884 11112 3893
rect 11980 3884 12032 3936
rect 12348 3884 12400 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 2688 3680 2740 3732
rect 3240 3680 3292 3732
rect 6828 3680 6880 3732
rect 7196 3680 7248 3732
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 8576 3680 8628 3732
rect 9496 3680 9548 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 13176 3680 13228 3732
rect 5080 3612 5132 3664
rect 6000 3655 6052 3664
rect 3424 3544 3476 3596
rect 4712 3544 4764 3596
rect 6000 3621 6009 3655
rect 6009 3621 6043 3655
rect 6043 3621 6052 3655
rect 6000 3612 6052 3621
rect 6736 3612 6788 3664
rect 2688 3476 2740 3528
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3332 3476 3384 3528
rect 5448 3476 5500 3528
rect 7840 3612 7892 3664
rect 8852 3655 8904 3664
rect 8852 3621 8861 3655
rect 8861 3621 8895 3655
rect 8895 3621 8904 3655
rect 8852 3612 8904 3621
rect 11980 3612 12032 3664
rect 8392 3544 8444 3596
rect 8760 3544 8812 3596
rect 10416 3476 10468 3528
rect 10692 3519 10744 3528
rect 10692 3485 10701 3519
rect 10701 3485 10735 3519
rect 10735 3485 10744 3519
rect 10692 3476 10744 3485
rect 10876 3476 10928 3528
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 5356 3408 5408 3460
rect 7012 3408 7064 3460
rect 7564 3408 7616 3460
rect 10968 3408 11020 3460
rect 4160 3340 4212 3392
rect 5080 3340 5132 3392
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 2872 3136 2924 3188
rect 6828 3136 6880 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 8208 3136 8260 3188
rect 8392 3136 8444 3188
rect 8760 3136 8812 3188
rect 9680 3136 9732 3188
rect 10416 3136 10468 3188
rect 11336 3136 11388 3188
rect 4712 3068 4764 3120
rect 10232 3068 10284 3120
rect 10968 3068 11020 3120
rect 11060 3068 11112 3120
rect 12716 3136 12768 3188
rect 4896 3000 4948 3052
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6828 3000 6880 3052
rect 13452 3000 13504 3052
rect 1676 2932 1728 2984
rect 3240 2932 3292 2984
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5264 2932 5316 2941
rect 7932 2932 7984 2984
rect 8208 2932 8260 2984
rect 1952 2907 2004 2916
rect 1952 2873 1961 2907
rect 1961 2873 1995 2907
rect 1995 2873 2004 2907
rect 1952 2864 2004 2873
rect 4436 2864 4488 2916
rect 6092 2864 6144 2916
rect 7840 2864 7892 2916
rect 8852 2932 8904 2984
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 13820 2975 13872 2984
rect 13820 2941 13829 2975
rect 13829 2941 13863 2975
rect 13863 2941 13872 2975
rect 13820 2932 13872 2941
rect 9588 2864 9640 2916
rect 13728 2864 13780 2916
rect 3516 2839 3568 2848
rect 3516 2805 3525 2839
rect 3525 2805 3559 2839
rect 3559 2805 3568 2839
rect 3516 2796 3568 2805
rect 13452 2839 13504 2848
rect 13452 2805 13461 2839
rect 13461 2805 13495 2839
rect 13495 2805 13504 2839
rect 13452 2796 13504 2805
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 2412 2635 2464 2644
rect 2412 2601 2421 2635
rect 2421 2601 2455 2635
rect 2455 2601 2464 2635
rect 2412 2592 2464 2601
rect 3332 2592 3384 2644
rect 3424 2592 3476 2644
rect 5172 2592 5224 2644
rect 6828 2592 6880 2644
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 4344 2567 4396 2576
rect 4344 2533 4353 2567
rect 4353 2533 4387 2567
rect 4387 2533 4396 2567
rect 4344 2524 4396 2533
rect 6092 2524 6144 2576
rect 10784 2592 10836 2644
rect 11980 2592 12032 2644
rect 12808 2592 12860 2644
rect 9128 2524 9180 2576
rect 10692 2524 10744 2576
rect 13084 2592 13136 2644
rect 13820 2592 13872 2644
rect 7932 2456 7984 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 9680 2456 9732 2508
rect 13636 2524 13688 2576
rect 4620 2388 4672 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 13452 2388 13504 2440
rect 2964 2320 3016 2372
rect 3332 2252 3384 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 5816 552 5868 604
rect 6920 552 6972 604
rect 7380 552 7432 604
rect 8024 552 8076 604
rect 10324 552 10376 604
rect 10600 552 10652 604
rect 12164 552 12216 604
rect 12348 552 12400 604
rect 12992 552 13044 604
rect 13268 552 13320 604
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39520 10194 40000
rect 10598 39520 10654 40000
rect 10966 39522 11022 40000
rect 11334 39522 11390 40000
rect 10704 39520 11022 39522
rect 11256 39520 11390 39522
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39520 13782 40000
rect 14186 39520 14242 40000
rect 14554 39520 14610 40000
rect 14922 39520 14978 40000
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 35834 244 39520
rect 204 35828 256 35834
rect 204 35770 256 35776
rect 584 34746 612 39520
rect 572 34740 624 34746
rect 572 34682 624 34688
rect 952 33658 980 39520
rect 1308 35828 1360 35834
rect 1308 35770 1360 35776
rect 1320 34218 1348 35770
rect 1412 34678 1440 39520
rect 1780 35290 1808 39520
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 2042 35184 2098 35193
rect 2042 35119 2098 35128
rect 1490 34912 1546 34921
rect 1490 34847 1546 34856
rect 1400 34672 1452 34678
rect 1400 34614 1452 34620
rect 1320 34202 1440 34218
rect 1320 34196 1452 34202
rect 1320 34190 1400 34196
rect 1400 34138 1452 34144
rect 940 33652 992 33658
rect 940 33594 992 33600
rect 1504 33046 1532 34847
rect 2056 34746 2084 35119
rect 2044 34740 2096 34746
rect 2044 34682 2096 34688
rect 2056 34542 2084 34682
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 2148 34202 2176 39520
rect 2412 35148 2464 35154
rect 2412 35090 2464 35096
rect 2424 34610 2452 35090
rect 2608 34746 2636 39520
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 2412 34604 2464 34610
rect 2412 34546 2464 34552
rect 2596 34604 2648 34610
rect 2596 34546 2648 34552
rect 2136 34196 2188 34202
rect 2136 34138 2188 34144
rect 1952 34060 2004 34066
rect 1952 34002 2004 34008
rect 1964 33658 1992 34002
rect 1952 33652 2004 33658
rect 1952 33594 2004 33600
rect 1964 33153 1992 33594
rect 2412 33312 2464 33318
rect 2412 33254 2464 33260
rect 1950 33144 2006 33153
rect 1950 33079 2006 33088
rect 1492 33040 1544 33046
rect 2424 33017 2452 33254
rect 1492 32982 1544 32988
rect 1674 33008 1730 33017
rect 2410 33008 2466 33017
rect 1674 32943 1730 32952
rect 1768 32972 1820 32978
rect 1688 31958 1716 32943
rect 2410 32943 2466 32952
rect 1768 32914 1820 32920
rect 1780 32230 1808 32914
rect 2608 32337 2636 34546
rect 2976 33658 3004 39520
rect 3146 38992 3202 39001
rect 3146 38927 3202 38936
rect 2964 33652 3016 33658
rect 2964 33594 3016 33600
rect 2780 33448 2832 33454
rect 2780 33390 2832 33396
rect 2792 33114 2820 33390
rect 2780 33108 2832 33114
rect 2832 33068 3004 33096
rect 2780 33050 2832 33056
rect 2594 32328 2650 32337
rect 2594 32263 2650 32272
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1676 31952 1728 31958
rect 1676 31894 1728 31900
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31414 1716 31758
rect 1676 31408 1728 31414
rect 1676 31350 1728 31356
rect 1688 31249 1716 31350
rect 1674 31240 1730 31249
rect 1674 31175 1730 31184
rect 1582 30968 1638 30977
rect 1582 30903 1638 30912
rect 1596 30258 1624 30903
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1400 29504 1452 29510
rect 1400 29446 1452 29452
rect 1412 29102 1440 29446
rect 1400 29096 1452 29102
rect 1400 29038 1452 29044
rect 1492 29028 1544 29034
rect 1492 28970 1544 28976
rect 1398 27976 1454 27985
rect 1398 27911 1454 27920
rect 1412 27538 1440 27911
rect 1400 27532 1452 27538
rect 1400 27474 1452 27480
rect 1412 27130 1440 27474
rect 1400 27124 1452 27130
rect 1400 27066 1452 27072
rect 1504 24993 1532 28970
rect 1674 28928 1730 28937
rect 1674 28863 1730 28872
rect 1584 28620 1636 28626
rect 1584 28562 1636 28568
rect 1596 28014 1624 28562
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1688 27606 1716 28863
rect 1676 27600 1728 27606
rect 1676 27542 1728 27548
rect 1582 27024 1638 27033
rect 1582 26959 1638 26968
rect 1596 25906 1624 26959
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1490 24984 1546 24993
rect 1490 24919 1546 24928
rect 1780 23089 1808 32166
rect 2226 30832 2282 30841
rect 2226 30767 2282 30776
rect 2240 30326 2268 30767
rect 2228 30320 2280 30326
rect 2228 30262 2280 30268
rect 2780 29776 2832 29782
rect 2780 29718 2832 29724
rect 2792 28762 2820 29718
rect 2976 29714 3004 33068
rect 2964 29708 3016 29714
rect 2964 29650 3016 29656
rect 2872 29640 2924 29646
rect 2872 29582 2924 29588
rect 3056 29640 3108 29646
rect 3056 29582 3108 29588
rect 2884 29306 2912 29582
rect 2872 29300 2924 29306
rect 2872 29242 2924 29248
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2884 28694 2912 29242
rect 3068 29238 3096 29582
rect 3056 29232 3108 29238
rect 3056 29174 3108 29180
rect 2872 28688 2924 28694
rect 2872 28630 2924 28636
rect 3160 28490 3188 38927
rect 3344 34610 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4016 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3422 36952 3478 36961
rect 3622 36944 3918 36964
rect 3422 36887 3478 36896
rect 3436 35057 3464 36887
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3988 35290 4016 37182
rect 3976 35284 4028 35290
rect 3976 35226 4028 35232
rect 4068 35148 4120 35154
rect 4068 35090 4120 35096
rect 3422 35048 3478 35057
rect 3422 34983 3478 34992
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3332 34604 3384 34610
rect 3332 34546 3384 34552
rect 3240 34536 3292 34542
rect 3240 34478 3292 34484
rect 3252 33561 3280 34478
rect 4080 34406 4108 35090
rect 4172 35018 4200 39520
rect 4540 35873 4568 39520
rect 4526 35864 4582 35873
rect 4526 35799 4582 35808
rect 4434 35184 4490 35193
rect 4434 35119 4490 35128
rect 4160 35012 4212 35018
rect 4160 34954 4212 34960
rect 4160 34604 4212 34610
rect 4160 34546 4212 34552
rect 4068 34400 4120 34406
rect 4068 34342 4120 34348
rect 4172 34202 4200 34546
rect 4344 34468 4396 34474
rect 4344 34410 4396 34416
rect 4160 34196 4212 34202
rect 4160 34138 4212 34144
rect 3332 34060 3384 34066
rect 3332 34002 3384 34008
rect 4068 34060 4120 34066
rect 4068 34002 4120 34008
rect 3238 33552 3294 33561
rect 3238 33487 3294 33496
rect 3344 33318 3372 34002
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3422 33552 3478 33561
rect 3422 33487 3478 33496
rect 3332 33312 3384 33318
rect 3332 33254 3384 33260
rect 3148 28484 3200 28490
rect 3148 28426 3200 28432
rect 2410 28112 2466 28121
rect 2410 28047 2412 28056
rect 2464 28047 2466 28056
rect 2412 28018 2464 28024
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2228 25696 2280 25702
rect 2226 25664 2228 25673
rect 2280 25664 2282 25673
rect 2226 25599 2282 25608
rect 1766 23080 1822 23089
rect 1766 23015 1822 23024
rect 2504 22976 2556 22982
rect 2318 22944 2374 22953
rect 2504 22918 2556 22924
rect 2318 22879 2374 22888
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 1674 21040 1730 21049
rect 2148 21010 2176 21830
rect 2332 21078 2360 22879
rect 2516 22642 2544 22918
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2412 21344 2464 21350
rect 2412 21286 2464 21292
rect 2424 21185 2452 21286
rect 2410 21176 2466 21185
rect 2410 21111 2466 21120
rect 2320 21072 2372 21078
rect 2320 21014 2372 21020
rect 1674 20975 1730 20984
rect 2136 21004 2188 21010
rect 1582 19000 1638 19009
rect 1582 18935 1638 18944
rect 1398 17232 1454 17241
rect 1596 17202 1624 18935
rect 1688 18902 1716 20975
rect 2136 20946 2188 20952
rect 2148 20602 2176 20946
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2608 19378 2636 19654
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2608 18970 2636 19314
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 1676 18896 1728 18902
rect 1676 18838 1728 18844
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1688 18358 1716 18702
rect 1676 18352 1728 18358
rect 1674 18320 1676 18329
rect 1728 18320 1730 18329
rect 1674 18255 1730 18264
rect 2608 18222 2636 18906
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2608 17610 2636 18158
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1398 17167 1454 17176
rect 1584 17196 1636 17202
rect 1412 17134 1440 17167
rect 1584 17138 1636 17144
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1412 16794 1440 17070
rect 1582 16960 1638 16969
rect 1582 16895 1638 16904
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1596 15026 1624 16895
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1768 14952 1820 14958
rect 1674 14920 1730 14929
rect 1768 14894 1820 14900
rect 1674 14855 1730 14864
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1398 12336 1454 12345
rect 1398 12271 1400 12280
rect 1452 12271 1454 12280
rect 1400 12242 1452 12248
rect 1596 11762 1624 12951
rect 1688 12374 1716 14855
rect 1780 14278 1808 14894
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1780 13977 1808 14214
rect 1766 13968 1822 13977
rect 1766 13903 1822 13912
rect 1872 13818 1900 17478
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2410 14920 2466 14929
rect 2410 14855 2466 14864
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1964 14074 1992 14282
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2240 13938 2268 14214
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 1780 13790 1900 13818
rect 1676 12368 1728 12374
rect 1676 12310 1728 12316
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1780 11354 1808 13790
rect 2424 13734 2452 14855
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 14414 2544 14758
rect 2608 14618 2636 15846
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2594 14376 2650 14385
rect 2516 14074 2544 14350
rect 2594 14311 2650 14320
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2608 13870 2636 14311
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2320 13524 2372 13530
rect 2424 13512 2452 13670
rect 2608 13512 2636 13670
rect 2372 13484 2452 13512
rect 2516 13484 2636 13512
rect 2320 13466 2372 13472
rect 2516 13410 2544 13484
rect 2240 13382 2544 13410
rect 2596 13388 2648 13394
rect 2240 12850 2268 13382
rect 2596 13330 2648 13336
rect 2608 13297 2636 13330
rect 2594 13288 2650 13297
rect 2424 13246 2594 13274
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2042 12336 2098 12345
rect 2042 12271 2098 12280
rect 2056 11354 2084 12271
rect 2240 11914 2268 12786
rect 2424 12102 2452 13246
rect 2594 13223 2650 13232
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2240 11898 2360 11914
rect 2240 11892 2372 11898
rect 2240 11886 2320 11892
rect 2320 11834 2372 11840
rect 2424 11370 2452 12038
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2240 11342 2452 11370
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1596 10674 1624 10911
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1780 10606 1808 11290
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 8430 1440 9862
rect 1688 9722 1716 10066
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2056 9722 2084 9998
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8498 1624 8871
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 7546 1440 8366
rect 1688 8090 1716 9658
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 9042 1808 9318
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1780 7954 1808 8978
rect 2056 8634 2084 9658
rect 2148 9586 2176 9862
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 9110 2176 9522
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2240 8922 2268 11342
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2148 8894 2268 8922
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 2148 6866 2176 8894
rect 2332 7410 2360 9862
rect 2424 9382 2452 9930
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2516 9178 2544 12650
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2516 7478 2544 9114
rect 2608 8022 2636 10678
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2320 7404 2372 7410
rect 2240 7364 2320 7392
rect 2240 7002 2268 7364
rect 2320 7346 2372 7352
rect 2608 7342 2636 7958
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2318 7032 2374 7041
rect 2228 6996 2280 7002
rect 2318 6967 2374 6976
rect 2228 6938 2280 6944
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 940 6656 992 6662
rect 940 6598 992 6604
rect 570 5672 626 5681
rect 570 5607 626 5616
rect 202 4176 258 4185
rect 202 4111 258 4120
rect 216 480 244 4111
rect 584 480 612 5607
rect 952 480 980 6598
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1412 480 1440 6326
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1582 4992 1638 5001
rect 1582 4927 1638 4936
rect 1596 4146 1624 4927
rect 2148 4826 2176 5102
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1688 4078 1716 4422
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1688 3641 1716 4014
rect 1766 3768 1822 3777
rect 1766 3703 1822 3712
rect 1674 3632 1730 3641
rect 1674 3567 1730 3576
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 2650 1716 2926
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1780 480 1808 3703
rect 1950 2952 2006 2961
rect 1950 2887 1952 2896
rect 2004 2887 2006 2896
rect 1952 2858 2004 2864
rect 2240 2802 2268 5510
rect 2332 5234 2360 6967
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 6118 2544 6802
rect 2504 6112 2556 6118
rect 2502 6080 2504 6089
rect 2556 6080 2558 6089
rect 2502 6015 2558 6024
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2700 3890 2728 27814
rect 3344 24154 3372 33254
rect 3436 29050 3464 33487
rect 4080 33318 4108 34002
rect 4068 33312 4120 33318
rect 4068 33254 4120 33260
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3976 32360 4028 32366
rect 3976 32302 4028 32308
rect 3988 31890 4016 32302
rect 3976 31884 4028 31890
rect 3976 31826 4028 31832
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 4252 31476 4304 31482
rect 4252 31418 4304 31424
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 4172 29866 4200 30534
rect 4080 29838 4200 29866
rect 4080 29782 4108 29838
rect 4068 29776 4120 29782
rect 4068 29718 4120 29724
rect 4160 29708 4212 29714
rect 4160 29650 4212 29656
rect 4066 29608 4122 29617
rect 4066 29543 4122 29552
rect 3516 29504 3568 29510
rect 3516 29446 3568 29452
rect 3528 29186 3556 29446
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3528 29158 3648 29186
rect 3620 29102 3648 29158
rect 3608 29096 3660 29102
rect 3436 29022 3556 29050
rect 3608 29038 3660 29044
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3436 28422 3464 28902
rect 3424 28416 3476 28422
rect 3424 28358 3476 28364
rect 3436 27674 3464 28358
rect 3424 27668 3476 27674
rect 3424 27610 3476 27616
rect 3528 27538 3556 29022
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3516 27532 3568 27538
rect 3516 27474 3568 27480
rect 3528 27130 3556 27474
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3988 26042 4016 26930
rect 4080 26858 4108 29543
rect 4172 29306 4200 29650
rect 4264 29646 4292 31418
rect 4252 29640 4304 29646
rect 4252 29582 4304 29588
rect 4160 29300 4212 29306
rect 4160 29242 4212 29248
rect 4252 29232 4304 29238
rect 4252 29174 4304 29180
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 4068 26240 4120 26246
rect 4068 26182 4120 26188
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 4080 25838 4108 26182
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 4080 25362 4108 25774
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 4080 24954 4108 25298
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 4172 24614 4200 25298
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 3344 24126 3464 24154
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 2792 21894 2820 22918
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2976 22030 3004 22374
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 2884 21350 2912 21422
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2884 20913 2912 21286
rect 2976 21146 3004 21966
rect 3252 21622 3280 22034
rect 3332 21956 3384 21962
rect 3332 21898 3384 21904
rect 3240 21616 3292 21622
rect 3240 21558 3292 21564
rect 3252 21146 3280 21558
rect 3344 21146 3372 21898
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 2870 20904 2926 20913
rect 2870 20839 2926 20848
rect 3436 17882 3464 24126
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 4068 22500 4120 22506
rect 4068 22442 4120 22448
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3976 21072 4028 21078
rect 3976 21014 4028 21020
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3988 20602 4016 21014
rect 4080 20942 4108 22442
rect 4172 22438 4200 24550
rect 4264 24274 4292 29174
rect 4356 28914 4384 34410
rect 4448 29617 4476 35119
rect 4896 34672 4948 34678
rect 4896 34614 4948 34620
rect 4908 34082 4936 34614
rect 5000 34202 5028 39520
rect 5172 35148 5224 35154
rect 5172 35090 5224 35096
rect 5184 34474 5212 35090
rect 5368 34649 5396 39520
rect 5736 36258 5764 39520
rect 5552 36230 5764 36258
rect 5552 35306 5580 36230
rect 5460 35290 5580 35306
rect 5448 35284 5580 35290
rect 5500 35278 5580 35284
rect 5448 35226 5500 35232
rect 5724 34944 5776 34950
rect 5724 34886 5776 34892
rect 5354 34640 5410 34649
rect 5354 34575 5410 34584
rect 5736 34542 5764 34886
rect 6196 34746 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6656 34746 6684 37726
rect 6932 35834 6960 39520
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 7392 35290 7420 39520
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 6736 35148 6788 35154
rect 6736 35090 6788 35096
rect 7472 35148 7524 35154
rect 7472 35090 7524 35096
rect 6184 34740 6236 34746
rect 6184 34682 6236 34688
rect 6644 34740 6696 34746
rect 6644 34682 6696 34688
rect 6748 34542 6776 35090
rect 7484 34746 7512 35090
rect 7472 34740 7524 34746
rect 7472 34682 7524 34688
rect 7484 34649 7512 34682
rect 6918 34640 6974 34649
rect 6918 34575 6974 34584
rect 7470 34640 7526 34649
rect 7470 34575 7526 34584
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 5172 34468 5224 34474
rect 5172 34410 5224 34416
rect 5264 34400 5316 34406
rect 5264 34342 5316 34348
rect 4988 34196 5040 34202
rect 4988 34138 5040 34144
rect 4908 34054 5028 34082
rect 4712 33312 4764 33318
rect 4712 33254 4764 33260
rect 4528 30796 4580 30802
rect 4528 30738 4580 30744
rect 4434 29608 4490 29617
rect 4434 29543 4490 29552
rect 4540 29306 4568 30738
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4632 29850 4660 30670
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4632 29073 4660 29582
rect 4618 29064 4674 29073
rect 4618 28999 4674 29008
rect 4356 28886 4476 28914
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4448 23322 4476 28886
rect 4632 28762 4660 28999
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 4528 27464 4580 27470
rect 4528 27406 4580 27412
rect 4540 27130 4568 27406
rect 4528 27124 4580 27130
rect 4528 27066 4580 27072
rect 4540 26586 4568 27066
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4528 26240 4580 26246
rect 4632 26228 4660 26726
rect 4580 26200 4660 26228
rect 4528 26182 4580 26188
rect 4540 24070 4568 26182
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4620 22704 4672 22710
rect 4620 22646 4672 22652
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4264 22250 4292 22578
rect 4172 22222 4292 22250
rect 4172 22166 4200 22222
rect 4160 22160 4212 22166
rect 4160 22102 4212 22108
rect 4172 21570 4200 22102
rect 4172 21542 4292 21570
rect 4264 21486 4292 21542
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4252 21480 4304 21486
rect 4252 21422 4304 21428
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 4080 20534 4108 20878
rect 4172 20874 4200 21286
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 4172 20602 4200 20810
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 4264 20466 4292 21422
rect 4434 21176 4490 21185
rect 4434 21111 4436 21120
rect 4488 21111 4490 21120
rect 4436 21082 4488 21088
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4448 20058 4476 21082
rect 4540 20942 4568 21490
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 4436 19712 4488 19718
rect 4540 19700 4568 20198
rect 4488 19672 4568 19700
rect 4436 19654 4488 19660
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3528 18426 3556 19178
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3988 17814 4016 19110
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2792 17338 2820 17682
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2884 16794 2912 17614
rect 3344 17270 3372 17614
rect 3424 17604 3476 17610
rect 3424 17546 3476 17552
rect 3332 17264 3384 17270
rect 3332 17206 3384 17212
rect 3436 16794 3464 17546
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 17202 3556 17478
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 4080 17202 4108 18362
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 4356 17202 4384 18090
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2884 16250 2912 16526
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2884 15910 2912 16186
rect 2976 16114 3004 16526
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 3252 15910 3280 16594
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3436 14618 3464 16730
rect 4080 16726 4108 17138
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4172 16794 4200 17002
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 4080 14618 4108 15846
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 2792 13530 2820 14418
rect 3252 14074 3280 14418
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3436 14006 3464 14554
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 3436 13870 3464 13942
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2884 12986 2912 13330
rect 3528 13190 3556 13738
rect 4080 13530 4108 14350
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 3528 12646 3556 13126
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 2976 12238 3004 12582
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 3252 12102 3280 12310
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3252 11762 3280 12038
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3606 11792 3662 11801
rect 3240 11756 3292 11762
rect 3606 11727 3662 11736
rect 3240 11698 3292 11704
rect 3620 11694 3648 11727
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3160 11393 3188 11494
rect 3146 11384 3202 11393
rect 3146 11319 3202 11328
rect 3528 11257 3556 11494
rect 3620 11354 3648 11630
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 2884 10062 2912 10610
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3344 10266 3372 10474
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10266 3464 10406
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 4080 9654 4108 10610
rect 4158 10160 4214 10169
rect 4158 10095 4214 10104
rect 4172 10062 4200 10095
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8974 2820 9318
rect 3436 9178 3464 9454
rect 4172 9382 4200 9998
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3436 9042 3464 9114
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2792 8362 2820 8910
rect 3436 8498 3464 8978
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3056 8424 3108 8430
rect 3054 8392 3056 8401
rect 3108 8392 3110 8401
rect 2780 8356 2832 8362
rect 3054 8327 3110 8336
rect 2780 8298 2832 8304
rect 2792 7818 2820 8298
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3712 8090 3740 8230
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2792 7002 2820 7754
rect 2976 7206 3004 7958
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7342 3372 7890
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 4080 7546 4108 7822
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3332 7336 3384 7342
rect 3330 7304 3332 7313
rect 3384 7304 3386 7313
rect 3330 7239 3386 7248
rect 2964 7200 3016 7206
rect 2962 7168 2964 7177
rect 3016 7168 3018 7177
rect 2962 7103 3018 7112
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2792 5778 2820 6831
rect 3344 6458 3372 7239
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3608 6384 3660 6390
rect 3606 6352 3608 6361
rect 3660 6352 3662 6361
rect 3606 6287 3662 6296
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2792 5370 2820 5714
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2148 2774 2268 2802
rect 2516 3862 2728 3890
rect 2148 480 2176 2774
rect 2410 2680 2466 2689
rect 2410 2615 2412 2624
rect 2464 2615 2466 2624
rect 2412 2586 2464 2592
rect 2516 1057 2544 3862
rect 2792 3754 2820 4626
rect 2872 4616 2924 4622
rect 2870 4584 2872 4593
rect 2924 4584 2926 4593
rect 2870 4519 2926 4528
rect 3160 4185 3188 6054
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3528 4826 3556 5102
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3146 4176 3202 4185
rect 3146 4111 3202 4120
rect 3148 4072 3200 4078
rect 3252 4060 3280 4762
rect 3988 4622 4016 5034
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3988 4282 4016 4558
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3330 4176 3386 4185
rect 3330 4111 3386 4120
rect 3344 4078 3372 4111
rect 3200 4032 3280 4060
rect 3148 4014 3200 4020
rect 2700 3738 2820 3754
rect 3252 3738 3280 4032
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 2688 3732 2820 3738
rect 2740 3726 2820 3732
rect 3240 3732 3292 3738
rect 2688 3674 2740 3680
rect 3240 3674 3292 3680
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2700 2825 2728 3470
rect 2884 3194 2912 3470
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3252 2990 3280 3674
rect 3344 3534 3372 4014
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 2686 2816 2742 2825
rect 2686 2751 2742 2760
rect 3344 2650 3372 3470
rect 3436 2650 3464 3538
rect 4172 3398 4200 9318
rect 4264 7478 4292 16934
rect 4356 16590 4384 17138
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 14482 4384 16526
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4448 13297 4476 19654
rect 4528 17060 4580 17066
rect 4528 17002 4580 17008
rect 4540 16794 4568 17002
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4540 16250 4568 16730
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4528 13456 4580 13462
rect 4526 13424 4528 13433
rect 4580 13424 4582 13433
rect 4526 13359 4582 13368
rect 4434 13288 4490 13297
rect 4434 13223 4490 13232
rect 4540 12986 4568 13359
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 8090 4568 12650
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4252 7472 4304 7478
rect 4356 7449 4384 7890
rect 4632 7562 4660 22646
rect 4724 16017 4752 33254
rect 4896 32292 4948 32298
rect 4896 32234 4948 32240
rect 4908 30734 4936 32234
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4804 30116 4856 30122
rect 4804 30058 4856 30064
rect 4816 29646 4844 30058
rect 4908 30054 4936 30670
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4908 29170 4936 29990
rect 5000 29617 5028 34054
rect 5080 31952 5132 31958
rect 5080 31894 5132 31900
rect 5092 31482 5120 31894
rect 5080 31476 5132 31482
rect 5080 31418 5132 31424
rect 4986 29608 5042 29617
rect 4986 29543 5042 29552
rect 4896 29164 4948 29170
rect 4896 29106 4948 29112
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4816 28404 4844 29038
rect 5000 28506 5028 29543
rect 5172 29504 5224 29510
rect 5172 29446 5224 29452
rect 5184 29102 5212 29446
rect 5276 29238 5304 34342
rect 5448 34060 5500 34066
rect 5448 34002 5500 34008
rect 5460 33318 5488 34002
rect 5448 33312 5500 33318
rect 5500 33272 5580 33300
rect 5448 33254 5500 33260
rect 5356 32224 5408 32230
rect 5356 32166 5408 32172
rect 5368 31958 5396 32166
rect 5356 31952 5408 31958
rect 5356 31894 5408 31900
rect 5448 31952 5500 31958
rect 5448 31894 5500 31900
rect 5460 31142 5488 31894
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5460 30326 5488 31078
rect 5448 30320 5500 30326
rect 5448 30262 5500 30268
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5264 29232 5316 29238
rect 5264 29174 5316 29180
rect 5368 29170 5396 29582
rect 5552 29170 5580 33272
rect 5736 29714 5764 34478
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6644 34060 6696 34066
rect 6644 34002 6696 34008
rect 6090 33416 6146 33425
rect 6090 33351 6146 33360
rect 5814 33144 5870 33153
rect 5814 33079 5870 33088
rect 5828 32978 5856 33079
rect 5816 32972 5868 32978
rect 5816 32914 5868 32920
rect 5828 32502 5856 32914
rect 5816 32496 5868 32502
rect 5816 32438 5868 32444
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5828 29345 5856 32438
rect 5908 32020 5960 32026
rect 5908 31962 5960 31968
rect 5814 29336 5870 29345
rect 5814 29271 5870 29280
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 5540 29164 5592 29170
rect 5540 29106 5592 29112
rect 5172 29096 5224 29102
rect 5172 29038 5224 29044
rect 5184 28762 5212 29038
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 5000 28478 5304 28506
rect 5172 28416 5224 28422
rect 4816 28376 5120 28404
rect 5092 27169 5120 28376
rect 5172 28358 5224 28364
rect 5184 27470 5212 28358
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 5078 27160 5134 27169
rect 5078 27095 5134 27104
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 5000 24721 5028 26794
rect 4986 24712 5042 24721
rect 4986 24647 5042 24656
rect 4896 23316 4948 23322
rect 4896 23258 4948 23264
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4816 21146 4844 22918
rect 4908 22778 4936 23258
rect 4896 22772 4948 22778
rect 4896 22714 4948 22720
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 4802 20904 4858 20913
rect 4802 20839 4858 20848
rect 4816 16794 4844 20839
rect 4908 17338 4936 22714
rect 5000 21350 5028 24647
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 4986 20360 5042 20369
rect 4986 20295 5042 20304
rect 5000 20262 5028 20295
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4908 17134 4936 17274
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4816 16182 4844 16730
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4710 16008 4766 16017
rect 4710 15943 4766 15952
rect 4724 14618 4752 15943
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4724 14074 4752 14554
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4724 12646 4752 13330
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12481 4752 12582
rect 4710 12472 4766 12481
rect 4710 12407 4766 12416
rect 4816 12186 4844 16118
rect 4448 7534 4660 7562
rect 4724 12158 4844 12186
rect 4252 7414 4304 7420
rect 4342 7440 4398 7449
rect 4342 7375 4398 7384
rect 4356 7206 4384 7375
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4356 5778 4384 7142
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4250 5672 4306 5681
rect 4250 5607 4252 5616
rect 4304 5607 4306 5616
rect 4252 5578 4304 5584
rect 4356 4826 4384 5714
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 4250 3224 4306 3233
rect 4250 3159 4306 3168
rect 3974 3088 4030 3097
rect 3974 3023 4030 3032
rect 3514 2952 3570 2961
rect 3514 2887 3570 2896
rect 3528 2854 3556 2887
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2594 1456 2650 1465
rect 2594 1391 2650 1400
rect 2502 1048 2558 1057
rect 2502 983 2558 992
rect 2608 480 2636 1391
rect 2976 480 3004 2314
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 480 3372 2246
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3988 1442 4016 3023
rect 3804 1414 4016 1442
rect 3804 480 3832 1414
rect 4264 1034 4292 3159
rect 4448 2922 4476 7534
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 5166 4568 7142
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4540 4826 4568 5102
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4526 3496 4582 3505
rect 4526 3431 4582 3440
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4342 2816 4398 2825
rect 4342 2751 4398 2760
rect 4356 2582 4384 2751
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4172 1006 4292 1034
rect 4172 480 4200 1006
rect 4540 480 4568 3431
rect 4632 2446 4660 7414
rect 4724 6866 4752 12158
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4816 11762 4844 12038
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4908 11234 4936 17070
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 16250 5028 16526
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5000 14074 5028 14350
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5092 12714 5120 27095
rect 5170 25664 5226 25673
rect 5170 25599 5226 25608
rect 5184 24954 5212 25599
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 21690 5212 22374
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5276 20330 5304 28478
rect 5368 28422 5396 29106
rect 5448 28688 5500 28694
rect 5828 28665 5856 29271
rect 5920 28762 5948 31962
rect 6000 30592 6052 30598
rect 6000 30534 6052 30540
rect 6012 30190 6040 30534
rect 6000 30184 6052 30190
rect 6000 30126 6052 30132
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 6012 29034 6040 29650
rect 6104 29102 6132 33351
rect 6656 33318 6684 34002
rect 6644 33312 6696 33318
rect 6644 33254 6696 33260
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6644 31204 6696 31210
rect 6644 31146 6696 31152
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6656 30666 6684 31146
rect 6748 30977 6776 34478
rect 6932 34202 6960 34575
rect 7196 34536 7248 34542
rect 7196 34478 7248 34484
rect 6920 34196 6972 34202
rect 6920 34138 6972 34144
rect 6828 33856 6880 33862
rect 6828 33798 6880 33804
rect 6840 33522 6868 33798
rect 6828 33516 6880 33522
rect 6828 33458 6880 33464
rect 6826 33144 6882 33153
rect 6826 33079 6828 33088
rect 6880 33079 6882 33088
rect 6828 33050 6880 33056
rect 6840 32570 6868 33050
rect 6918 33008 6974 33017
rect 6918 32943 6974 32952
rect 6828 32564 6880 32570
rect 6828 32506 6880 32512
rect 6932 32366 6960 32943
rect 7012 32768 7064 32774
rect 7012 32710 7064 32716
rect 6920 32360 6972 32366
rect 6920 32302 6972 32308
rect 6828 32224 6880 32230
rect 6828 32166 6880 32172
rect 6840 31958 6868 32166
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6840 31482 6868 31894
rect 6932 31890 6960 32302
rect 7024 31890 7052 32710
rect 7208 32348 7236 34478
rect 7760 34202 7788 39520
rect 8220 35578 8248 39520
rect 8482 35864 8538 35873
rect 8482 35799 8484 35808
rect 8536 35799 8538 35808
rect 8484 35770 8536 35776
rect 7852 35550 8248 35578
rect 7748 34196 7800 34202
rect 7748 34138 7800 34144
rect 7564 34060 7616 34066
rect 7564 34002 7616 34008
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7288 33312 7340 33318
rect 7288 33254 7340 33260
rect 7116 32320 7236 32348
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 7012 31884 7064 31890
rect 7012 31826 7064 31832
rect 6932 31793 6960 31826
rect 6918 31784 6974 31793
rect 6918 31719 6974 31728
rect 7024 31482 7052 31826
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 7116 31362 7144 32320
rect 7300 32178 7328 33254
rect 7392 32910 7420 33322
rect 7576 33114 7604 34002
rect 7852 33153 7880 35550
rect 8024 35488 8076 35494
rect 8024 35430 8076 35436
rect 7932 34536 7984 34542
rect 7932 34478 7984 34484
rect 7944 33862 7972 34478
rect 7932 33856 7984 33862
rect 7932 33798 7984 33804
rect 7838 33144 7894 33153
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7760 33102 7838 33130
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7392 32434 7420 32846
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7470 32328 7526 32337
rect 7380 32292 7432 32298
rect 7470 32263 7526 32272
rect 7380 32234 7432 32240
rect 6932 31334 7144 31362
rect 7208 32150 7328 32178
rect 6734 30968 6790 30977
rect 6734 30903 6790 30912
rect 6644 30660 6696 30666
rect 6644 30602 6696 30608
rect 6184 30252 6236 30258
rect 6184 30194 6236 30200
rect 6092 29096 6144 29102
rect 6092 29038 6144 29044
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 5908 28756 5960 28762
rect 5908 28698 5960 28704
rect 5448 28630 5500 28636
rect 5814 28656 5870 28665
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5460 28218 5488 28630
rect 5814 28591 5870 28600
rect 5816 28552 5868 28558
rect 5816 28494 5868 28500
rect 5632 28416 5684 28422
rect 5632 28358 5684 28364
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5460 26790 5488 27406
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5460 26042 5488 26726
rect 5448 26036 5500 26042
rect 5448 25978 5500 25984
rect 5448 25832 5500 25838
rect 5448 25774 5500 25780
rect 5460 25498 5488 25774
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5552 23225 5580 27474
rect 5644 24818 5672 28358
rect 5828 28218 5856 28494
rect 5920 28218 5948 28698
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 5908 28212 5960 28218
rect 5908 28154 5960 28160
rect 5828 26586 5856 28154
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5644 24410 5672 24754
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5644 23526 5672 24142
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5538 23216 5594 23225
rect 5538 23151 5594 23160
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5368 22778 5396 23054
rect 5816 22976 5868 22982
rect 5816 22918 5868 22924
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5828 22642 5856 22918
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 5540 22568 5592 22574
rect 5538 22536 5540 22545
rect 5592 22536 5594 22545
rect 5538 22471 5594 22480
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5460 21554 5488 21830
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5264 20324 5316 20330
rect 5264 20266 5316 20272
rect 5368 18737 5396 21286
rect 5644 21010 5672 21966
rect 5920 21894 5948 22374
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 6012 21298 6040 28970
rect 5736 21270 6040 21298
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5644 20602 5672 20946
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5630 18864 5686 18873
rect 5630 18799 5686 18808
rect 5354 18728 5410 18737
rect 5354 18663 5410 18672
rect 5368 18426 5396 18663
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5368 18222 5396 18362
rect 5356 18216 5408 18222
rect 5552 18193 5580 18566
rect 5356 18158 5408 18164
rect 5538 18184 5594 18193
rect 5538 18119 5540 18128
rect 5592 18119 5594 18128
rect 5540 18090 5592 18096
rect 5448 18080 5500 18086
rect 5500 18028 5580 18034
rect 5448 18022 5580 18028
rect 5460 18006 5580 18022
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5184 15502 5212 17818
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16153 5488 16934
rect 5552 16794 5580 18006
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5446 16144 5502 16153
rect 5552 16114 5580 16730
rect 5446 16079 5502 16088
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12850 5212 13126
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5000 12102 5028 12582
rect 5184 12442 5212 12786
rect 5460 12782 5488 15846
rect 5644 15450 5672 18799
rect 5552 15422 5672 15450
rect 5552 14550 5580 15422
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5644 14618 5672 15302
rect 5736 15201 5764 21270
rect 6000 21072 6052 21078
rect 6000 21014 6052 21020
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5828 19938 5856 20266
rect 6012 20262 6040 21014
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6012 19990 6040 20198
rect 6000 19984 6052 19990
rect 5828 19910 5948 19938
rect 6000 19926 6052 19932
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 15978 5856 18566
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5920 15688 5948 19910
rect 6012 19514 6040 19926
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18902 6040 19110
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 18290 6040 18702
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 6012 17542 6040 18226
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 6012 16726 6040 17478
rect 6104 17270 6132 29038
rect 6196 27606 6224 30194
rect 6644 30184 6696 30190
rect 6644 30126 6696 30132
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 6288 29238 6316 29650
rect 6276 29232 6328 29238
rect 6274 29200 6276 29209
rect 6328 29200 6330 29209
rect 6274 29135 6330 29144
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6184 27600 6236 27606
rect 6184 27542 6236 27548
rect 6656 27402 6684 30126
rect 6828 28960 6880 28966
rect 6828 28902 6880 28908
rect 6840 28694 6868 28902
rect 6828 28688 6880 28694
rect 6828 28630 6880 28636
rect 6734 27568 6790 27577
rect 6734 27503 6736 27512
rect 6788 27503 6790 27512
rect 6736 27474 6788 27480
rect 6644 27396 6696 27402
rect 6644 27338 6696 27344
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6196 24954 6224 26522
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6656 25498 6684 27338
rect 6748 27130 6776 27474
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6736 26240 6788 26246
rect 6736 26182 6788 26188
rect 6644 25492 6696 25498
rect 6644 25434 6696 25440
rect 6748 25158 6776 26182
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6184 24948 6236 24954
rect 6184 24890 6236 24896
rect 6196 24342 6224 24890
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6184 24336 6236 24342
rect 6184 24278 6236 24284
rect 6196 23866 6224 24278
rect 6644 24268 6696 24274
rect 6644 24210 6696 24216
rect 6184 23860 6236 23866
rect 6184 23802 6236 23808
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6182 23216 6238 23225
rect 6182 23151 6238 23160
rect 6196 18970 6224 23151
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 6288 21690 6316 22034
rect 6276 21684 6328 21690
rect 6276 21626 6328 21632
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6366 19952 6422 19961
rect 6276 19916 6328 19922
rect 6366 19887 6368 19896
rect 6276 19858 6328 19864
rect 6420 19887 6422 19896
rect 6368 19858 6420 19864
rect 6288 19242 6316 19858
rect 6380 19310 6408 19858
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 6276 19236 6328 19242
rect 6276 19178 6328 19184
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6196 18426 6224 18906
rect 6552 18896 6604 18902
rect 6656 18873 6684 24210
rect 6748 23526 6776 25094
rect 6840 24698 6868 26726
rect 6932 25838 6960 31334
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7012 30728 7064 30734
rect 7116 30705 7144 30738
rect 7012 30670 7064 30676
rect 7102 30696 7158 30705
rect 7024 30394 7052 30670
rect 7102 30631 7158 30640
rect 7012 30388 7064 30394
rect 7012 30330 7064 30336
rect 7116 30138 7144 30631
rect 7024 30110 7144 30138
rect 7024 29782 7052 30110
rect 7104 30048 7156 30054
rect 7104 29990 7156 29996
rect 7116 29850 7144 29990
rect 7104 29844 7156 29850
rect 7104 29786 7156 29792
rect 7012 29776 7064 29782
rect 7208 29730 7236 32150
rect 7392 31822 7420 32234
rect 7380 31816 7432 31822
rect 7380 31758 7432 31764
rect 7484 31634 7512 32263
rect 7576 32201 7604 33050
rect 7562 32192 7618 32201
rect 7562 32127 7618 32136
rect 7760 32065 7788 33102
rect 7838 33079 7894 33088
rect 7932 32768 7984 32774
rect 7932 32710 7984 32716
rect 7840 32428 7892 32434
rect 7840 32370 7892 32376
rect 7852 32230 7880 32370
rect 7840 32224 7892 32230
rect 7840 32166 7892 32172
rect 7746 32056 7802 32065
rect 7746 31991 7802 32000
rect 7852 31754 7880 32166
rect 7840 31748 7892 31754
rect 7840 31690 7892 31696
rect 7392 31606 7512 31634
rect 7288 29844 7340 29850
rect 7288 29786 7340 29792
rect 7012 29718 7064 29724
rect 7116 29702 7236 29730
rect 7010 27976 7066 27985
rect 7010 27911 7066 27920
rect 7024 27878 7052 27911
rect 7012 27872 7064 27878
rect 7012 27814 7064 27820
rect 7116 26042 7144 29702
rect 7196 29504 7248 29510
rect 7196 29446 7248 29452
rect 7208 29170 7236 29446
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7208 27130 7236 28698
rect 7300 28694 7328 29786
rect 7288 28688 7340 28694
rect 7288 28630 7340 28636
rect 7196 27124 7248 27130
rect 7196 27066 7248 27072
rect 7300 26976 7328 28630
rect 7392 27962 7420 31606
rect 7472 31476 7524 31482
rect 7472 31418 7524 31424
rect 7484 29170 7512 31418
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7564 31136 7616 31142
rect 7564 31078 7616 31084
rect 7576 30841 7604 31078
rect 7668 30870 7696 31282
rect 7656 30864 7708 30870
rect 7562 30832 7618 30841
rect 7656 30806 7708 30812
rect 7562 30767 7618 30776
rect 7564 30048 7616 30054
rect 7564 29990 7616 29996
rect 7472 29164 7524 29170
rect 7472 29106 7524 29112
rect 7484 28762 7512 29106
rect 7472 28756 7524 28762
rect 7472 28698 7524 28704
rect 7576 28218 7604 29990
rect 7654 29880 7710 29889
rect 7654 29815 7656 29824
rect 7708 29815 7710 29824
rect 7656 29786 7708 29792
rect 7852 29646 7880 31690
rect 7944 31278 7972 32710
rect 7932 31272 7984 31278
rect 7932 31214 7984 31220
rect 7656 29640 7708 29646
rect 7654 29608 7656 29617
rect 7840 29640 7892 29646
rect 7708 29608 7710 29617
rect 7840 29582 7892 29588
rect 7654 29543 7710 29552
rect 7668 29306 7696 29543
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7564 28212 7616 28218
rect 7564 28154 7616 28160
rect 7392 27934 7604 27962
rect 7380 27872 7432 27878
rect 7380 27814 7432 27820
rect 7392 27674 7420 27814
rect 7380 27668 7432 27674
rect 7380 27610 7432 27616
rect 7208 26948 7328 26976
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 6920 25696 6972 25702
rect 6920 25638 6972 25644
rect 6932 24818 6960 25638
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 7024 24954 7052 25298
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6840 24682 6960 24698
rect 6840 24676 6972 24682
rect 6840 24670 6920 24676
rect 6920 24618 6972 24624
rect 6932 24410 6960 24618
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 7024 24138 7052 24890
rect 7102 24576 7158 24585
rect 7102 24511 7158 24520
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6748 22098 6776 23462
rect 7116 22658 7144 24511
rect 7208 22778 7236 26948
rect 7286 26888 7342 26897
rect 7286 26823 7288 26832
rect 7340 26823 7342 26832
rect 7288 26794 7340 26800
rect 7286 25800 7342 25809
rect 7286 25735 7288 25744
rect 7340 25735 7342 25744
rect 7288 25706 7340 25712
rect 7286 24848 7342 24857
rect 7286 24783 7342 24792
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 6920 22636 6972 22642
rect 7116 22630 7236 22658
rect 6920 22578 6972 22584
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 20058 6776 21830
rect 6932 21146 6960 22578
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6840 20058 6868 20402
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 7010 19272 7066 19281
rect 7010 19207 7066 19216
rect 6828 19168 6880 19174
rect 7024 19156 7052 19207
rect 6880 19128 7052 19156
rect 6828 19110 6880 19116
rect 6552 18838 6604 18844
rect 6642 18864 6698 18873
rect 6564 18714 6592 18838
rect 6642 18799 6698 18808
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6564 18686 6684 18714
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16794 6132 16934
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6092 16788 6144 16794
rect 6656 16776 6684 18686
rect 6748 18086 6776 18770
rect 6736 18080 6788 18086
rect 6734 18048 6736 18057
rect 6788 18048 6790 18057
rect 6734 17983 6790 17992
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6092 16730 6144 16736
rect 6564 16748 6684 16776
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 6012 16114 6040 16390
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6012 15706 6040 16050
rect 6196 15910 6224 16662
rect 6564 16250 6592 16748
rect 6642 16552 6698 16561
rect 6642 16487 6698 16496
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 5828 15660 5948 15688
rect 6000 15700 6052 15706
rect 5722 15192 5778 15201
rect 5722 15127 5778 15136
rect 5828 14634 5856 15660
rect 6000 15642 6052 15648
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5920 15162 5948 15506
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5736 14606 5856 14634
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5552 12714 5580 14214
rect 5644 13530 5672 14554
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5448 12640 5500 12646
rect 5736 12594 5764 14606
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5828 14074 5856 14486
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5920 13274 5948 15098
rect 6012 14396 6040 15642
rect 6196 15502 6224 15846
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6104 14958 6132 15438
rect 6380 15162 6408 15438
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6092 14408 6144 14414
rect 6012 14368 6092 14396
rect 6092 14350 6144 14356
rect 6104 14074 6132 14350
rect 6092 14068 6144 14074
rect 6144 14028 6224 14056
rect 6092 14010 6144 14016
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6104 13530 6132 13738
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5816 13252 5868 13258
rect 5920 13246 6132 13274
rect 5816 13194 5868 13200
rect 5448 12582 5500 12588
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5092 11354 5120 12242
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5184 12102 5212 12174
rect 5460 12102 5488 12582
rect 5552 12566 5764 12594
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5184 11354 5212 12038
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 4908 11206 5028 11234
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4816 9994 4844 10542
rect 4908 10470 4936 11086
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4816 8974 4844 9930
rect 4908 9178 4936 10406
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8650 4844 8910
rect 4816 8634 4936 8650
rect 4816 8628 4948 8634
rect 4816 8622 4896 8628
rect 4896 8570 4948 8576
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4816 7886 4844 8298
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7342 4844 7822
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4712 6248 4764 6254
rect 4710 6216 4712 6225
rect 4764 6216 4766 6225
rect 4710 6151 4766 6160
rect 4816 5370 4844 7278
rect 5000 6474 5028 11206
rect 5092 9654 5120 11290
rect 5170 11248 5226 11257
rect 5170 11183 5226 11192
rect 5184 10266 5212 11183
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5092 7546 5120 9590
rect 5184 9518 5212 10202
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5184 9217 5212 9454
rect 5170 9208 5226 9217
rect 5276 9178 5304 9454
rect 5368 9194 5396 11630
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5460 11354 5488 11562
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 9738 5580 12566
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5644 11150 5672 12378
rect 5724 12368 5776 12374
rect 5828 12345 5856 13194
rect 5724 12310 5776 12316
rect 5814 12336 5870 12345
rect 5736 11898 5764 12310
rect 5814 12271 5870 12280
rect 6104 12186 6132 13246
rect 6196 12374 6224 14028
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6472 12714 6500 13398
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6104 12158 6224 12186
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 10810 5672 11086
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5460 9710 5580 9738
rect 5460 9330 5488 9710
rect 5644 9636 5672 10746
rect 5736 10742 5764 11834
rect 5906 11384 5962 11393
rect 5906 11319 5908 11328
rect 5960 11319 5962 11328
rect 5908 11290 5960 11296
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 10810 5856 11154
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5828 9994 5856 10746
rect 5920 10266 5948 11290
rect 5998 11248 6054 11257
rect 5998 11183 6054 11192
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5644 9608 5764 9636
rect 5460 9302 5672 9330
rect 5368 9178 5580 9194
rect 5170 9143 5226 9152
rect 5264 9172 5316 9178
rect 5368 9172 5592 9178
rect 5368 9166 5540 9172
rect 5264 9114 5316 9120
rect 5540 9114 5592 9120
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5184 8090 5212 8978
rect 5644 8956 5672 9302
rect 5736 9110 5764 9608
rect 5906 9344 5962 9353
rect 5906 9279 5962 9288
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5644 8928 5856 8956
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5092 7342 5120 7482
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5184 7206 5212 8026
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5630 7168 5686 7177
rect 5630 7103 5686 7112
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 4908 6446 5028 6474
rect 5184 6458 5212 6802
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5172 6452 5224 6458
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4724 3369 4752 3538
rect 4710 3360 4766 3369
rect 4710 3295 4766 3304
rect 4724 3126 4752 3295
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4908 3058 4936 6446
rect 5172 6394 5224 6400
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5000 480 5028 6326
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5092 4010 5120 4626
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5092 3670 5120 3946
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 2689 5120 3334
rect 5078 2680 5134 2689
rect 5184 2650 5212 6394
rect 5262 5672 5318 5681
rect 5262 5607 5318 5616
rect 5276 3346 5304 5607
rect 5354 4448 5410 4457
rect 5354 4383 5410 4392
rect 5368 3466 5396 4383
rect 5460 3618 5488 6598
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 4690 5580 5510
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5644 4321 5672 7103
rect 5828 6780 5856 8928
rect 5920 6905 5948 9279
rect 5906 6896 5962 6905
rect 5906 6831 5962 6840
rect 5828 6752 5948 6780
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5722 5128 5778 5137
rect 5722 5063 5724 5072
rect 5776 5063 5778 5072
rect 5724 5034 5776 5040
rect 5630 4312 5686 4321
rect 5630 4247 5686 4256
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3777 5764 3878
rect 5722 3768 5778 3777
rect 5722 3703 5778 3712
rect 5460 3590 5764 3618
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5276 3318 5396 3346
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5078 2615 5134 2624
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5276 2009 5304 2926
rect 5262 2000 5318 2009
rect 5262 1935 5318 1944
rect 5368 480 5396 3318
rect 5460 3058 5488 3470
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5460 2446 5488 2994
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5736 480 5764 3590
rect 5828 610 5856 6054
rect 5920 5778 5948 6752
rect 6012 6390 6040 11183
rect 6196 11098 6224 12158
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6104 11070 6224 11098
rect 6104 9353 6132 11070
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6196 10538 6224 10950
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6196 10198 6224 10474
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6196 9722 6224 10134
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6090 9344 6146 9353
rect 6090 9279 6146 9288
rect 6196 9160 6224 9658
rect 6460 9648 6512 9654
rect 6458 9616 6460 9625
rect 6512 9616 6514 9625
rect 6458 9551 6514 9560
rect 6656 9518 6684 16487
rect 6748 11014 6776 17206
rect 6840 16794 6868 17614
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6840 16538 6868 16730
rect 6840 16510 6960 16538
rect 6932 16250 6960 16510
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6840 14385 6868 16186
rect 6826 14376 6882 14385
rect 6826 14311 6882 14320
rect 6840 13818 6868 14311
rect 6932 13938 6960 16186
rect 7024 14906 7052 19128
rect 7116 18970 7144 20266
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7104 18352 7156 18358
rect 7102 18320 7104 18329
rect 7156 18320 7158 18329
rect 7102 18255 7158 18264
rect 7102 14920 7158 14929
rect 7024 14878 7102 14906
rect 7102 14855 7158 14864
rect 7116 14362 7144 14855
rect 7208 14482 7236 22630
rect 7300 15570 7328 24783
rect 7392 22778 7420 27610
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 7484 26586 7512 26930
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7484 25906 7512 26522
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 7484 25430 7512 25842
rect 7472 25424 7524 25430
rect 7472 25366 7524 25372
rect 7576 25265 7604 27934
rect 7562 25256 7618 25265
rect 7562 25191 7618 25200
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7484 24342 7512 24754
rect 7472 24336 7524 24342
rect 7472 24278 7524 24284
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7668 22642 7696 22918
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7392 21554 7420 22034
rect 7668 21690 7696 22578
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7470 20496 7526 20505
rect 7470 20431 7526 20440
rect 7484 18170 7512 20431
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7576 18290 7604 18566
rect 7668 18290 7696 18906
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7484 18142 7604 18170
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7392 17202 7420 17682
rect 7484 17542 7512 18022
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7484 17338 7512 17478
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7576 14634 7604 18142
rect 7668 17882 7696 18226
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7760 17649 7788 28970
rect 7852 28762 7880 29582
rect 7840 28756 7892 28762
rect 7840 28698 7892 28704
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7852 24585 7880 28154
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 7944 26790 7972 27474
rect 8036 26874 8064 35430
rect 8116 34944 8168 34950
rect 8116 34886 8168 34892
rect 8128 34474 8156 34886
rect 8300 34740 8352 34746
rect 8220 34700 8300 34728
rect 8116 34468 8168 34474
rect 8116 34410 8168 34416
rect 8220 34354 8248 34700
rect 8300 34682 8352 34688
rect 8588 34626 8616 39520
rect 8956 37210 8984 39520
rect 8772 37182 8984 37210
rect 8496 34598 8616 34626
rect 8666 34640 8722 34649
rect 8496 34513 8524 34598
rect 8666 34575 8722 34584
rect 8482 34504 8538 34513
rect 8482 34439 8538 34448
rect 8576 34468 8628 34474
rect 8576 34410 8628 34416
rect 8128 34326 8248 34354
rect 8128 31346 8156 34326
rect 8300 33856 8352 33862
rect 8300 33798 8352 33804
rect 8208 33312 8260 33318
rect 8208 33254 8260 33260
rect 8220 31754 8248 33254
rect 8208 31748 8260 31754
rect 8208 31690 8260 31696
rect 8220 31482 8248 31690
rect 8208 31476 8260 31482
rect 8208 31418 8260 31424
rect 8116 31340 8168 31346
rect 8116 31282 8168 31288
rect 8206 30968 8262 30977
rect 8206 30903 8262 30912
rect 8220 30802 8248 30903
rect 8208 30796 8260 30802
rect 8208 30738 8260 30744
rect 8220 30054 8248 30738
rect 8312 30190 8340 33798
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 8404 32026 8432 32914
rect 8588 32910 8616 34410
rect 8484 32904 8536 32910
rect 8484 32846 8536 32852
rect 8576 32904 8628 32910
rect 8576 32846 8628 32852
rect 8496 32570 8524 32846
rect 8484 32564 8536 32570
rect 8484 32506 8536 32512
rect 8484 32292 8536 32298
rect 8484 32234 8536 32240
rect 8392 32020 8444 32026
rect 8392 31962 8444 31968
rect 8404 31482 8432 31962
rect 8392 31476 8444 31482
rect 8392 31418 8444 31424
rect 8496 30938 8524 32234
rect 8588 31668 8616 32846
rect 8680 32502 8708 34575
rect 8668 32496 8720 32502
rect 8668 32438 8720 32444
rect 8772 32298 8800 37182
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 9310 34504 9366 34513
rect 9310 34439 9366 34448
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9324 32858 9352 34439
rect 9416 32994 9444 39520
rect 9678 34776 9734 34785
rect 9678 34711 9734 34720
rect 9692 33425 9720 34711
rect 9678 33416 9734 33425
rect 9678 33351 9734 33360
rect 9416 32966 9720 32994
rect 9324 32830 9628 32858
rect 9404 32768 9456 32774
rect 9404 32710 9456 32716
rect 9494 32736 9550 32745
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8850 32464 8906 32473
rect 9416 32434 9444 32710
rect 9494 32671 9550 32680
rect 9508 32434 9536 32671
rect 8850 32399 8906 32408
rect 9404 32428 9456 32434
rect 8760 32292 8812 32298
rect 8760 32234 8812 32240
rect 8666 32192 8722 32201
rect 8666 32127 8722 32136
rect 8680 31906 8708 32127
rect 8680 31878 8800 31906
rect 8668 31680 8720 31686
rect 8588 31640 8668 31668
rect 8668 31622 8720 31628
rect 8576 31136 8628 31142
rect 8576 31078 8628 31084
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8208 30048 8260 30054
rect 8208 29990 8260 29996
rect 8312 29850 8340 30126
rect 8300 29844 8352 29850
rect 8300 29786 8352 29792
rect 8496 29714 8524 30874
rect 8588 30734 8616 31078
rect 8576 30728 8628 30734
rect 8576 30670 8628 30676
rect 8588 30122 8616 30670
rect 8680 30326 8708 31622
rect 8668 30320 8720 30326
rect 8668 30262 8720 30268
rect 8576 30116 8628 30122
rect 8576 30058 8628 30064
rect 8484 29708 8536 29714
rect 8484 29650 8536 29656
rect 8666 29336 8722 29345
rect 8666 29271 8668 29280
rect 8720 29271 8722 29280
rect 8668 29242 8720 29248
rect 8390 29200 8446 29209
rect 8390 29135 8446 29144
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8116 27872 8168 27878
rect 8114 27840 8116 27849
rect 8168 27840 8170 27849
rect 8114 27775 8170 27784
rect 8312 27577 8340 28358
rect 8298 27568 8354 27577
rect 8298 27503 8354 27512
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 8036 26846 8156 26874
rect 7932 26784 7984 26790
rect 7930 26752 7932 26761
rect 7984 26752 7986 26761
rect 7930 26687 7986 26696
rect 7838 24576 7894 24585
rect 7838 24511 7894 24520
rect 7944 22710 7972 26687
rect 8024 26036 8076 26042
rect 8024 25978 8076 25984
rect 7932 22704 7984 22710
rect 7932 22646 7984 22652
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7944 22273 7972 22374
rect 7930 22264 7986 22273
rect 7930 22199 7986 22208
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7746 17640 7802 17649
rect 7746 17575 7802 17584
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7760 15706 7788 15982
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7760 14906 7788 15642
rect 7852 15065 7880 19178
rect 7838 15056 7894 15065
rect 7838 14991 7894 15000
rect 7760 14878 7880 14906
rect 7748 14816 7800 14822
rect 7746 14784 7748 14793
rect 7800 14784 7802 14793
rect 7746 14719 7802 14728
rect 7576 14606 7788 14634
rect 7656 14544 7708 14550
rect 7576 14492 7656 14498
rect 7576 14486 7708 14492
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7576 14470 7696 14486
rect 7472 14408 7524 14414
rect 7194 14376 7250 14385
rect 7012 14340 7064 14346
rect 7116 14334 7194 14362
rect 7472 14350 7524 14356
rect 7194 14311 7250 14320
rect 7012 14282 7064 14288
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 7024 13870 7052 14282
rect 7012 13864 7064 13870
rect 6840 13790 6960 13818
rect 7012 13806 7064 13812
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6748 10062 6776 10678
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10266 6868 10406
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6932 9654 6960 13790
rect 7208 13716 7236 14311
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7024 13688 7236 13716
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6104 9132 6224 9160
rect 6104 6866 6132 9132
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8634 6224 8978
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6656 8090 6684 9454
rect 7024 9450 7052 13688
rect 7300 13512 7328 14214
rect 7116 13484 7328 13512
rect 7116 12442 7144 13484
rect 7484 13462 7512 14350
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7208 12442 7236 13330
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7300 12986 7328 13262
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7116 11694 7144 12378
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7116 11082 7144 11494
rect 7208 11354 7236 12378
rect 7300 11898 7328 12922
rect 7484 12918 7512 13262
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6748 8634 6776 9114
rect 7024 9110 7052 9386
rect 7116 9178 7144 11018
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6840 7886 6868 8366
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7546 6868 7822
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6104 6458 6132 6802
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 6090 6080 6146 6089
rect 6090 6015 6146 6024
rect 6104 5914 6132 6015
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5920 5137 5948 5714
rect 6104 5370 6132 5850
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5160 6052 5166
rect 5906 5128 5962 5137
rect 6000 5102 6052 5108
rect 5906 5063 5962 5072
rect 6012 4758 6040 5102
rect 6000 4752 6052 4758
rect 6104 4729 6132 5306
rect 6000 4694 6052 4700
rect 6090 4720 6146 4729
rect 6012 4146 6040 4694
rect 6090 4655 6146 4664
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6012 3670 6040 4082
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6092 2916 6144 2922
rect 6092 2858 6144 2864
rect 6104 2582 6132 2858
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 5816 604 5868 610
rect 5816 546 5868 552
rect 6196 480 6224 6598
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5166 6868 5510
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6932 4978 6960 7142
rect 7024 6361 7052 9046
rect 7300 8974 7328 9318
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7954 7236 8230
rect 7300 8090 7328 8910
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7208 7002 7236 7890
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7010 6352 7066 6361
rect 7010 6287 7066 6296
rect 7024 5953 7052 6287
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7010 5944 7066 5953
rect 7010 5879 7066 5888
rect 7208 5681 7236 6054
rect 7194 5672 7250 5681
rect 7012 5636 7064 5642
rect 7194 5607 7250 5616
rect 7012 5578 7064 5584
rect 6656 4950 6960 4978
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6380 4185 6408 4490
rect 6366 4176 6422 4185
rect 6366 4111 6422 4120
rect 6276 4072 6328 4078
rect 6274 4040 6276 4049
rect 6328 4040 6330 4049
rect 6274 3975 6330 3984
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6656 1034 6684 4950
rect 7024 4826 7052 5578
rect 7392 5273 7420 9454
rect 7470 7848 7526 7857
rect 7470 7783 7526 7792
rect 7484 7546 7512 7783
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7484 7342 7512 7482
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7576 6458 7604 14470
rect 7760 14396 7788 14606
rect 7668 14368 7788 14396
rect 7668 11506 7696 14368
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 12238 7788 14214
rect 7852 13530 7880 14878
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 13297 7880 13330
rect 7838 13288 7894 13297
rect 7838 13223 7840 13232
rect 7892 13223 7894 13232
rect 7840 13194 7892 13200
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7852 11762 7880 12786
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7668 11478 7788 11506
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7576 6254 7604 6394
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7562 5944 7618 5953
rect 7562 5879 7618 5888
rect 7378 5264 7434 5273
rect 7208 5208 7378 5216
rect 7208 5199 7434 5208
rect 7208 5188 7420 5199
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6748 3670 6776 3946
rect 7208 3738 7236 5188
rect 7392 5139 7420 5188
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7288 4480 7340 4486
rect 7286 4448 7288 4457
rect 7340 4448 7342 4457
rect 7286 4383 7342 4392
rect 7392 4078 7420 4966
rect 7470 4584 7526 4593
rect 7470 4519 7472 4528
rect 7524 4519 7526 4528
rect 7472 4490 7524 4496
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6840 3194 6868 3674
rect 7576 3466 7604 5879
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7024 3194 7052 3402
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6840 2650 6868 2994
rect 7668 2825 7696 11222
rect 7760 6225 7788 11478
rect 7944 11286 7972 21286
rect 8036 18834 8064 25978
rect 8128 21350 8156 26846
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 8220 26042 8248 26386
rect 8312 26382 8340 26998
rect 8404 26790 8432 29135
rect 8666 29064 8722 29073
rect 8666 28999 8722 29008
rect 8576 28484 8628 28490
rect 8576 28426 8628 28432
rect 8484 28076 8536 28082
rect 8484 28018 8536 28024
rect 8496 27674 8524 28018
rect 8588 28014 8616 28426
rect 8576 28008 8628 28014
rect 8576 27950 8628 27956
rect 8484 27668 8536 27674
rect 8484 27610 8536 27616
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8208 25832 8260 25838
rect 8208 25774 8260 25780
rect 8220 25401 8248 25774
rect 8206 25392 8262 25401
rect 8206 25327 8262 25336
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8220 24410 8248 25230
rect 8312 24818 8340 26318
rect 8404 25294 8432 26726
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8404 24818 8432 25094
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8208 24404 8260 24410
rect 8208 24346 8260 24352
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8220 22166 8248 24006
rect 8298 23216 8354 23225
rect 8298 23151 8354 23160
rect 8312 22778 8340 23151
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8312 22234 8340 22578
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8208 21480 8260 21486
rect 8206 21448 8208 21457
rect 8260 21448 8262 21457
rect 8206 21383 8262 21392
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8220 21146 8248 21383
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 19854 8248 20198
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8312 19700 8340 21966
rect 8220 19672 8340 19700
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 8114 18728 8170 18737
rect 8114 18663 8170 18672
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8036 15706 8064 16730
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8036 14074 8064 14418
rect 8128 14278 8156 18663
rect 8220 18193 8248 19672
rect 8496 19258 8524 27406
rect 8574 27160 8630 27169
rect 8574 27095 8576 27104
rect 8628 27095 8630 27104
rect 8576 27066 8628 27072
rect 8574 26616 8630 26625
rect 8574 26551 8630 26560
rect 8588 19281 8616 26551
rect 8680 26466 8708 28999
rect 8772 27470 8800 31878
rect 8864 29073 8892 32399
rect 9404 32370 9456 32376
rect 9496 32428 9548 32434
rect 9496 32370 9548 32376
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 8944 32224 8996 32230
rect 9324 32212 9352 32302
rect 9416 32280 9444 32370
rect 9416 32252 9536 32280
rect 9324 32184 9444 32212
rect 8944 32166 8996 32172
rect 8956 31958 8984 32166
rect 9310 32056 9366 32065
rect 9310 31991 9366 32000
rect 8944 31952 8996 31958
rect 8944 31894 8996 31900
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 9220 29232 9272 29238
rect 9220 29174 9272 29180
rect 8850 29064 8906 29073
rect 8850 28999 8906 29008
rect 8852 28620 8904 28626
rect 8852 28562 8904 28568
rect 8864 28422 8892 28562
rect 9232 28529 9260 29174
rect 9324 29102 9352 31991
rect 9312 29096 9364 29102
rect 9312 29038 9364 29044
rect 9218 28520 9274 28529
rect 9218 28455 9274 28464
rect 8852 28416 8904 28422
rect 8852 28358 8904 28364
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8772 26586 8800 27270
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8680 26438 8800 26466
rect 8668 25492 8720 25498
rect 8668 25434 8720 25440
rect 8680 23866 8708 25434
rect 8668 23860 8720 23866
rect 8668 23802 8720 23808
rect 8772 23746 8800 26438
rect 8680 23718 8800 23746
rect 8680 21894 8708 23718
rect 8760 23656 8812 23662
rect 8760 23598 8812 23604
rect 8772 22982 8800 23598
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8758 21448 8814 21457
rect 8758 21383 8814 21392
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8312 19230 8524 19258
rect 8574 19272 8630 19281
rect 8206 18184 8262 18193
rect 8206 18119 8262 18128
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15162 8248 15438
rect 8312 15162 8340 19230
rect 8574 19207 8630 19216
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 16561 8432 19110
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8496 18086 8524 18770
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18426 8616 18702
rect 8680 18698 8708 19654
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16794 8524 16934
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8390 16552 8446 16561
rect 8390 16487 8446 16496
rect 8588 16046 8616 18362
rect 8680 18222 8708 18634
rect 8772 18442 8800 21383
rect 8864 19174 8892 28358
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 9416 27985 9444 32184
rect 9508 31754 9536 32252
rect 9496 31748 9548 31754
rect 9496 31690 9548 31696
rect 9508 31142 9536 31690
rect 9496 31136 9548 31142
rect 9496 31078 9548 31084
rect 9508 30394 9536 31078
rect 9496 30388 9548 30394
rect 9496 30330 9548 30336
rect 9496 29708 9548 29714
rect 9496 29650 9548 29656
rect 9402 27976 9458 27985
rect 9402 27911 9458 27920
rect 9508 27470 9536 29650
rect 9600 29238 9628 32830
rect 9692 32570 9720 32966
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9692 32473 9720 32506
rect 9678 32464 9734 32473
rect 9678 32399 9734 32408
rect 9784 31278 9812 39520
rect 10048 35624 10100 35630
rect 10048 35566 10100 35572
rect 9864 35216 9916 35222
rect 9864 35158 9916 35164
rect 9876 34746 9904 35158
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9876 34202 9904 34682
rect 9956 34536 10008 34542
rect 9954 34504 9956 34513
rect 10008 34504 10010 34513
rect 9954 34439 10010 34448
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 9862 33552 9918 33561
rect 9862 33487 9918 33496
rect 9876 33386 9904 33487
rect 9864 33380 9916 33386
rect 9864 33322 9916 33328
rect 10060 32230 10088 35566
rect 10152 33402 10180 39520
rect 10322 35184 10378 35193
rect 10322 35119 10378 35128
rect 10336 34746 10364 35119
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10508 34400 10560 34406
rect 10612 34377 10640 39520
rect 10704 39494 11008 39520
rect 11256 39494 11376 39520
rect 10508 34342 10560 34348
rect 10598 34368 10654 34377
rect 10520 33522 10548 34342
rect 10598 34303 10654 34312
rect 10508 33516 10560 33522
rect 10508 33458 10560 33464
rect 10152 33374 10272 33402
rect 10140 33312 10192 33318
rect 10140 33254 10192 33260
rect 10152 32910 10180 33254
rect 10140 32904 10192 32910
rect 10140 32846 10192 32852
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 10060 32065 10088 32166
rect 10046 32056 10102 32065
rect 10046 31991 10102 32000
rect 10152 31958 10180 32846
rect 10140 31952 10192 31958
rect 10140 31894 10192 31900
rect 10048 31884 10100 31890
rect 10048 31826 10100 31832
rect 10060 31482 10088 31826
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 9772 31272 9824 31278
rect 9772 31214 9824 31220
rect 10048 31272 10100 31278
rect 10048 31214 10100 31220
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9678 30696 9734 30705
rect 9678 30631 9680 30640
rect 9732 30631 9734 30640
rect 9680 30602 9732 30608
rect 9680 30116 9732 30122
rect 9680 30058 9732 30064
rect 9588 29232 9640 29238
rect 9588 29174 9640 29180
rect 9588 29096 9640 29102
rect 9588 29038 9640 29044
rect 9496 27464 9548 27470
rect 9496 27406 9548 27412
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9324 25786 9352 26522
rect 9416 26042 9444 27270
rect 9496 26988 9548 26994
rect 9496 26930 9548 26936
rect 9508 26586 9536 26930
rect 9600 26790 9628 29038
rect 9692 28966 9720 30058
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9678 27840 9734 27849
rect 9678 27775 9734 27784
rect 9692 27674 9720 27775
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9588 26784 9640 26790
rect 9588 26726 9640 26732
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9692 26450 9720 27406
rect 9680 26444 9732 26450
rect 9680 26386 9732 26392
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9496 26240 9548 26246
rect 9496 26182 9548 26188
rect 9404 26036 9456 26042
rect 9404 25978 9456 25984
rect 9508 25922 9536 26182
rect 9232 25758 9352 25786
rect 9416 25894 9536 25922
rect 9416 25770 9444 25894
rect 9496 25832 9548 25838
rect 9600 25786 9628 26318
rect 9548 25780 9628 25786
rect 9496 25774 9628 25780
rect 9404 25764 9456 25770
rect 9232 25498 9260 25758
rect 9404 25706 9456 25712
rect 9508 25758 9628 25774
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9220 25492 9272 25498
rect 9220 25434 9272 25440
rect 9324 25158 9352 25638
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9324 24954 9352 25094
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 8944 24744 8996 24750
rect 8942 24712 8944 24721
rect 8996 24712 8998 24721
rect 8942 24647 8998 24656
rect 9310 24712 9366 24721
rect 9310 24647 9366 24656
rect 9324 24614 9352 24647
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9324 24070 9352 24550
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9324 23322 9352 23598
rect 9312 23316 9364 23322
rect 9312 23258 9364 23264
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 9324 20942 9352 22918
rect 9416 22778 9444 25706
rect 9508 23526 9536 25758
rect 9692 25702 9720 26386
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9600 24818 9628 25434
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9508 21894 9536 22374
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 9324 20466 9352 20878
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9324 20058 9352 20402
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 8772 18414 8892 18442
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8588 15706 8616 15982
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8482 15600 8538 15609
rect 8392 15564 8444 15570
rect 8482 15535 8484 15544
rect 8392 15506 8444 15512
rect 8536 15535 8538 15544
rect 8484 15506 8536 15512
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8312 14618 8340 14962
rect 8404 14793 8432 15506
rect 8588 15502 8616 15642
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8390 14784 8446 14793
rect 8390 14719 8446 14728
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8036 13841 8064 14010
rect 8022 13832 8078 13841
rect 8022 13767 8078 13776
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8128 12714 8156 13466
rect 8312 12782 8340 13670
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7852 10266 7880 11154
rect 8036 11150 8064 11698
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7944 10810 7972 11086
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 8036 10130 8064 11086
rect 8128 10470 8156 12310
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11558 8248 12174
rect 8404 11762 8432 12650
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11098 8248 11494
rect 8404 11286 8432 11698
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8220 11070 8340 11098
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7852 9586 7880 9930
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 8294 7880 9522
rect 8206 9344 8262 9353
rect 8206 9279 8262 9288
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7206 7880 7686
rect 8220 7342 8248 9279
rect 8312 8022 8340 11070
rect 8496 10169 8524 15370
rect 8588 15026 8616 15438
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8588 13870 8616 14350
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8588 10674 8616 13806
rect 8680 12753 8708 18022
rect 8772 17542 8800 18226
rect 8760 17536 8812 17542
rect 8864 17524 8892 18414
rect 9416 18222 9444 19110
rect 9508 18902 9536 19246
rect 9496 18896 9548 18902
rect 9496 18838 9548 18844
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9508 18222 9536 18566
rect 9404 18216 9456 18222
rect 9310 18184 9366 18193
rect 9404 18158 9456 18164
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9310 18119 9366 18128
rect 9324 17746 9352 18119
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 8864 17496 9352 17524
rect 8760 17478 8812 17484
rect 8772 17202 8800 17478
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8772 16250 8800 17138
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8864 16658 8892 16934
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8864 15162 8892 16594
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 9324 14958 9352 17496
rect 9416 16794 9444 18158
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9508 17338 9536 17750
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8666 12744 8722 12753
rect 8666 12679 8722 12688
rect 8772 12646 8800 13262
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8680 12442 8708 12582
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8680 11558 8708 12378
rect 8772 11694 8800 12582
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8482 10160 8538 10169
rect 8392 10124 8444 10130
rect 8482 10095 8538 10104
rect 8392 10066 8444 10072
rect 8404 9722 8432 10066
rect 8588 10062 8616 10610
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8496 9450 8524 9998
rect 8588 9518 8616 9998
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8588 8974 8616 9454
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8090 8616 8910
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8300 8016 8352 8022
rect 8352 7964 8432 7970
rect 8300 7958 8432 7964
rect 8312 7942 8432 7958
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7746 6216 7802 6225
rect 7746 6151 7802 6160
rect 7760 4298 7788 6151
rect 7852 5914 7880 7142
rect 8220 7002 8248 7278
rect 8312 7041 8340 7754
rect 8404 7177 8432 7942
rect 8680 7449 8708 11494
rect 8772 11354 8800 11630
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8772 8634 8800 8978
rect 8864 8634 8892 14894
rect 9324 14618 9352 14894
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 9324 9042 9352 13126
rect 9508 12714 9536 17002
rect 9600 15434 9628 24346
rect 9692 22522 9720 25638
rect 9784 23186 9812 31078
rect 9864 30796 9916 30802
rect 9864 30738 9916 30744
rect 9876 30122 9904 30738
rect 9864 30116 9916 30122
rect 9864 30058 9916 30064
rect 9864 29776 9916 29782
rect 9864 29718 9916 29724
rect 9876 29170 9904 29718
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9876 29034 9904 29106
rect 9864 29028 9916 29034
rect 9864 28970 9916 28976
rect 9876 28762 9904 28970
rect 9864 28756 9916 28762
rect 9864 28698 9916 28704
rect 9876 28218 9904 28698
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9876 26625 9904 26726
rect 9862 26616 9918 26625
rect 9862 26551 9918 26560
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9968 25702 9996 26318
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9876 22642 9904 23258
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9968 22545 9996 25638
rect 10060 25480 10088 31214
rect 10152 31142 10180 31758
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10140 30932 10192 30938
rect 10140 30874 10192 30880
rect 10152 30054 10180 30874
rect 10244 30818 10272 33374
rect 10508 32972 10560 32978
rect 10508 32914 10560 32920
rect 10324 32768 10376 32774
rect 10324 32710 10376 32716
rect 10336 31346 10364 32710
rect 10520 32570 10548 32914
rect 10508 32564 10560 32570
rect 10508 32506 10560 32512
rect 10506 31784 10562 31793
rect 10704 31770 10732 39494
rect 11152 34944 11204 34950
rect 11152 34886 11204 34892
rect 10874 34640 10930 34649
rect 11164 34610 11192 34886
rect 10874 34575 10930 34584
rect 11152 34604 11204 34610
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10796 33114 10824 33458
rect 10784 33108 10836 33114
rect 10784 33050 10836 33056
rect 10796 32502 10824 33050
rect 10784 32496 10836 32502
rect 10784 32438 10836 32444
rect 10796 32026 10824 32438
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10888 31890 10916 34575
rect 11152 34546 11204 34552
rect 11164 34066 11192 34546
rect 11152 34060 11204 34066
rect 11152 34002 11204 34008
rect 11164 33658 11192 34002
rect 11152 33652 11204 33658
rect 11152 33594 11204 33600
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 11164 32026 11192 32846
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 10876 31884 10928 31890
rect 10876 31826 10928 31832
rect 10506 31719 10562 31728
rect 10612 31742 10732 31770
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10414 31240 10470 31249
rect 10414 31175 10470 31184
rect 10428 31142 10456 31175
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10520 30938 10548 31719
rect 10508 30932 10560 30938
rect 10508 30874 10560 30880
rect 10244 30790 10364 30818
rect 10232 30728 10284 30734
rect 10232 30670 10284 30676
rect 10244 30394 10272 30670
rect 10232 30388 10284 30394
rect 10232 30330 10284 30336
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10152 26382 10180 29990
rect 10244 29850 10272 30330
rect 10232 29844 10284 29850
rect 10232 29786 10284 29792
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10244 26761 10272 27406
rect 10230 26752 10286 26761
rect 10230 26687 10286 26696
rect 10244 26586 10272 26687
rect 10232 26580 10284 26586
rect 10232 26522 10284 26528
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10140 25492 10192 25498
rect 10060 25452 10140 25480
rect 10140 25434 10192 25440
rect 10046 25256 10102 25265
rect 10046 25191 10048 25200
rect 10100 25191 10102 25200
rect 10048 25162 10100 25168
rect 10060 24954 10088 25162
rect 10048 24948 10100 24954
rect 10048 24890 10100 24896
rect 10152 24070 10180 25434
rect 10336 24857 10364 30790
rect 10612 29209 10640 31742
rect 11164 31482 11192 31962
rect 11152 31476 11204 31482
rect 11152 31418 11204 31424
rect 10966 31376 11022 31385
rect 10876 31340 10928 31346
rect 10966 31311 10968 31320
rect 10876 31282 10928 31288
rect 11020 31311 11022 31320
rect 10968 31282 11020 31288
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10796 30666 10824 31078
rect 10888 30938 10916 31282
rect 10876 30932 10928 30938
rect 10876 30874 10928 30880
rect 10980 30870 11008 31282
rect 10968 30864 11020 30870
rect 10968 30806 11020 30812
rect 10784 30660 10836 30666
rect 10784 30602 10836 30608
rect 10796 30394 10824 30602
rect 10980 30410 11008 30806
rect 11164 30734 11192 31418
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 10784 30388 10836 30394
rect 10980 30382 11100 30410
rect 11164 30394 11192 30670
rect 10784 30330 10836 30336
rect 10784 29708 10836 29714
rect 10784 29650 10836 29656
rect 10598 29200 10654 29209
rect 10598 29135 10654 29144
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 10428 27130 10456 29038
rect 10796 28966 10824 29650
rect 10784 28960 10836 28966
rect 10784 28902 10836 28908
rect 11072 28694 11100 30382
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 10600 28620 10652 28626
rect 10600 28562 10652 28568
rect 10612 27878 10640 28562
rect 11072 28218 11100 28630
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10600 27872 10652 27878
rect 10600 27814 10652 27820
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 10980 27554 11008 27814
rect 10980 27526 11192 27554
rect 11164 27334 11192 27526
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10428 26926 10456 27066
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 10416 26920 10468 26926
rect 10416 26862 10468 26868
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10796 25906 10824 26726
rect 11072 26382 11100 26930
rect 11060 26376 11112 26382
rect 11060 26318 11112 26324
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10876 25968 10928 25974
rect 10876 25910 10928 25916
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 10520 25430 10548 25774
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10508 25424 10560 25430
rect 10508 25366 10560 25372
rect 10508 25220 10560 25226
rect 10508 25162 10560 25168
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10322 24848 10378 24857
rect 10322 24783 10378 24792
rect 10428 24682 10456 25094
rect 10416 24676 10468 24682
rect 10416 24618 10468 24624
rect 10324 24608 10376 24614
rect 10322 24576 10324 24585
rect 10376 24576 10378 24585
rect 10322 24511 10378 24520
rect 10428 24410 10456 24618
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10520 24290 10548 25162
rect 10612 24410 10640 25638
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10428 24262 10548 24290
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10060 23322 10088 24006
rect 10048 23316 10100 23322
rect 10048 23258 10100 23264
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 9954 22536 10010 22545
rect 9692 22494 9904 22522
rect 9678 22264 9734 22273
rect 9678 22199 9680 22208
rect 9732 22199 9734 22208
rect 9772 22228 9824 22234
rect 9680 22170 9732 22176
rect 9772 22170 9824 22176
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9692 19174 9720 19654
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 17882 9720 19110
rect 9784 18465 9812 22170
rect 9876 20369 9904 22494
rect 9954 22471 10010 22480
rect 10060 22234 10088 23122
rect 10048 22228 10100 22234
rect 10048 22170 10100 22176
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9968 21690 9996 22102
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9968 20505 9996 21626
rect 10060 21350 10088 22034
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 21146 10088 21286
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 9954 20496 10010 20505
rect 9954 20431 10010 20440
rect 9862 20360 9918 20369
rect 9862 20295 9918 20304
rect 9954 20224 10010 20233
rect 9954 20159 10010 20168
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9876 19446 9904 19654
rect 9864 19440 9916 19446
rect 9864 19382 9916 19388
rect 9876 19310 9904 19382
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9862 18864 9918 18873
rect 9862 18799 9864 18808
rect 9916 18799 9918 18808
rect 9864 18770 9916 18776
rect 9862 18728 9918 18737
rect 9862 18663 9918 18672
rect 9770 18456 9826 18465
rect 9770 18391 9826 18400
rect 9876 17882 9904 18663
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9784 17066 9812 17682
rect 9876 17338 9904 17818
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9968 17218 9996 20159
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9876 17190 9996 17218
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9678 16144 9734 16153
rect 9678 16079 9734 16088
rect 9692 16046 9720 16079
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9600 14249 9628 14826
rect 9678 14784 9734 14793
rect 9678 14719 9734 14728
rect 9692 14618 9720 14719
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9586 14240 9642 14249
rect 9586 14175 9642 14184
rect 9678 13696 9734 13705
rect 9678 13631 9734 13640
rect 9692 12986 9720 13631
rect 9784 13190 9812 15030
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9494 11792 9550 11801
rect 9494 11727 9550 11736
rect 9402 10976 9458 10985
rect 9402 10911 9458 10920
rect 9416 10606 9444 10911
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 9897 9444 10406
rect 9402 9888 9458 9897
rect 9402 9823 9458 9832
rect 9402 9752 9458 9761
rect 9402 9687 9458 9696
rect 9416 9450 9444 9687
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8772 8514 8800 8570
rect 8772 8486 8892 8514
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8666 7440 8722 7449
rect 8666 7375 8722 7384
rect 8484 7200 8536 7206
rect 8390 7168 8446 7177
rect 8484 7142 8536 7148
rect 8390 7103 8446 7112
rect 8298 7032 8354 7041
rect 8208 6996 8260 7002
rect 8298 6967 8354 6976
rect 8208 6938 8260 6944
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8404 6458 8432 6802
rect 8496 6798 8524 7142
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8496 5914 8524 6734
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8300 5704 8352 5710
rect 7930 5672 7986 5681
rect 8300 5646 8352 5652
rect 7930 5607 7986 5616
rect 7760 4270 7880 4298
rect 7746 4176 7802 4185
rect 7746 4111 7802 4120
rect 7654 2816 7710 2825
rect 7654 2751 7710 2760
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1465 7144 2246
rect 7102 1456 7158 1465
rect 7102 1391 7158 1400
rect 6564 1006 6684 1034
rect 6564 480 6592 1006
rect 6920 604 6972 610
rect 6920 546 6972 552
rect 7380 604 7432 610
rect 7380 546 7432 552
rect 6932 480 6960 546
rect 7392 480 7420 546
rect 7760 480 7788 4111
rect 7852 3670 7880 4270
rect 7944 3738 7972 5607
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 4214 8064 5034
rect 8220 4826 8248 5510
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8312 4486 8340 5646
rect 8404 4554 8432 5714
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8300 4480 8352 4486
rect 8128 4428 8300 4434
rect 8128 4422 8352 4428
rect 8128 4406 8340 4422
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7852 2922 7880 3606
rect 7944 2990 7972 3674
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7930 2816 7986 2825
rect 7930 2751 7986 2760
rect 7944 2650 7972 2751
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7944 2514 7972 2586
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8036 610 8064 3975
rect 8128 2650 8156 4406
rect 8404 4298 8432 4490
rect 8220 4270 8432 4298
rect 8220 3194 8248 4270
rect 8496 4078 8524 4558
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8588 3738 8616 6598
rect 8680 6118 8708 6734
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5710 8708 6054
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8680 5098 8708 5646
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8680 3618 8708 4626
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8588 3590 8708 3618
rect 8772 3602 8800 8366
rect 8864 6440 8892 8486
rect 9508 8430 9536 11727
rect 9496 8424 9548 8430
rect 9692 8401 9720 12271
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11218 9812 11494
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9784 10266 9812 11154
rect 9876 10470 9904 17190
rect 10060 17116 10088 19110
rect 10152 19009 10180 24006
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 22030 10272 23462
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10244 21690 10272 21966
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10244 19922 10272 20878
rect 10336 20058 10364 22510
rect 10324 20052 10376 20058
rect 10324 19994 10376 20000
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10336 19174 10364 19994
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10138 19000 10194 19009
rect 10138 18935 10194 18944
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10152 18086 10180 18838
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9968 17088 10088 17116
rect 9968 14090 9996 17088
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 15706 10088 16526
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10152 15008 10180 18022
rect 10244 17814 10272 18702
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18426 10364 18566
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10336 17241 10364 18022
rect 10322 17232 10378 17241
rect 10322 17167 10378 17176
rect 10428 17134 10456 24262
rect 10612 23254 10640 24346
rect 10704 24274 10732 24550
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10888 24206 10916 25910
rect 10980 25838 11008 26182
rect 11072 26042 11100 26318
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 11072 25684 11100 25978
rect 10980 25656 11100 25684
rect 10980 25294 11008 25656
rect 11164 25430 11192 27270
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10796 23866 10824 24142
rect 11072 23866 11100 24210
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 10796 23662 10824 23802
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 11164 23322 11192 24142
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 10600 23112 10652 23118
rect 10506 23080 10562 23089
rect 10600 23054 10652 23060
rect 10506 23015 10508 23024
rect 10560 23015 10562 23024
rect 10508 22986 10560 22992
rect 10612 22778 10640 23054
rect 10888 22778 10916 23258
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 10782 22536 10838 22545
rect 10782 22471 10838 22480
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10612 19156 10640 21830
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10704 19378 10732 20198
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10692 19168 10744 19174
rect 10612 19128 10692 19156
rect 10692 19110 10744 19116
rect 10704 18630 10732 19110
rect 10692 18624 10744 18630
rect 10690 18592 10692 18601
rect 10744 18592 10746 18601
rect 10690 18527 10746 18536
rect 10600 18216 10652 18222
rect 10598 18184 10600 18193
rect 10652 18184 10654 18193
rect 10598 18119 10654 18128
rect 10690 17640 10746 17649
rect 10690 17575 10746 17584
rect 10704 17338 10732 17575
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10796 17218 10824 22471
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10980 20618 11008 20946
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 10980 20602 11100 20618
rect 10980 20596 11112 20602
rect 10980 20590 11060 20596
rect 11060 20538 11112 20544
rect 11072 20074 11100 20538
rect 11164 20330 11192 20742
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 10888 20058 11100 20074
rect 10888 20052 11112 20058
rect 10888 20046 11060 20052
rect 10888 18290 10916 20046
rect 11060 19994 11112 20000
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10980 19292 11008 19926
rect 11164 19378 11192 20266
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11060 19304 11112 19310
rect 10980 19264 11060 19292
rect 11060 19246 11112 19252
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18834 11100 19110
rect 11164 18970 11192 19314
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10888 17882 10916 18226
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10980 17626 11008 18362
rect 11072 18086 11100 18770
rect 11164 18766 11192 18906
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11256 18578 11284 39494
rect 11808 37754 11836 39520
rect 11532 37726 11836 37754
rect 11428 36168 11480 36174
rect 11428 36110 11480 36116
rect 11440 35562 11468 36110
rect 11428 35556 11480 35562
rect 11428 35498 11480 35504
rect 11440 35154 11468 35498
rect 11428 35148 11480 35154
rect 11428 35090 11480 35096
rect 11440 33862 11468 35090
rect 11428 33856 11480 33862
rect 11428 33798 11480 33804
rect 11440 33318 11468 33798
rect 11428 33312 11480 33318
rect 11428 33254 11480 33260
rect 11336 32224 11388 32230
rect 11334 32192 11336 32201
rect 11388 32192 11390 32201
rect 11334 32127 11390 32136
rect 11440 31890 11468 33254
rect 11428 31884 11480 31890
rect 11428 31826 11480 31832
rect 11440 28966 11468 31826
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 11440 28642 11468 28902
rect 11348 28626 11468 28642
rect 11336 28620 11468 28626
rect 11388 28614 11468 28620
rect 11336 28562 11388 28568
rect 11440 28218 11468 28614
rect 11428 28212 11480 28218
rect 11428 28154 11480 28160
rect 11440 27674 11468 28154
rect 11428 27668 11480 27674
rect 11348 27628 11428 27656
rect 11348 26586 11376 27628
rect 11428 27610 11480 27616
rect 11426 27568 11482 27577
rect 11426 27503 11428 27512
rect 11480 27503 11482 27512
rect 11428 27474 11480 27480
rect 11440 27130 11468 27474
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 11348 25226 11376 25842
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 11348 24818 11376 25162
rect 11336 24812 11388 24818
rect 11388 24772 11468 24800
rect 11336 24754 11388 24760
rect 11336 24676 11388 24682
rect 11336 24618 11388 24624
rect 11348 23746 11376 24618
rect 11440 24410 11468 24772
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11440 23866 11468 24346
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11348 23718 11468 23746
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11348 22778 11376 23190
rect 11440 22778 11468 23718
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11532 22658 11560 37726
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11612 36236 11664 36242
rect 11612 36178 11664 36184
rect 11624 35834 11652 36178
rect 11612 35828 11664 35834
rect 11612 35770 11664 35776
rect 11980 35828 12032 35834
rect 11980 35770 12032 35776
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11992 34202 12020 35770
rect 11980 34196 12032 34202
rect 11980 34138 12032 34144
rect 11992 33522 12020 34138
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11992 32858 12020 33458
rect 12176 32881 12204 39520
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12256 33312 12308 33318
rect 12256 33254 12308 33260
rect 12268 33046 12296 33254
rect 12256 33040 12308 33046
rect 12452 32994 12480 35974
rect 12256 32982 12308 32988
rect 12360 32966 12480 32994
rect 12256 32904 12308 32910
rect 12162 32872 12218 32881
rect 11992 32842 12112 32858
rect 11992 32836 12124 32842
rect 11992 32830 12072 32836
rect 12360 32858 12388 32966
rect 12308 32852 12388 32858
rect 12256 32846 12388 32852
rect 12268 32830 12388 32846
rect 12162 32807 12218 32816
rect 12072 32778 12124 32784
rect 11980 32768 12032 32774
rect 11980 32710 12032 32716
rect 12084 32722 12112 32778
rect 12346 32736 12402 32745
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11796 30864 11848 30870
rect 11888 30864 11940 30870
rect 11848 30824 11888 30852
rect 11796 30806 11848 30812
rect 11888 30806 11940 30812
rect 11808 30394 11836 30806
rect 11992 30802 12020 32710
rect 12084 32694 12204 32722
rect 12072 32292 12124 32298
rect 12072 32234 12124 32240
rect 11980 30796 12032 30802
rect 11980 30738 12032 30744
rect 11992 30394 12020 30738
rect 11796 30388 11848 30394
rect 11796 30330 11848 30336
rect 11980 30388 12032 30394
rect 11980 30330 12032 30336
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11992 27606 12020 28358
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 11992 27062 12020 27542
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 12084 26874 12112 32234
rect 12176 31482 12204 32694
rect 12346 32671 12402 32680
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 12268 31482 12296 31826
rect 12164 31476 12216 31482
rect 12164 31418 12216 31424
rect 12256 31476 12308 31482
rect 12256 31418 12308 31424
rect 12360 31090 12388 32671
rect 12544 32298 12572 39520
rect 12532 32292 12584 32298
rect 12532 32234 12584 32240
rect 12440 32224 12492 32230
rect 12440 32166 12492 32172
rect 12268 31062 12388 31090
rect 12162 30016 12218 30025
rect 12162 29951 12218 29960
rect 12176 28121 12204 29951
rect 12162 28112 12218 28121
rect 12162 28047 12218 28056
rect 12162 27976 12218 27985
rect 12162 27911 12218 27920
rect 11992 26846 12112 26874
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11348 22630 11560 22658
rect 11348 18902 11376 22630
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 11256 18550 11376 18578
rect 11242 18456 11298 18465
rect 11242 18391 11298 18400
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10704 17190 10824 17218
rect 10888 17598 11008 17626
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10428 16697 10456 16730
rect 10414 16688 10470 16697
rect 10324 16652 10376 16658
rect 10414 16623 10470 16632
rect 10324 16594 10376 16600
rect 10336 15162 10364 16594
rect 10598 16008 10654 16017
rect 10598 15943 10600 15952
rect 10652 15943 10654 15952
rect 10600 15914 10652 15920
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10152 14980 10364 15008
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10060 14385 10088 14758
rect 10244 14521 10272 14758
rect 10230 14512 10286 14521
rect 10230 14447 10286 14456
rect 10046 14376 10102 14385
rect 10046 14311 10102 14320
rect 10232 14340 10284 14346
rect 10060 14278 10088 14311
rect 10232 14282 10284 14288
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9968 14062 10088 14090
rect 10060 13394 10088 14062
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9968 12442 9996 13262
rect 10060 12646 10088 13330
rect 10244 13297 10272 14282
rect 10230 13288 10286 13297
rect 10230 13223 10286 13232
rect 10048 12640 10100 12646
rect 10046 12608 10048 12617
rect 10100 12608 10102 12617
rect 10046 12543 10102 12552
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9968 12170 9996 12378
rect 10138 12336 10194 12345
rect 10138 12271 10194 12280
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10060 11898 10088 12174
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9956 11212 10008 11218
rect 10060 11200 10088 11834
rect 10008 11172 10088 11200
rect 9956 11154 10008 11160
rect 9968 10810 9996 11154
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 10060 9518 10088 9551
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9864 9376 9916 9382
rect 9862 9344 9864 9353
rect 9916 9344 9918 9353
rect 9862 9279 9918 9288
rect 10152 8922 10180 12271
rect 10336 11801 10364 14980
rect 10428 14414 10456 15506
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10612 13410 10640 15914
rect 10704 15706 10732 17190
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10704 15094 10732 15642
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10796 13433 10824 17070
rect 10428 13382 10640 13410
rect 10782 13424 10838 13433
rect 10428 12481 10456 13382
rect 10782 13359 10838 13368
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10414 12472 10470 12481
rect 10414 12407 10470 12416
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10322 11792 10378 11801
rect 10322 11727 10378 11736
rect 10428 11286 10456 12242
rect 10520 12238 10548 13126
rect 10612 12986 10640 13262
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10796 12594 10824 13359
rect 10888 13274 10916 17598
rect 11072 17542 11100 18022
rect 11164 17610 11192 18090
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11060 17536 11112 17542
rect 10980 17496 11060 17524
rect 10980 17202 11008 17496
rect 11060 17478 11112 17484
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10980 16590 11008 17138
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16658 11100 17070
rect 11164 16998 11192 17274
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10980 16182 11008 16526
rect 11072 16250 11100 16594
rect 11164 16454 11192 16934
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 15026 11100 15438
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11072 14618 11100 14962
rect 11164 14822 11192 15506
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10888 13246 11100 13274
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12850 11008 13126
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10612 12566 10824 12594
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11898 10548 12174
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10506 11792 10562 11801
rect 10506 11727 10562 11736
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10428 10810 10456 11222
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10520 10538 10548 11727
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10152 8894 10364 8922
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8498 10272 8774
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10140 8424 10192 8430
rect 9496 8366 9548 8372
rect 9678 8392 9734 8401
rect 10140 8366 10192 8372
rect 9678 8327 9734 8336
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9220 7472 9272 7478
rect 9218 7440 9220 7449
rect 9272 7440 9274 7449
rect 9218 7375 9274 7384
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 7002 9168 7278
rect 9220 7200 9272 7206
rect 9324 7188 9352 7686
rect 9272 7160 9352 7188
rect 9220 7142 9272 7148
rect 9416 7154 9444 8230
rect 9508 7818 9536 8230
rect 9692 8106 9720 8327
rect 9692 8078 9996 8106
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9232 7002 9260 7142
rect 9416 7126 9536 7154
rect 9402 7032 9458 7041
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9324 6990 9402 7018
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8864 6412 8984 6440
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8864 3670 8892 5782
rect 8956 5710 8984 6412
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 4690 9352 6990
rect 9402 6967 9458 6976
rect 9508 6848 9536 7126
rect 9416 6820 9536 6848
rect 9416 6322 9444 6820
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5817 9444 6054
rect 9508 5914 9536 6666
rect 9600 6322 9628 7482
rect 9692 7342 9720 7686
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9680 7200 9732 7206
rect 9678 7168 9680 7177
rect 9784 7188 9812 7822
rect 9876 7478 9904 7890
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9732 7168 9812 7188
rect 9734 7160 9812 7168
rect 9678 7103 9734 7112
rect 9968 6866 9996 8078
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9968 6458 9996 6802
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5846 9628 6258
rect 9588 5840 9640 5846
rect 9402 5808 9458 5817
rect 9588 5782 9640 5788
rect 9402 5743 9458 5752
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8760 3596 8812 3602
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8312 3097 8340 3334
rect 8404 3194 8432 3538
rect 8482 3360 8538 3369
rect 8482 3295 8538 3304
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8298 3088 8354 3097
rect 8298 3023 8354 3032
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8024 604 8076 610
rect 8024 546 8076 552
rect 8220 480 8248 2926
rect 8496 2825 8524 3295
rect 8482 2816 8538 2825
rect 8482 2751 8538 2760
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8496 2417 8524 2450
rect 8482 2408 8538 2417
rect 8482 2343 8538 2352
rect 8588 480 8616 3590
rect 8760 3538 8812 3544
rect 8760 3188 8812 3194
rect 8864 3176 8892 3606
rect 9140 3482 9168 3946
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3641 9352 3878
rect 9310 3632 9366 3641
rect 9416 3618 9444 5646
rect 9692 5556 9720 6394
rect 9508 5528 9720 5556
rect 9508 4078 9536 5528
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 3738 9536 3878
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9416 3590 9536 3618
rect 9310 3567 9366 3576
rect 9140 3454 9444 3482
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8812 3148 8892 3176
rect 8760 3130 8812 3136
rect 8772 2446 8800 3130
rect 8864 2990 8892 3148
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 9126 2952 9182 2961
rect 9126 2887 9182 2896
rect 8850 2816 8906 2825
rect 8850 2751 8906 2760
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8864 1442 8892 2751
rect 9140 2582 9168 2887
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8864 1414 8984 1442
rect 8956 480 8984 1414
rect 9416 480 9444 3454
rect 9508 2825 9536 3590
rect 9600 3176 9628 5034
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9692 4078 9720 4762
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9680 3188 9732 3194
rect 9600 3148 9680 3176
rect 9680 3130 9732 3136
rect 9678 2952 9734 2961
rect 9600 2922 9678 2938
rect 9588 2916 9678 2922
rect 9640 2910 9678 2916
rect 9678 2887 9734 2896
rect 9588 2858 9640 2864
rect 9494 2816 9550 2825
rect 9494 2751 9550 2760
rect 9692 2514 9720 2887
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9784 480 9812 4218
rect 9876 3738 9904 4655
rect 10060 4486 10088 5102
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10060 2961 10088 4422
rect 10046 2952 10102 2961
rect 10046 2887 10102 2896
rect 10152 480 10180 8366
rect 10244 7886 10272 8434
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10244 7274 10272 7822
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 6730 10272 7210
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10336 4690 10364 8894
rect 10428 5817 10456 10406
rect 10520 9926 10548 10474
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10520 7313 10548 9862
rect 10506 7304 10562 7313
rect 10506 7239 10562 7248
rect 10520 7002 10548 7239
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10520 6458 10548 6938
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10414 5808 10470 5817
rect 10414 5743 10470 5752
rect 10414 5128 10470 5137
rect 10414 5063 10470 5072
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10230 4584 10286 4593
rect 10230 4519 10286 4528
rect 10244 3126 10272 4519
rect 10336 3913 10364 4626
rect 10322 3904 10378 3913
rect 10322 3839 10378 3848
rect 10428 3754 10456 5063
rect 10612 4826 10640 12566
rect 10782 12472 10838 12481
rect 10782 12407 10838 12416
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11830 10732 12174
rect 10796 12073 10824 12407
rect 10888 12084 10916 12582
rect 10980 12442 11008 12786
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11072 12238 11100 13246
rect 11164 13161 11192 14758
rect 11150 13152 11206 13161
rect 11150 13087 11206 13096
rect 11164 12850 11192 13087
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11152 12096 11204 12102
rect 10782 12064 10838 12073
rect 10888 12056 11152 12084
rect 11152 12038 11204 12044
rect 10782 11999 10838 12008
rect 11164 11898 11192 12038
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 11060 11688 11112 11694
rect 10980 11636 11060 11642
rect 11256 11642 11284 18391
rect 11348 16046 11376 18550
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11348 15502 11376 15846
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11348 14890 11376 15438
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 11348 13326 11376 14826
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11348 12918 11376 13262
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11348 12238 11376 12854
rect 11440 12374 11468 22510
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11532 21350 11560 21966
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 20262 11560 21286
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11532 19922 11560 20198
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11532 18766 11560 19858
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11532 18426 11560 18702
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11900 16046 11928 16526
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11532 12374 11560 12922
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11992 12458 12020 26846
rect 12070 25392 12126 25401
rect 12070 25327 12126 25336
rect 12084 24886 12112 25327
rect 12072 24880 12124 24886
rect 12072 24822 12124 24828
rect 12176 24426 12204 27911
rect 12268 24682 12296 31062
rect 12452 30870 12480 32166
rect 12808 31680 12860 31686
rect 12808 31622 12860 31628
rect 12820 31385 12848 31622
rect 12806 31376 12862 31385
rect 12806 31311 12862 31320
rect 12440 30864 12492 30870
rect 12440 30806 12492 30812
rect 12900 28960 12952 28966
rect 12900 28902 12952 28908
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12256 24676 12308 24682
rect 12256 24618 12308 24624
rect 12176 24398 12296 24426
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 12084 23186 12112 23258
rect 12176 23186 12204 23598
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12084 22438 12112 23122
rect 12176 22778 12204 23122
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12268 22658 12296 24398
rect 12360 23662 12388 25094
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 23338 12480 23462
rect 12360 23322 12480 23338
rect 12348 23316 12480 23322
rect 12400 23310 12480 23316
rect 12348 23258 12400 23264
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12176 22630 12296 22658
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 12176 22012 12204 22630
rect 12360 22098 12388 22918
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 12084 21984 12204 22012
rect 12084 19242 12112 21984
rect 12360 21690 12388 22034
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12164 21480 12216 21486
rect 12544 21457 12572 26930
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12728 25362 12756 25638
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12728 24954 12756 25298
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12728 23662 12756 24550
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12636 23526 12664 23598
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12636 21690 12664 22374
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12164 21422 12216 21428
rect 12530 21448 12586 21457
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 12084 18970 12112 19178
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12070 18456 12126 18465
rect 12070 18391 12126 18400
rect 12084 18358 12112 18391
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12084 16794 12112 17750
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12084 16250 12112 16594
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12084 16114 12112 16186
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 12084 15706 12112 16050
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 12084 12646 12112 13398
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11983 12442 12020 12458
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11978 12336 12034 12345
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11334 12064 11390 12073
rect 11334 11999 11390 12008
rect 10980 11630 11112 11636
rect 10980 11614 11100 11630
rect 11164 11614 11284 11642
rect 10980 9382 11008 11614
rect 11058 9752 11114 9761
rect 11164 9738 11192 11614
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11286 11284 11494
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11242 9888 11298 9897
rect 11242 9823 11298 9832
rect 11114 9710 11192 9738
rect 11058 9687 11114 9696
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10704 7342 10732 8230
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10782 7304 10838 7313
rect 10782 7239 10838 7248
rect 10796 6458 10824 7239
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 11072 6322 11100 9687
rect 11256 6746 11284 9823
rect 11348 6848 11376 11999
rect 11440 7041 11468 12106
rect 11532 11762 11560 12310
rect 11978 12271 12034 12280
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 11354 11560 11698
rect 11624 11626 11652 12174
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11694 11836 12038
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11532 11150 11560 11290
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10810 11560 11086
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9382 11560 10066
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11992 8401 12020 12271
rect 12084 11830 12112 12582
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12084 10062 12112 10746
rect 12072 10056 12124 10062
rect 12176 10033 12204 21422
rect 12530 21383 12586 21392
rect 12636 21350 12664 21626
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12820 20913 12848 26862
rect 12912 22234 12940 28902
rect 13004 25809 13032 39520
rect 13084 32768 13136 32774
rect 13084 32710 13136 32716
rect 13096 32434 13124 32710
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 12990 25800 13046 25809
rect 12990 25735 13046 25744
rect 13096 25226 13124 27270
rect 13372 26994 13400 39520
rect 13634 36680 13690 36689
rect 13634 36615 13690 36624
rect 13450 35048 13506 35057
rect 13450 34983 13506 34992
rect 13464 34542 13492 34983
rect 13648 34746 13676 36615
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 13452 34536 13504 34542
rect 13452 34478 13504 34484
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13556 32881 13584 32914
rect 13542 32872 13598 32881
rect 13542 32807 13598 32816
rect 13556 32570 13584 32807
rect 13544 32564 13596 32570
rect 13544 32506 13596 32512
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 13556 26874 13584 32506
rect 13740 26926 13768 39520
rect 14200 37346 14228 39520
rect 13832 37318 14228 37346
rect 13832 34785 13860 37318
rect 14568 37210 14596 39520
rect 13924 37182 14596 37210
rect 13818 34776 13874 34785
rect 13818 34711 13874 34720
rect 13372 26846 13584 26874
rect 13728 26920 13780 26926
rect 13924 26897 13952 37182
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14936 31754 14964 39520
rect 15396 34649 15424 39520
rect 15382 34640 15438 34649
rect 15382 34575 15438 34584
rect 15764 32881 15792 39520
rect 15750 32872 15806 32881
rect 15750 32807 15806 32816
rect 14004 31748 14056 31754
rect 14004 31690 14056 31696
rect 14924 31748 14976 31754
rect 14924 31690 14976 31696
rect 14016 28966 14044 31690
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14004 28960 14056 28966
rect 14004 28902 14056 28908
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 13728 26862 13780 26868
rect 13910 26888 13966 26897
rect 13176 25356 13228 25362
rect 13176 25298 13228 25304
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 13096 24818 13124 25162
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13188 24682 13216 25298
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13004 23730 13032 24006
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12806 20904 12862 20913
rect 12806 20839 12862 20848
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12348 19168 12400 19174
rect 12268 19128 12348 19156
rect 12268 17814 12296 19128
rect 12348 19110 12400 19116
rect 12452 18290 12480 19790
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19378 12572 19654
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12438 18184 12494 18193
rect 12438 18119 12494 18128
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12360 17882 12388 18022
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12268 17338 12296 17614
rect 12452 17338 12480 18119
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 16674 12572 19314
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12636 18630 12664 19246
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18970 12756 19110
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12912 18086 12940 18294
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 13004 17678 13032 18566
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12728 16794 12756 17478
rect 12820 17270 12848 17478
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12820 17134 12848 17206
rect 13004 17202 13032 17614
rect 13096 17610 13124 18226
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12912 16697 12940 16934
rect 12898 16688 12954 16697
rect 12544 16646 12756 16674
rect 12254 15056 12310 15065
rect 12254 14991 12310 15000
rect 12072 9998 12124 10004
rect 12162 10024 12218 10033
rect 12084 9722 12112 9998
rect 12162 9959 12218 9968
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11978 8392 12034 8401
rect 11978 8327 12034 8336
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11532 7342 11560 7686
rect 11992 7546 12020 7890
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11426 7032 11482 7041
rect 11426 6967 11482 6976
rect 11532 6882 11560 7278
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11532 6854 11652 6882
rect 11348 6820 11468 6848
rect 11256 6718 11376 6746
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11256 6118 11284 6598
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 10690 5944 10746 5953
rect 10690 5879 10692 5888
rect 10744 5879 10746 5888
rect 10692 5850 10744 5856
rect 10704 5302 10732 5850
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10796 5370 10824 5646
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10692 5296 10744 5302
rect 10796 5273 10824 5306
rect 10692 5238 10744 5244
rect 10782 5264 10838 5273
rect 10782 5199 10838 5208
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10612 4282 10640 4762
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10704 4214 10732 4966
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10796 4282 10824 4626
rect 10888 4622 10916 5646
rect 11164 5642 11192 6054
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11072 4690 11100 5578
rect 11256 4826 11284 6054
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10336 3726 10456 3754
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10336 610 10364 3726
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10428 3194 10456 3470
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10428 2825 10456 3130
rect 10414 2816 10470 2825
rect 10414 2751 10470 2760
rect 10704 2582 10732 3470
rect 10796 2650 10824 4014
rect 10888 3534 10916 4558
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10980 3466 11008 4558
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 3505 11100 3878
rect 11058 3496 11114 3505
rect 10968 3460 11020 3466
rect 11058 3431 11114 3440
rect 10968 3402 11020 3408
rect 11348 3194 11376 6718
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 10968 3120 11020 3126
rect 11060 3120 11112 3126
rect 10968 3062 11020 3068
rect 11058 3088 11060 3097
rect 11112 3088 11114 3097
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10324 604 10376 610
rect 10324 546 10376 552
rect 10600 604 10652 610
rect 10600 546 10652 552
rect 10612 480 10640 546
rect 10980 480 11008 3062
rect 11058 3023 11114 3032
rect 11244 2984 11296 2990
rect 11348 2972 11376 3130
rect 11296 2944 11376 2972
rect 11244 2926 11296 2932
rect 11440 2836 11468 6820
rect 11624 6662 11652 6854
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11520 6112 11572 6118
rect 11624 6100 11652 6598
rect 11716 6458 11744 6802
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11572 6072 11652 6100
rect 11520 6054 11572 6060
rect 11532 5794 11560 6054
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11532 5766 11652 5794
rect 11992 5778 12020 6122
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 4049 11560 5510
rect 11624 5166 11652 5766
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 5370 12020 5714
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11886 4312 11942 4321
rect 11886 4247 11888 4256
rect 11940 4247 11942 4256
rect 11888 4218 11940 4224
rect 11992 4078 12020 4422
rect 12084 4146 12112 9318
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11980 4072 12032 4078
rect 11518 4040 11574 4049
rect 11980 4014 12032 4020
rect 11518 3975 11574 3984
rect 11992 3942 12020 4014
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11992 3670 12020 3878
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11624 3233 11652 3470
rect 11610 3224 11666 3233
rect 11610 3159 11666 3168
rect 11164 2808 11468 2836
rect 11164 2666 11192 2808
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11164 2638 11376 2666
rect 11992 2650 12020 3606
rect 12268 3505 12296 14991
rect 12346 14240 12402 14249
rect 12346 14175 12402 14184
rect 12360 11234 12388 14175
rect 12530 12744 12586 12753
rect 12530 12679 12586 12688
rect 12544 11626 12572 12679
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12636 11286 12664 11834
rect 12624 11280 12676 11286
rect 12360 11206 12480 11234
rect 12728 11257 12756 16646
rect 12898 16623 12954 16632
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 11354 12848 11494
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12624 11222 12676 11228
rect 12714 11248 12770 11257
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12360 10266 12388 11018
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12452 10130 12480 11206
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12544 10674 12572 11154
rect 12636 10792 12664 11222
rect 12714 11183 12770 11192
rect 12716 10804 12768 10810
rect 12636 10764 12716 10792
rect 12716 10746 12768 10752
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12360 9654 12388 10066
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12360 8945 12388 9590
rect 12346 8936 12402 8945
rect 12346 8871 12402 8880
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5681 12480 6054
rect 12530 5808 12586 5817
rect 12530 5743 12586 5752
rect 12438 5672 12494 5681
rect 12348 5636 12400 5642
rect 12438 5607 12494 5616
rect 12348 5578 12400 5584
rect 12360 4282 12388 5578
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12452 4078 12480 4558
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12254 3496 12310 3505
rect 12254 3431 12310 3440
rect 11348 480 11376 2638
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11794 2544 11850 2553
rect 11794 2479 11850 2488
rect 11808 480 11836 2479
rect 12360 610 12388 3878
rect 12164 604 12216 610
rect 12164 546 12216 552
rect 12348 604 12400 610
rect 12348 546 12400 552
rect 12176 480 12204 546
rect 12544 480 12572 5743
rect 12636 5370 12664 7142
rect 12728 6882 12756 10746
rect 12912 7478 12940 16390
rect 13084 13184 13136 13190
rect 13082 13152 13084 13161
rect 13136 13152 13138 13161
rect 13082 13087 13138 13096
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11762 13032 12038
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11082 13032 11494
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 13096 10198 13124 12378
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13188 7857 13216 24618
rect 13372 15609 13400 26846
rect 13910 26823 13966 26832
rect 13542 25800 13598 25809
rect 13542 25735 13598 25744
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13464 21486 13492 21830
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13556 19718 13584 25735
rect 13924 25362 13952 26823
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 13912 25356 13964 25362
rect 13912 25298 13964 25304
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13634 23352 13690 23361
rect 13634 23287 13690 23296
rect 13648 21690 13676 23287
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13358 15600 13414 15609
rect 13358 15535 13414 15544
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 13870 13308 14418
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13174 7848 13230 7857
rect 13174 7783 13230 7792
rect 13280 7546 13308 13806
rect 13372 11898 13400 15535
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12820 7002 12848 7346
rect 12898 7304 12954 7313
rect 12898 7239 12900 7248
rect 12952 7239 12954 7248
rect 12900 7210 12952 7216
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12728 6854 12940 6882
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12728 5098 12756 5510
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12728 3194 12756 5034
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12820 2650 12848 4966
rect 12912 4690 12940 6854
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12912 4146 12940 4490
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 13096 2650 13124 5646
rect 13188 5642 13216 6190
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13188 5234 13216 5578
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13188 3738 13216 5170
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13280 610 13308 7346
rect 12992 604 13044 610
rect 12992 546 13044 552
rect 13268 604 13320 610
rect 13268 546 13320 552
rect 13004 480 13032 546
rect 13372 480 13400 11562
rect 13464 10985 13492 18906
rect 13542 16688 13598 16697
rect 13542 16623 13598 16632
rect 13556 14550 13584 16623
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13450 10976 13506 10985
rect 13450 10911 13506 10920
rect 13464 10713 13492 10911
rect 13450 10704 13506 10713
rect 13450 10639 13506 10648
rect 13740 9194 13768 24550
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 15382 10704 15438 10713
rect 15382 10639 15438 10648
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 13464 9166 13768 9194
rect 13464 5234 13492 9166
rect 13726 9072 13782 9081
rect 13726 9007 13782 9016
rect 13634 7848 13690 7857
rect 13634 7783 13690 7792
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13464 4282 13492 4626
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13556 4185 13584 4422
rect 13542 4176 13598 4185
rect 13452 4140 13504 4146
rect 13542 4111 13598 4120
rect 13452 4082 13504 4088
rect 13464 3058 13492 4082
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13464 2854 13492 2994
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13464 2446 13492 2790
rect 13648 2582 13676 7783
rect 13740 5522 13768 9007
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 13740 5494 14228 5522
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13740 4049 13768 5170
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 13740 2922 13768 3975
rect 13818 3224 13874 3233
rect 13818 3159 13874 3168
rect 13832 2990 13860 3159
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13832 2650 13860 2926
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13726 2000 13782 2009
rect 13726 1935 13782 1944
rect 13740 480 13768 1935
rect 14200 480 14228 5494
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14646 4040 14702 4049
rect 14646 3975 14702 3984
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 1986 14688 3975
rect 14922 2408 14978 2417
rect 14922 2343 14978 2352
rect 14568 1958 14688 1986
rect 14568 480 14596 1958
rect 14936 480 14964 2343
rect 15396 480 15424 10639
rect 15750 8936 15806 8945
rect 15750 8871 15806 8880
rect 15764 480 15792 8871
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 2042 35128 2098 35184
rect 1490 34856 1546 34912
rect 1950 33088 2006 33144
rect 1674 32952 1730 33008
rect 2410 32952 2466 33008
rect 3146 38936 3202 38992
rect 2594 32272 2650 32328
rect 1674 31184 1730 31240
rect 1582 30912 1638 30968
rect 1398 27920 1454 27976
rect 1674 28872 1730 28928
rect 1582 26968 1638 27024
rect 1490 24928 1546 24984
rect 2226 30776 2282 30832
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3422 36896 3478 36952
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3422 34992 3478 35048
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 4526 35808 4582 35864
rect 4434 35128 4490 35184
rect 3238 33496 3294 33552
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3422 33496 3478 33552
rect 2410 28076 2466 28112
rect 2410 28056 2412 28076
rect 2412 28056 2464 28076
rect 2464 28056 2466 28076
rect 2226 25644 2228 25664
rect 2228 25644 2280 25664
rect 2280 25644 2282 25664
rect 2226 25608 2282 25644
rect 1766 23024 1822 23080
rect 2318 22888 2374 22944
rect 1674 20984 1730 21040
rect 2410 21120 2466 21176
rect 1582 18944 1638 19000
rect 1398 17176 1454 17232
rect 1674 18300 1676 18320
rect 1676 18300 1728 18320
rect 1728 18300 1730 18320
rect 1674 18264 1730 18300
rect 1582 16904 1638 16960
rect 1674 14864 1730 14920
rect 1582 12960 1638 13016
rect 1398 12300 1454 12336
rect 1398 12280 1400 12300
rect 1400 12280 1452 12300
rect 1452 12280 1454 12300
rect 1766 13912 1822 13968
rect 2410 14864 2466 14920
rect 2594 14320 2650 14376
rect 2042 12280 2098 12336
rect 2594 13232 2650 13288
rect 1582 10920 1638 10976
rect 1582 8880 1638 8936
rect 2318 6976 2374 7032
rect 570 5616 626 5672
rect 202 4120 258 4176
rect 1582 4936 1638 4992
rect 1766 3712 1822 3768
rect 1674 3576 1730 3632
rect 1950 2916 2006 2952
rect 1950 2896 1952 2916
rect 1952 2896 2004 2916
rect 2004 2896 2006 2916
rect 2502 6060 2504 6080
rect 2504 6060 2556 6080
rect 2556 6060 2558 6080
rect 2502 6024 2558 6060
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 4066 29552 4122 29608
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 2870 20848 2926 20904
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 5354 34584 5410 34640
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6918 34584 6974 34640
rect 7470 34584 7526 34640
rect 4434 29552 4490 29608
rect 4618 29008 4674 29064
rect 4434 21140 4490 21176
rect 4434 21120 4436 21140
rect 4436 21120 4488 21140
rect 4488 21120 4490 21140
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3606 11736 3662 11792
rect 3146 11328 3202 11384
rect 3514 11192 3570 11248
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 4158 10104 4214 10160
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3054 8372 3056 8392
rect 3056 8372 3108 8392
rect 3108 8372 3110 8392
rect 3054 8336 3110 8372
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3330 7284 3332 7304
rect 3332 7284 3384 7304
rect 3384 7284 3386 7304
rect 3330 7248 3386 7284
rect 2962 7148 2964 7168
rect 2964 7148 3016 7168
rect 3016 7148 3018 7168
rect 2962 7112 3018 7148
rect 2778 6840 2834 6896
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3606 6332 3608 6352
rect 3608 6332 3660 6352
rect 3660 6332 3662 6352
rect 3606 6296 3662 6332
rect 2410 2644 2466 2680
rect 2410 2624 2412 2644
rect 2412 2624 2464 2644
rect 2464 2624 2466 2644
rect 2870 4564 2872 4584
rect 2872 4564 2924 4584
rect 2924 4564 2926 4584
rect 2870 4528 2926 4564
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3146 4120 3202 4176
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3330 4120 3386 4176
rect 2686 2760 2742 2816
rect 4526 13404 4528 13424
rect 4528 13404 4580 13424
rect 4580 13404 4582 13424
rect 4526 13368 4582 13404
rect 4434 13232 4490 13288
rect 4986 29552 5042 29608
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6090 33360 6146 33416
rect 5814 33088 5870 33144
rect 5814 29280 5870 29336
rect 5078 27104 5134 27160
rect 4986 24656 5042 24712
rect 4802 20848 4858 20904
rect 4986 20304 5042 20360
rect 4710 15952 4766 16008
rect 4710 12416 4766 12472
rect 4342 7384 4398 7440
rect 4250 5636 4306 5672
rect 4250 5616 4252 5636
rect 4252 5616 4304 5636
rect 4304 5616 4306 5636
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 4250 3168 4306 3224
rect 3974 3032 4030 3088
rect 3514 2896 3570 2952
rect 2594 1400 2650 1456
rect 2502 992 2558 1048
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 4526 3440 4582 3496
rect 4342 2760 4398 2816
rect 5170 25608 5226 25664
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6826 33108 6882 33144
rect 6826 33088 6828 33108
rect 6828 33088 6880 33108
rect 6880 33088 6882 33108
rect 6918 32952 6974 33008
rect 8482 35828 8538 35864
rect 8482 35808 8484 35828
rect 8484 35808 8536 35828
rect 8536 35808 8538 35828
rect 6918 31728 6974 31784
rect 7470 32272 7526 32328
rect 6734 30912 6790 30968
rect 5814 28600 5870 28656
rect 5538 23160 5594 23216
rect 5538 22516 5540 22536
rect 5540 22516 5592 22536
rect 5592 22516 5594 22536
rect 5538 22480 5594 22516
rect 5630 18808 5686 18864
rect 5354 18672 5410 18728
rect 5538 18148 5594 18184
rect 5538 18128 5540 18148
rect 5540 18128 5592 18148
rect 5592 18128 5594 18148
rect 5446 16088 5502 16144
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6274 29180 6276 29200
rect 6276 29180 6328 29200
rect 6328 29180 6330 29200
rect 6274 29144 6330 29180
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6734 27532 6790 27568
rect 6734 27512 6736 27532
rect 6736 27512 6788 27532
rect 6788 27512 6790 27532
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6182 23160 6238 23216
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6366 19916 6422 19952
rect 6366 19896 6368 19916
rect 6368 19896 6420 19916
rect 6420 19896 6422 19916
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 7102 30640 7158 30696
rect 7562 32136 7618 32192
rect 7838 33088 7894 33144
rect 7746 32000 7802 32056
rect 7010 27920 7066 27976
rect 7562 30776 7618 30832
rect 7654 29844 7710 29880
rect 7654 29824 7656 29844
rect 7656 29824 7708 29844
rect 7708 29824 7710 29844
rect 7654 29588 7656 29608
rect 7656 29588 7708 29608
rect 7708 29588 7710 29608
rect 7654 29552 7710 29588
rect 7102 24520 7158 24576
rect 7286 26852 7342 26888
rect 7286 26832 7288 26852
rect 7288 26832 7340 26852
rect 7340 26832 7342 26852
rect 7286 25764 7342 25800
rect 7286 25744 7288 25764
rect 7288 25744 7340 25764
rect 7340 25744 7342 25764
rect 7286 24792 7342 24848
rect 7010 19216 7066 19272
rect 6642 18808 6698 18864
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6734 18028 6736 18048
rect 6736 18028 6788 18048
rect 6788 18028 6790 18048
rect 6734 17992 6790 18028
rect 6642 16496 6698 16552
rect 5722 15136 5778 15192
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 4710 6196 4712 6216
rect 4712 6196 4764 6216
rect 4764 6196 4766 6216
rect 4710 6160 4766 6196
rect 5170 11192 5226 11248
rect 5170 9152 5226 9208
rect 5814 12280 5870 12336
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 5906 11348 5962 11384
rect 5906 11328 5908 11348
rect 5908 11328 5960 11348
rect 5960 11328 5962 11348
rect 5998 11192 6054 11248
rect 5906 9288 5962 9344
rect 5630 7112 5686 7168
rect 4710 3304 4766 3360
rect 5078 2624 5134 2680
rect 5262 5616 5318 5672
rect 5354 4392 5410 4448
rect 5906 6840 5962 6896
rect 5722 5092 5778 5128
rect 5722 5072 5724 5092
rect 5724 5072 5776 5092
rect 5776 5072 5778 5092
rect 5630 4256 5686 4312
rect 5722 3712 5778 3768
rect 5262 1944 5318 2000
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6090 9288 6146 9344
rect 6458 9596 6460 9616
rect 6460 9596 6512 9616
rect 6512 9596 6514 9616
rect 6458 9560 6514 9596
rect 6826 14320 6882 14376
rect 7102 18300 7104 18320
rect 7104 18300 7156 18320
rect 7156 18300 7158 18320
rect 7102 18264 7158 18300
rect 7102 14864 7158 14920
rect 7562 25200 7618 25256
rect 7470 20440 7526 20496
rect 8666 34584 8722 34640
rect 8482 34448 8538 34504
rect 8206 30912 8262 30968
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 9310 34448 9366 34504
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 9678 34720 9734 34776
rect 9678 33360 9734 33416
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8850 32408 8906 32464
rect 9494 32680 9550 32736
rect 8666 32136 8722 32192
rect 8666 29300 8722 29336
rect 8666 29280 8668 29300
rect 8668 29280 8720 29300
rect 8720 29280 8722 29300
rect 8390 29144 8446 29200
rect 8114 27820 8116 27840
rect 8116 27820 8168 27840
rect 8168 27820 8170 27840
rect 8114 27784 8170 27820
rect 8298 27512 8354 27568
rect 7930 26732 7932 26752
rect 7932 26732 7984 26752
rect 7984 26732 7986 26752
rect 7930 26696 7986 26732
rect 7838 24520 7894 24576
rect 7930 22208 7986 22264
rect 7746 17584 7802 17640
rect 7838 15000 7894 15056
rect 7746 14764 7748 14784
rect 7748 14764 7800 14784
rect 7800 14764 7802 14784
rect 7746 14728 7802 14764
rect 7194 14320 7250 14376
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6090 6024 6146 6080
rect 5906 5072 5962 5128
rect 6090 4664 6146 4720
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 7010 6296 7066 6352
rect 7010 5888 7066 5944
rect 7194 5616 7250 5672
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6366 4120 6422 4176
rect 6274 4020 6276 4040
rect 6276 4020 6328 4040
rect 6328 4020 6330 4040
rect 6274 3984 6330 4020
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 7470 7792 7526 7848
rect 7838 13252 7894 13288
rect 7838 13232 7840 13252
rect 7840 13232 7892 13252
rect 7892 13232 7894 13252
rect 7562 5888 7618 5944
rect 7378 5208 7434 5264
rect 7286 4428 7288 4448
rect 7288 4428 7340 4448
rect 7340 4428 7342 4448
rect 7286 4392 7342 4428
rect 7470 4548 7526 4584
rect 7470 4528 7472 4548
rect 7472 4528 7524 4548
rect 7524 4528 7526 4548
rect 8666 29008 8722 29064
rect 8206 25336 8262 25392
rect 8298 23160 8354 23216
rect 8206 21428 8208 21448
rect 8208 21428 8260 21448
rect 8260 21428 8262 21448
rect 8206 21392 8262 21428
rect 8114 18672 8170 18728
rect 8574 27124 8630 27160
rect 8574 27104 8576 27124
rect 8576 27104 8628 27124
rect 8628 27104 8630 27124
rect 8574 26560 8630 26616
rect 9310 32000 9366 32056
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8850 29008 8906 29064
rect 9218 28464 9274 28520
rect 8758 21392 8814 21448
rect 8206 18128 8262 18184
rect 8574 19216 8630 19272
rect 8390 16496 8446 16552
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 9402 27920 9458 27976
rect 9678 32408 9734 32464
rect 9954 34484 9956 34504
rect 9956 34484 10008 34504
rect 10008 34484 10010 34504
rect 9954 34448 10010 34484
rect 9862 33496 9918 33552
rect 10322 35128 10378 35184
rect 10598 34312 10654 34368
rect 10046 32000 10102 32056
rect 9678 30660 9734 30696
rect 9678 30640 9680 30660
rect 9680 30640 9732 30660
rect 9732 30640 9734 30660
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 9678 27784 9734 27840
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8942 24692 8944 24712
rect 8944 24692 8996 24712
rect 8996 24692 8998 24712
rect 8942 24656 8998 24692
rect 9310 24656 9366 24712
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8482 15564 8538 15600
rect 8482 15544 8484 15564
rect 8484 15544 8536 15564
rect 8536 15544 8538 15564
rect 8390 14728 8446 14784
rect 8022 13776 8078 13832
rect 8206 9288 8262 9344
rect 9310 18128 9366 18184
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8666 12688 8722 12744
rect 8482 10104 8538 10160
rect 7746 6160 7802 6216
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 9862 26560 9918 26616
rect 10506 31728 10562 31784
rect 10874 34584 10930 34640
rect 10414 31184 10470 31240
rect 10230 26696 10286 26752
rect 10046 25220 10102 25256
rect 10046 25200 10048 25220
rect 10048 25200 10100 25220
rect 10100 25200 10102 25220
rect 10966 31340 11022 31376
rect 10966 31320 10968 31340
rect 10968 31320 11020 31340
rect 11020 31320 11022 31340
rect 10598 29144 10654 29200
rect 10322 24792 10378 24848
rect 10322 24556 10324 24576
rect 10324 24556 10376 24576
rect 10376 24556 10378 24576
rect 10322 24520 10378 24556
rect 9678 22228 9734 22264
rect 9678 22208 9680 22228
rect 9680 22208 9732 22228
rect 9732 22208 9734 22228
rect 9954 22480 10010 22536
rect 9954 20440 10010 20496
rect 9862 20304 9918 20360
rect 9954 20168 10010 20224
rect 9862 18828 9918 18864
rect 9862 18808 9864 18828
rect 9864 18808 9916 18828
rect 9916 18808 9918 18828
rect 9862 18672 9918 18728
rect 9770 18400 9826 18456
rect 9678 16088 9734 16144
rect 9678 14728 9734 14784
rect 9586 14184 9642 14240
rect 9678 13640 9734 13696
rect 9678 12280 9734 12336
rect 9494 11736 9550 11792
rect 9402 10920 9458 10976
rect 9402 9832 9458 9888
rect 9402 9696 9458 9752
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8666 7384 8722 7440
rect 8390 7112 8446 7168
rect 8298 6976 8354 7032
rect 7930 5616 7986 5672
rect 7746 4120 7802 4176
rect 7654 2760 7710 2816
rect 7102 1400 7158 1456
rect 8022 3984 8078 4040
rect 7930 2760 7986 2816
rect 10138 18944 10194 19000
rect 10322 17176 10378 17232
rect 10506 23044 10562 23080
rect 10506 23024 10508 23044
rect 10508 23024 10560 23044
rect 10560 23024 10562 23044
rect 10782 22480 10838 22536
rect 10690 18572 10692 18592
rect 10692 18572 10744 18592
rect 10744 18572 10746 18592
rect 10690 18536 10746 18572
rect 10598 18164 10600 18184
rect 10600 18164 10652 18184
rect 10652 18164 10654 18184
rect 10598 18128 10654 18164
rect 10690 17584 10746 17640
rect 11334 32172 11336 32192
rect 11336 32172 11388 32192
rect 11388 32172 11390 32192
rect 11334 32136 11390 32172
rect 11426 27532 11482 27568
rect 11426 27512 11428 27532
rect 11428 27512 11480 27532
rect 11480 27512 11482 27532
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 12162 32816 12218 32872
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 12346 32680 12402 32736
rect 12162 29960 12218 30016
rect 12162 28056 12218 28112
rect 12162 27920 12218 27976
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11242 18400 11298 18456
rect 10414 16632 10470 16688
rect 10598 15972 10654 16008
rect 10598 15952 10600 15972
rect 10600 15952 10652 15972
rect 10652 15952 10654 15972
rect 10230 14456 10286 14512
rect 10046 14320 10102 14376
rect 10230 13232 10286 13288
rect 10046 12588 10048 12608
rect 10048 12588 10100 12608
rect 10100 12588 10102 12608
rect 10046 12552 10102 12588
rect 10138 12280 10194 12336
rect 10046 9560 10102 9616
rect 9862 9324 9864 9344
rect 9864 9324 9916 9344
rect 9916 9324 9918 9344
rect 9862 9288 9918 9324
rect 10782 13368 10838 13424
rect 10414 12416 10470 12472
rect 10322 11736 10378 11792
rect 10506 11736 10562 11792
rect 9678 8336 9734 8392
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 9218 7420 9220 7440
rect 9220 7420 9272 7440
rect 9272 7420 9274 7440
rect 9218 7384 9274 7420
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 9402 6976 9458 7032
rect 9678 7148 9680 7168
rect 9680 7148 9732 7168
rect 9732 7148 9734 7168
rect 9678 7112 9734 7148
rect 9402 5752 9458 5808
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8482 3304 8538 3360
rect 8298 3032 8354 3088
rect 8482 2760 8538 2816
rect 8482 2352 8538 2408
rect 9310 3576 9366 3632
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9126 2896 9182 2952
rect 8850 2760 8906 2816
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9862 4664 9918 4720
rect 9678 2896 9734 2952
rect 9494 2760 9550 2816
rect 10046 2896 10102 2952
rect 10506 7248 10562 7304
rect 10414 5752 10470 5808
rect 10414 5072 10470 5128
rect 10230 4528 10286 4584
rect 10322 3848 10378 3904
rect 10782 12416 10838 12472
rect 11150 13096 11206 13152
rect 10782 12008 10838 12064
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 12070 25336 12126 25392
rect 12806 31320 12862 31376
rect 12070 18400 12126 18456
rect 11334 12008 11390 12064
rect 11058 9696 11114 9752
rect 11242 9832 11298 9888
rect 10782 7248 10838 7304
rect 11978 12280 12034 12336
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 12530 21392 12586 21448
rect 12990 25744 13046 25800
rect 13634 36624 13690 36680
rect 13450 34992 13506 35048
rect 13542 32816 13598 32872
rect 13818 34720 13874 34776
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 15382 34584 15438 34640
rect 15750 32816 15806 32872
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 12806 20848 12862 20904
rect 12438 18128 12494 18184
rect 12254 15000 12310 15056
rect 12162 9968 12218 10024
rect 11978 8336 12034 8392
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11426 6976 11482 7032
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 10690 5908 10746 5944
rect 10690 5888 10692 5908
rect 10692 5888 10744 5908
rect 10744 5888 10746 5908
rect 10782 5208 10838 5264
rect 10414 2760 10470 2816
rect 11058 3440 11114 3496
rect 11058 3068 11060 3088
rect 11060 3068 11112 3088
rect 11112 3068 11114 3088
rect 11058 3032 11114 3068
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11886 4276 11942 4312
rect 11886 4256 11888 4276
rect 11888 4256 11940 4276
rect 11940 4256 11942 4276
rect 11518 3984 11574 4040
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11610 3168 11666 3224
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12346 14184 12402 14240
rect 12530 12688 12586 12744
rect 12898 16632 12954 16688
rect 12714 11192 12770 11248
rect 12346 8880 12402 8936
rect 12530 5752 12586 5808
rect 12438 5616 12494 5672
rect 12254 3440 12310 3496
rect 11794 2488 11850 2544
rect 13082 13132 13084 13152
rect 13084 13132 13136 13152
rect 13136 13132 13138 13152
rect 13082 13096 13138 13132
rect 13910 26832 13966 26888
rect 13542 25744 13598 25800
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 13634 23296 13690 23352
rect 13358 15544 13414 15600
rect 13174 7792 13230 7848
rect 12898 7268 12954 7304
rect 12898 7248 12900 7268
rect 12900 7248 12952 7268
rect 12952 7248 12954 7268
rect 13542 16632 13598 16688
rect 13450 10920 13506 10976
rect 13450 10648 13506 10704
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 15382 10648 15438 10704
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 13726 9016 13782 9072
rect 13634 7792 13690 7848
rect 13542 4120 13598 4176
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 13726 3984 13782 4040
rect 13818 3168 13874 3224
rect 13726 1944 13782 2000
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14646 3984 14702 4040
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 14922 2352 14978 2408
rect 15750 8880 15806 8936
<< metal3 >>
rect 0 38994 480 39024
rect 3141 38994 3207 38997
rect 0 38992 3207 38994
rect 0 38936 3146 38992
rect 3202 38936 3207 38992
rect 0 38934 3207 38936
rect 0 38904 480 38934
rect 3141 38931 3207 38934
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 0 36954 480 36984
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 3417 36954 3483 36957
rect 0 36952 3483 36954
rect 0 36896 3422 36952
rect 3478 36896 3483 36952
rect 0 36894 3483 36896
rect 0 36864 480 36894
rect 3417 36891 3483 36894
rect 13629 36682 13695 36685
rect 15520 36682 16000 36712
rect 13629 36680 16000 36682
rect 13629 36624 13634 36680
rect 13690 36624 16000 36680
rect 13629 36622 16000 36624
rect 13629 36619 13695 36622
rect 15520 36592 16000 36622
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 4521 35866 4587 35869
rect 8477 35866 8543 35869
rect 4521 35864 8543 35866
rect 4521 35808 4526 35864
rect 4582 35808 8482 35864
rect 8538 35808 8543 35864
rect 4521 35806 8543 35808
rect 4521 35803 4587 35806
rect 8477 35803 8543 35806
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 2037 35186 2103 35189
rect 4429 35186 4495 35189
rect 10317 35186 10383 35189
rect 2037 35184 10383 35186
rect 2037 35128 2042 35184
rect 2098 35128 4434 35184
rect 4490 35128 10322 35184
rect 10378 35128 10383 35184
rect 2037 35126 10383 35128
rect 2037 35123 2103 35126
rect 4429 35123 4495 35126
rect 10317 35123 10383 35126
rect 3417 35050 3483 35053
rect 13445 35050 13511 35053
rect 3417 35048 13511 35050
rect 3417 34992 3422 35048
rect 3478 34992 13450 35048
rect 13506 34992 13511 35048
rect 3417 34990 13511 34992
rect 3417 34987 3483 34990
rect 13445 34987 13511 34990
rect 0 34914 480 34944
rect 1485 34914 1551 34917
rect 0 34912 1551 34914
rect 0 34856 1490 34912
rect 1546 34856 1551 34912
rect 0 34854 1551 34856
rect 0 34824 480 34854
rect 1485 34851 1551 34854
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 9673 34778 9739 34781
rect 13813 34778 13879 34781
rect 9673 34776 13879 34778
rect 9673 34720 9678 34776
rect 9734 34720 13818 34776
rect 13874 34720 13879 34776
rect 9673 34718 13879 34720
rect 9673 34715 9739 34718
rect 13813 34715 13879 34718
rect 5349 34642 5415 34645
rect 6913 34642 6979 34645
rect 5349 34640 6979 34642
rect 5349 34584 5354 34640
rect 5410 34584 6918 34640
rect 6974 34584 6979 34640
rect 5349 34582 6979 34584
rect 5349 34579 5415 34582
rect 6913 34579 6979 34582
rect 7465 34642 7531 34645
rect 8661 34642 8727 34645
rect 7465 34640 8727 34642
rect 7465 34584 7470 34640
rect 7526 34584 8666 34640
rect 8722 34584 8727 34640
rect 7465 34582 8727 34584
rect 7465 34579 7531 34582
rect 8661 34579 8727 34582
rect 10869 34642 10935 34645
rect 15377 34642 15443 34645
rect 10869 34640 15443 34642
rect 10869 34584 10874 34640
rect 10930 34584 15382 34640
rect 15438 34584 15443 34640
rect 10869 34582 15443 34584
rect 10869 34579 10935 34582
rect 15377 34579 15443 34582
rect 8477 34506 8543 34509
rect 9305 34506 9371 34509
rect 9949 34506 10015 34509
rect 8477 34504 10015 34506
rect 8477 34448 8482 34504
rect 8538 34448 9310 34504
rect 9366 34448 9954 34504
rect 10010 34448 10015 34504
rect 8477 34446 10015 34448
rect 8477 34443 8543 34446
rect 9305 34443 9371 34446
rect 9949 34443 10015 34446
rect 8150 34308 8156 34372
rect 8220 34370 8226 34372
rect 10593 34370 10659 34373
rect 8220 34368 10659 34370
rect 8220 34312 10598 34368
rect 10654 34312 10659 34368
rect 8220 34310 10659 34312
rect 8220 34308 8226 34310
rect 10593 34307 10659 34310
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 3233 33554 3299 33557
rect 3417 33554 3483 33557
rect 9857 33554 9923 33557
rect 3233 33552 9923 33554
rect 3233 33496 3238 33552
rect 3294 33496 3422 33552
rect 3478 33496 9862 33552
rect 9918 33496 9923 33552
rect 3233 33494 9923 33496
rect 3233 33491 3299 33494
rect 3417 33491 3483 33494
rect 9857 33491 9923 33494
rect 6085 33418 6151 33421
rect 9673 33418 9739 33421
rect 6085 33416 9739 33418
rect 6085 33360 6090 33416
rect 6146 33360 9678 33416
rect 9734 33360 9739 33416
rect 6085 33358 9739 33360
rect 6085 33355 6151 33358
rect 9673 33355 9739 33358
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 1945 33146 2011 33149
rect 5809 33146 5875 33149
rect 1945 33144 5875 33146
rect 1945 33088 1950 33144
rect 2006 33088 5814 33144
rect 5870 33088 5875 33144
rect 1945 33086 5875 33088
rect 1945 33083 2011 33086
rect 5809 33083 5875 33086
rect 6821 33146 6887 33149
rect 7833 33146 7899 33149
rect 6821 33144 7899 33146
rect 6821 33088 6826 33144
rect 6882 33088 7838 33144
rect 7894 33088 7899 33144
rect 6821 33086 7899 33088
rect 6821 33083 6887 33086
rect 7833 33083 7899 33086
rect 0 33010 480 33040
rect 1669 33010 1735 33013
rect 0 33008 1735 33010
rect 0 32952 1674 33008
rect 1730 32952 1735 33008
rect 0 32950 1735 32952
rect 0 32920 480 32950
rect 1669 32947 1735 32950
rect 2405 33010 2471 33013
rect 6913 33010 6979 33013
rect 2405 33008 6979 33010
rect 2405 32952 2410 33008
rect 2466 32952 6918 33008
rect 6974 32952 6979 33008
rect 2405 32950 6979 32952
rect 2405 32947 2471 32950
rect 6913 32947 6979 32950
rect 12157 32874 12223 32877
rect 13537 32874 13603 32877
rect 15745 32874 15811 32877
rect 12157 32872 12266 32874
rect 12157 32816 12162 32872
rect 12218 32816 12266 32872
rect 12157 32811 12266 32816
rect 13537 32872 15811 32874
rect 13537 32816 13542 32872
rect 13598 32816 15750 32872
rect 15806 32816 15811 32872
rect 13537 32814 15811 32816
rect 13537 32811 13603 32814
rect 15745 32811 15811 32814
rect 9489 32738 9555 32741
rect 12206 32738 12266 32811
rect 12341 32738 12407 32741
rect 9489 32736 12407 32738
rect 9489 32680 9494 32736
rect 9550 32680 12346 32736
rect 12402 32680 12407 32736
rect 9489 32678 12407 32680
rect 9489 32675 9555 32678
rect 12341 32675 12407 32678
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 8845 32466 8911 32469
rect 9673 32466 9739 32469
rect 8845 32464 9739 32466
rect 8845 32408 8850 32464
rect 8906 32408 9678 32464
rect 9734 32408 9739 32464
rect 8845 32406 9739 32408
rect 8845 32403 8911 32406
rect 9673 32403 9739 32406
rect 2589 32330 2655 32333
rect 7465 32330 7531 32333
rect 2589 32328 7531 32330
rect 2589 32272 2594 32328
rect 2650 32272 7470 32328
rect 7526 32272 7531 32328
rect 2589 32270 7531 32272
rect 2589 32267 2655 32270
rect 7465 32267 7531 32270
rect 7557 32194 7623 32197
rect 8661 32194 8727 32197
rect 11329 32194 11395 32197
rect 7557 32192 11395 32194
rect 7557 32136 7562 32192
rect 7618 32136 8666 32192
rect 8722 32136 11334 32192
rect 11390 32136 11395 32192
rect 7557 32134 11395 32136
rect 7557 32131 7623 32134
rect 8661 32131 8727 32134
rect 11329 32131 11395 32134
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 7741 32058 7807 32061
rect 9305 32058 9371 32061
rect 10041 32060 10107 32061
rect 7741 32056 9371 32058
rect 7741 32000 7746 32056
rect 7802 32000 9310 32056
rect 9366 32000 9371 32056
rect 7741 31998 9371 32000
rect 7741 31995 7807 31998
rect 9305 31995 9371 31998
rect 9990 31996 9996 32060
rect 10060 32058 10107 32060
rect 10060 32056 10152 32058
rect 10102 32000 10152 32056
rect 10060 31998 10152 32000
rect 10060 31996 10107 31998
rect 10041 31995 10107 31996
rect 6913 31786 6979 31789
rect 10501 31786 10567 31789
rect 6913 31784 10567 31786
rect 6913 31728 6918 31784
rect 6974 31728 10506 31784
rect 10562 31728 10567 31784
rect 6913 31726 10567 31728
rect 6913 31723 6979 31726
rect 10501 31723 10567 31726
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 10961 31378 11027 31381
rect 12801 31378 12867 31381
rect 10961 31376 12867 31378
rect 10961 31320 10966 31376
rect 11022 31320 12806 31376
rect 12862 31320 12867 31376
rect 10961 31318 12867 31320
rect 10961 31315 11027 31318
rect 12801 31315 12867 31318
rect 1669 31242 1735 31245
rect 10409 31242 10475 31245
rect 1669 31240 10475 31242
rect 1669 31184 1674 31240
rect 1730 31184 10414 31240
rect 10470 31184 10475 31240
rect 1669 31182 10475 31184
rect 1669 31179 1735 31182
rect 10409 31179 10475 31182
rect 6277 31040 6597 31041
rect 0 30970 480 31000
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 1577 30970 1643 30973
rect 0 30968 1643 30970
rect 0 30912 1582 30968
rect 1638 30912 1643 30968
rect 0 30910 1643 30912
rect 0 30880 480 30910
rect 1577 30907 1643 30910
rect 6729 30970 6795 30973
rect 8201 30970 8267 30973
rect 6729 30968 8267 30970
rect 6729 30912 6734 30968
rect 6790 30912 8206 30968
rect 8262 30912 8267 30968
rect 6729 30910 8267 30912
rect 6729 30907 6795 30910
rect 8201 30907 8267 30910
rect 2221 30834 2287 30837
rect 7557 30834 7623 30837
rect 2221 30832 7623 30834
rect 2221 30776 2226 30832
rect 2282 30776 7562 30832
rect 7618 30776 7623 30832
rect 2221 30774 7623 30776
rect 2221 30771 2287 30774
rect 7557 30771 7623 30774
rect 7097 30698 7163 30701
rect 9673 30698 9739 30701
rect 7097 30696 9739 30698
rect 7097 30640 7102 30696
rect 7158 30640 9678 30696
rect 9734 30640 9739 30696
rect 7097 30638 9739 30640
rect 7097 30635 7163 30638
rect 9673 30635 9739 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 12157 30018 12223 30021
rect 15520 30018 16000 30048
rect 12157 30016 16000 30018
rect 12157 29960 12162 30016
rect 12218 29960 16000 30016
rect 12157 29958 16000 29960
rect 12157 29955 12223 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 7649 29882 7715 29885
rect 8150 29882 8156 29884
rect 7649 29880 8156 29882
rect 7649 29824 7654 29880
rect 7710 29824 8156 29880
rect 7649 29822 8156 29824
rect 7649 29819 7715 29822
rect 8150 29820 8156 29822
rect 8220 29820 8226 29884
rect 4061 29610 4127 29613
rect 4429 29610 4495 29613
rect 4061 29608 4495 29610
rect 4061 29552 4066 29608
rect 4122 29552 4434 29608
rect 4490 29552 4495 29608
rect 4061 29550 4495 29552
rect 4061 29547 4127 29550
rect 4429 29547 4495 29550
rect 4981 29610 5047 29613
rect 7649 29610 7715 29613
rect 4981 29608 7715 29610
rect 4981 29552 4986 29608
rect 5042 29552 7654 29608
rect 7710 29552 7715 29608
rect 4981 29550 7715 29552
rect 4981 29547 5047 29550
rect 7649 29547 7715 29550
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 5809 29338 5875 29341
rect 8661 29338 8727 29341
rect 5809 29336 8727 29338
rect 5809 29280 5814 29336
rect 5870 29280 8666 29336
rect 8722 29280 8727 29336
rect 5809 29278 8727 29280
rect 5809 29275 5875 29278
rect 8661 29275 8727 29278
rect 6269 29202 6335 29205
rect 8385 29202 8451 29205
rect 10593 29202 10659 29205
rect 6269 29200 10659 29202
rect 6269 29144 6274 29200
rect 6330 29144 8390 29200
rect 8446 29144 10598 29200
rect 10654 29144 10659 29200
rect 6269 29142 10659 29144
rect 6269 29139 6335 29142
rect 8385 29139 8451 29142
rect 10593 29139 10659 29142
rect 4613 29066 4679 29069
rect 8661 29066 8727 29069
rect 8845 29066 8911 29069
rect 4613 29064 8911 29066
rect 4613 29008 4618 29064
rect 4674 29008 8666 29064
rect 8722 29008 8850 29064
rect 8906 29008 8911 29064
rect 4613 29006 8911 29008
rect 4613 29003 4679 29006
rect 8661 29003 8727 29006
rect 8845 29003 8911 29006
rect 9990 29004 9996 29068
rect 10060 29004 10066 29068
rect 0 28930 480 28960
rect 1669 28930 1735 28933
rect 9998 28932 10058 29004
rect 0 28928 1735 28930
rect 0 28872 1674 28928
rect 1730 28872 1735 28928
rect 0 28870 1735 28872
rect 0 28840 480 28870
rect 1669 28867 1735 28870
rect 9990 28868 9996 28932
rect 10060 28868 10066 28932
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 5809 28658 5875 28661
rect 6126 28658 6132 28660
rect 5809 28656 6132 28658
rect 5809 28600 5814 28656
rect 5870 28600 6132 28656
rect 5809 28598 6132 28600
rect 5809 28595 5875 28598
rect 6126 28596 6132 28598
rect 6196 28596 6202 28660
rect 9213 28522 9279 28525
rect 9438 28522 9444 28524
rect 9213 28520 9444 28522
rect 9213 28464 9218 28520
rect 9274 28464 9444 28520
rect 9213 28462 9444 28464
rect 9213 28459 9279 28462
rect 9438 28460 9444 28462
rect 9508 28460 9514 28524
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 2405 28114 2471 28117
rect 12157 28114 12223 28117
rect 2405 28112 12223 28114
rect 2405 28056 2410 28112
rect 2466 28056 12162 28112
rect 12218 28056 12223 28112
rect 2405 28054 12223 28056
rect 2405 28051 2471 28054
rect 12157 28051 12223 28054
rect 1393 27978 1459 27981
rect 7005 27978 7071 27981
rect 1393 27976 7071 27978
rect 1393 27920 1398 27976
rect 1454 27920 7010 27976
rect 7066 27920 7071 27976
rect 1393 27918 7071 27920
rect 1393 27915 1459 27918
rect 7005 27915 7071 27918
rect 9397 27978 9463 27981
rect 12157 27978 12223 27981
rect 9397 27976 12223 27978
rect 9397 27920 9402 27976
rect 9458 27920 12162 27976
rect 12218 27920 12223 27976
rect 9397 27918 12223 27920
rect 9397 27915 9463 27918
rect 12157 27915 12223 27918
rect 8109 27842 8175 27845
rect 9673 27842 9739 27845
rect 8109 27840 9739 27842
rect 8109 27784 8114 27840
rect 8170 27784 9678 27840
rect 9734 27784 9739 27840
rect 8109 27782 9739 27784
rect 8109 27779 8175 27782
rect 9673 27779 9739 27782
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 6729 27570 6795 27573
rect 8293 27570 8359 27573
rect 11421 27570 11487 27573
rect 6729 27568 11487 27570
rect 6729 27512 6734 27568
rect 6790 27512 8298 27568
rect 8354 27512 11426 27568
rect 11482 27512 11487 27568
rect 6729 27510 11487 27512
rect 6729 27507 6795 27510
rect 8293 27507 8359 27510
rect 11421 27507 11487 27510
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 5073 27162 5139 27165
rect 8569 27162 8635 27165
rect 5073 27160 8635 27162
rect 5073 27104 5078 27160
rect 5134 27104 8574 27160
rect 8630 27104 8635 27160
rect 5073 27102 8635 27104
rect 5073 27099 5139 27102
rect 8569 27099 8635 27102
rect 0 27026 480 27056
rect 1577 27026 1643 27029
rect 0 27024 1643 27026
rect 0 26968 1582 27024
rect 1638 26968 1643 27024
rect 0 26966 1643 26968
rect 0 26936 480 26966
rect 1577 26963 1643 26966
rect 7281 26890 7347 26893
rect 13905 26890 13971 26893
rect 7281 26888 13971 26890
rect 7281 26832 7286 26888
rect 7342 26832 13910 26888
rect 13966 26832 13971 26888
rect 7281 26830 13971 26832
rect 7281 26827 7347 26830
rect 13905 26827 13971 26830
rect 7925 26754 7991 26757
rect 10225 26754 10291 26757
rect 7925 26752 10291 26754
rect 7925 26696 7930 26752
rect 7986 26696 10230 26752
rect 10286 26696 10291 26752
rect 7925 26694 10291 26696
rect 7925 26691 7991 26694
rect 10225 26691 10291 26694
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 8569 26618 8635 26621
rect 9857 26618 9923 26621
rect 8569 26616 9923 26618
rect 8569 26560 8574 26616
rect 8630 26560 9862 26616
rect 9918 26560 9923 26616
rect 8569 26558 9923 26560
rect 8569 26555 8635 26558
rect 9857 26555 9923 26558
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 7281 25802 7347 25805
rect 12985 25802 13051 25805
rect 13537 25802 13603 25805
rect 7281 25800 13603 25802
rect 7281 25744 7286 25800
rect 7342 25744 12990 25800
rect 13046 25744 13542 25800
rect 13598 25744 13603 25800
rect 7281 25742 13603 25744
rect 7281 25739 7347 25742
rect 12985 25739 13051 25742
rect 13537 25739 13603 25742
rect 2221 25666 2287 25669
rect 5165 25666 5231 25669
rect 2221 25664 5231 25666
rect 2221 25608 2226 25664
rect 2282 25608 5170 25664
rect 5226 25608 5231 25664
rect 2221 25606 5231 25608
rect 2221 25603 2287 25606
rect 5165 25603 5231 25606
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 8201 25394 8267 25397
rect 12065 25394 12131 25397
rect 8201 25392 12131 25394
rect 8201 25336 8206 25392
rect 8262 25336 12070 25392
rect 12126 25336 12131 25392
rect 8201 25334 12131 25336
rect 8201 25331 8267 25334
rect 12065 25331 12131 25334
rect 7557 25258 7623 25261
rect 10041 25258 10107 25261
rect 7557 25256 10107 25258
rect 7557 25200 7562 25256
rect 7618 25200 10046 25256
rect 10102 25200 10107 25256
rect 7557 25198 10107 25200
rect 7557 25195 7623 25198
rect 10041 25195 10107 25198
rect 3610 25056 3930 25057
rect 0 24986 480 25016
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 1485 24986 1551 24989
rect 0 24984 1551 24986
rect 0 24928 1490 24984
rect 1546 24928 1551 24984
rect 0 24926 1551 24928
rect 0 24896 480 24926
rect 1485 24923 1551 24926
rect 7281 24850 7347 24853
rect 10317 24850 10383 24853
rect 7281 24848 10383 24850
rect 7281 24792 7286 24848
rect 7342 24792 10322 24848
rect 10378 24792 10383 24848
rect 7281 24790 10383 24792
rect 7281 24787 7347 24790
rect 10317 24787 10383 24790
rect 4981 24714 5047 24717
rect 8937 24714 9003 24717
rect 4981 24712 9003 24714
rect 4981 24656 4986 24712
rect 5042 24656 8942 24712
rect 8998 24656 9003 24712
rect 4981 24654 9003 24656
rect 4981 24651 5047 24654
rect 8937 24651 9003 24654
rect 9305 24714 9371 24717
rect 9438 24714 9444 24716
rect 9305 24712 9444 24714
rect 9305 24656 9310 24712
rect 9366 24656 9444 24712
rect 9305 24654 9444 24656
rect 9305 24651 9371 24654
rect 9438 24652 9444 24654
rect 9508 24652 9514 24716
rect 7097 24578 7163 24581
rect 7833 24578 7899 24581
rect 10317 24578 10383 24581
rect 7097 24576 10383 24578
rect 7097 24520 7102 24576
rect 7158 24520 7838 24576
rect 7894 24520 10322 24576
rect 10378 24520 10383 24576
rect 7097 24518 10383 24520
rect 7097 24515 7163 24518
rect 7833 24515 7899 24518
rect 10317 24515 10383 24518
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 13629 23354 13695 23357
rect 15520 23354 16000 23384
rect 13629 23352 16000 23354
rect 13629 23296 13634 23352
rect 13690 23296 16000 23352
rect 13629 23294 16000 23296
rect 13629 23291 13695 23294
rect 15520 23264 16000 23294
rect 5533 23218 5599 23221
rect 6177 23218 6243 23221
rect 8293 23218 8359 23221
rect 5533 23216 8359 23218
rect 5533 23160 5538 23216
rect 5594 23160 6182 23216
rect 6238 23160 8298 23216
rect 8354 23160 8359 23216
rect 5533 23158 8359 23160
rect 5533 23155 5599 23158
rect 6177 23155 6243 23158
rect 8293 23155 8359 23158
rect 1761 23082 1827 23085
rect 10501 23082 10567 23085
rect 1761 23080 10567 23082
rect 1761 23024 1766 23080
rect 1822 23024 10506 23080
rect 10562 23024 10567 23080
rect 1761 23022 10567 23024
rect 1761 23019 1827 23022
rect 10501 23019 10567 23022
rect 0 22946 480 22976
rect 2313 22946 2379 22949
rect 0 22944 2379 22946
rect 0 22888 2318 22944
rect 2374 22888 2379 22944
rect 0 22886 2379 22888
rect 0 22856 480 22886
rect 2313 22883 2379 22886
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 5533 22538 5599 22541
rect 9949 22538 10015 22541
rect 10777 22538 10843 22541
rect 5533 22536 10843 22538
rect 5533 22480 5538 22536
rect 5594 22480 9954 22536
rect 10010 22480 10782 22536
rect 10838 22480 10843 22536
rect 5533 22478 10843 22480
rect 5533 22475 5599 22478
rect 9949 22475 10015 22478
rect 10777 22475 10843 22478
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 7925 22266 7991 22269
rect 9673 22266 9739 22269
rect 7925 22264 9739 22266
rect 7925 22208 7930 22264
rect 7986 22208 9678 22264
rect 9734 22208 9739 22264
rect 7925 22206 9739 22208
rect 7925 22203 7991 22206
rect 9673 22203 9739 22206
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 8201 21450 8267 21453
rect 8753 21450 8819 21453
rect 12525 21450 12591 21453
rect 8201 21448 12591 21450
rect 8201 21392 8206 21448
rect 8262 21392 8758 21448
rect 8814 21392 12530 21448
rect 12586 21392 12591 21448
rect 8201 21390 12591 21392
rect 8201 21387 8267 21390
rect 8753 21387 8819 21390
rect 12525 21387 12591 21390
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 2405 21178 2471 21181
rect 4429 21178 4495 21181
rect 2405 21176 4495 21178
rect 2405 21120 2410 21176
rect 2466 21120 4434 21176
rect 4490 21120 4495 21176
rect 2405 21118 4495 21120
rect 2405 21115 2471 21118
rect 4429 21115 4495 21118
rect 0 21042 480 21072
rect 1669 21042 1735 21045
rect 0 21040 1735 21042
rect 0 20984 1674 21040
rect 1730 20984 1735 21040
rect 0 20982 1735 20984
rect 0 20952 480 20982
rect 1669 20979 1735 20982
rect 2865 20906 2931 20909
rect 4797 20906 4863 20909
rect 12801 20906 12867 20909
rect 2865 20904 12867 20906
rect 2865 20848 2870 20904
rect 2926 20848 4802 20904
rect 4858 20848 12806 20904
rect 12862 20848 12867 20904
rect 2865 20846 12867 20848
rect 2865 20843 2931 20846
rect 4797 20843 4863 20846
rect 12801 20843 12867 20846
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 7465 20498 7531 20501
rect 9949 20498 10015 20501
rect 7465 20496 10015 20498
rect 7465 20440 7470 20496
rect 7526 20440 9954 20496
rect 10010 20440 10015 20496
rect 7465 20438 10015 20440
rect 7465 20435 7531 20438
rect 9949 20435 10015 20438
rect 4981 20362 5047 20365
rect 9857 20362 9923 20365
rect 4981 20360 9923 20362
rect 4981 20304 4986 20360
rect 5042 20304 9862 20360
rect 9918 20304 9923 20360
rect 4981 20302 9923 20304
rect 4981 20299 5047 20302
rect 9857 20299 9923 20302
rect 9949 20228 10015 20229
rect 9949 20226 9996 20228
rect 9904 20224 9996 20226
rect 9904 20168 9954 20224
rect 9904 20166 9996 20168
rect 9949 20164 9996 20166
rect 10060 20164 10066 20228
rect 9949 20163 10015 20164
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 6126 19892 6132 19956
rect 6196 19954 6202 19956
rect 6361 19954 6427 19957
rect 6196 19952 6427 19954
rect 6196 19896 6366 19952
rect 6422 19896 6427 19952
rect 6196 19894 6427 19896
rect 6196 19892 6202 19894
rect 6361 19891 6427 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 7005 19274 7071 19277
rect 8569 19274 8635 19277
rect 7005 19272 8635 19274
rect 7005 19216 7010 19272
rect 7066 19216 8574 19272
rect 8630 19216 8635 19272
rect 7005 19214 8635 19216
rect 7005 19211 7071 19214
rect 8569 19211 8635 19214
rect 6277 19072 6597 19073
rect 0 19002 480 19032
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 1577 19002 1643 19005
rect 0 19000 1643 19002
rect 0 18944 1582 19000
rect 1638 18944 1643 19000
rect 0 18942 1643 18944
rect 0 18912 480 18942
rect 1577 18939 1643 18942
rect 9622 18940 9628 19004
rect 9692 19002 9698 19004
rect 10133 19002 10199 19005
rect 9692 19000 10199 19002
rect 9692 18944 10138 19000
rect 10194 18944 10199 19000
rect 9692 18942 10199 18944
rect 9692 18940 9698 18942
rect 10133 18939 10199 18942
rect 5625 18866 5691 18869
rect 6637 18866 6703 18869
rect 9857 18866 9923 18869
rect 5625 18864 9923 18866
rect 5625 18808 5630 18864
rect 5686 18808 6642 18864
rect 6698 18808 9862 18864
rect 9918 18808 9923 18864
rect 5625 18806 9923 18808
rect 5625 18803 5691 18806
rect 6637 18803 6703 18806
rect 9857 18803 9923 18806
rect 5349 18730 5415 18733
rect 8109 18730 8175 18733
rect 9857 18730 9923 18733
rect 5349 18728 9923 18730
rect 5349 18672 5354 18728
rect 5410 18672 8114 18728
rect 8170 18672 9862 18728
rect 9918 18672 9923 18728
rect 5349 18670 9923 18672
rect 5349 18667 5415 18670
rect 8109 18667 8175 18670
rect 9857 18667 9923 18670
rect 10542 18532 10548 18596
rect 10612 18594 10618 18596
rect 10685 18594 10751 18597
rect 10612 18592 10751 18594
rect 10612 18536 10690 18592
rect 10746 18536 10751 18592
rect 10612 18534 10751 18536
rect 10612 18532 10618 18534
rect 10685 18531 10751 18534
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 9765 18458 9831 18461
rect 11237 18458 11303 18461
rect 12065 18458 12131 18461
rect 9765 18456 12131 18458
rect 9765 18400 9770 18456
rect 9826 18400 11242 18456
rect 11298 18400 12070 18456
rect 12126 18400 12131 18456
rect 9765 18398 12131 18400
rect 9765 18395 9831 18398
rect 11237 18395 11303 18398
rect 12065 18395 12131 18398
rect 1669 18322 1735 18325
rect 7097 18322 7163 18325
rect 1669 18320 7163 18322
rect 1669 18264 1674 18320
rect 1730 18264 7102 18320
rect 7158 18264 7163 18320
rect 1669 18262 7163 18264
rect 1669 18259 1735 18262
rect 7097 18259 7163 18262
rect 5533 18186 5599 18189
rect 8201 18186 8267 18189
rect 9305 18186 9371 18189
rect 5533 18184 9371 18186
rect 5533 18128 5538 18184
rect 5594 18128 8206 18184
rect 8262 18128 9310 18184
rect 9366 18128 9371 18184
rect 5533 18126 9371 18128
rect 5533 18123 5599 18126
rect 8201 18123 8267 18126
rect 9305 18123 9371 18126
rect 10593 18186 10659 18189
rect 12433 18186 12499 18189
rect 10593 18184 12499 18186
rect 10593 18128 10598 18184
rect 10654 18128 12438 18184
rect 12494 18128 12499 18184
rect 10593 18126 12499 18128
rect 10593 18123 10659 18126
rect 12433 18123 12499 18126
rect 6729 18050 6795 18053
rect 10542 18050 10548 18052
rect 6729 18048 10548 18050
rect 6729 17992 6734 18048
rect 6790 17992 10548 18048
rect 6729 17990 10548 17992
rect 6729 17987 6795 17990
rect 10542 17988 10548 17990
rect 10612 17988 10618 18052
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 7741 17642 7807 17645
rect 10685 17642 10751 17645
rect 7741 17640 10751 17642
rect 7741 17584 7746 17640
rect 7802 17584 10690 17640
rect 10746 17584 10751 17640
rect 7741 17582 10751 17584
rect 7741 17579 7807 17582
rect 10685 17579 10751 17582
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 1393 17234 1459 17237
rect 10317 17234 10383 17237
rect 1393 17232 10383 17234
rect 1393 17176 1398 17232
rect 1454 17176 10322 17232
rect 10378 17176 10383 17232
rect 1393 17174 10383 17176
rect 1393 17171 1459 17174
rect 10317 17171 10383 17174
rect 0 16962 480 16992
rect 1577 16962 1643 16965
rect 0 16960 1643 16962
rect 0 16904 1582 16960
rect 1638 16904 1643 16960
rect 0 16902 1643 16904
rect 0 16872 480 16902
rect 1577 16899 1643 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 10409 16690 10475 16693
rect 12893 16690 12959 16693
rect 10409 16688 12959 16690
rect 10409 16632 10414 16688
rect 10470 16632 12898 16688
rect 12954 16632 12959 16688
rect 10409 16630 12959 16632
rect 10409 16627 10475 16630
rect 12893 16627 12959 16630
rect 13537 16690 13603 16693
rect 15520 16690 16000 16720
rect 13537 16688 16000 16690
rect 13537 16632 13542 16688
rect 13598 16632 16000 16688
rect 13537 16630 16000 16632
rect 13537 16627 13603 16630
rect 15520 16600 16000 16630
rect 6637 16554 6703 16557
rect 8385 16554 8451 16557
rect 6637 16552 8451 16554
rect 6637 16496 6642 16552
rect 6698 16496 8390 16552
rect 8446 16496 8451 16552
rect 6637 16494 8451 16496
rect 6637 16491 6703 16494
rect 8385 16491 8451 16494
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 5441 16146 5507 16149
rect 9673 16146 9739 16149
rect 5441 16144 9739 16146
rect 5441 16088 5446 16144
rect 5502 16088 9678 16144
rect 9734 16088 9739 16144
rect 5441 16086 9739 16088
rect 5441 16083 5507 16086
rect 9673 16083 9739 16086
rect 4705 16010 4771 16013
rect 10593 16010 10659 16013
rect 4705 16008 10659 16010
rect 4705 15952 4710 16008
rect 4766 15952 10598 16008
rect 10654 15952 10659 16008
rect 4705 15950 10659 15952
rect 4705 15947 4771 15950
rect 10593 15947 10659 15950
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 8477 15602 8543 15605
rect 13353 15602 13419 15605
rect 8477 15600 13419 15602
rect 8477 15544 8482 15600
rect 8538 15544 13358 15600
rect 13414 15544 13419 15600
rect 8477 15542 13419 15544
rect 8477 15539 8543 15542
rect 13353 15539 13419 15542
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 5206 15132 5212 15196
rect 5276 15194 5282 15196
rect 5717 15194 5783 15197
rect 5276 15192 5783 15194
rect 5276 15136 5722 15192
rect 5778 15136 5783 15192
rect 5276 15134 5783 15136
rect 5276 15132 5282 15134
rect 5717 15131 5783 15134
rect 7833 15058 7899 15061
rect 12249 15058 12315 15061
rect 7833 15056 12315 15058
rect 7833 15000 7838 15056
rect 7894 15000 12254 15056
rect 12310 15000 12315 15056
rect 7833 14998 12315 15000
rect 7833 14995 7899 14998
rect 12249 14995 12315 14998
rect 0 14922 480 14952
rect 1669 14922 1735 14925
rect 0 14920 1735 14922
rect 0 14864 1674 14920
rect 1730 14864 1735 14920
rect 0 14862 1735 14864
rect 0 14832 480 14862
rect 1669 14859 1735 14862
rect 2405 14922 2471 14925
rect 7097 14922 7163 14925
rect 2405 14920 7163 14922
rect 2405 14864 2410 14920
rect 2466 14864 7102 14920
rect 7158 14864 7163 14920
rect 2405 14862 7163 14864
rect 2405 14859 2471 14862
rect 7097 14859 7163 14862
rect 7741 14786 7807 14789
rect 8385 14786 8451 14789
rect 9673 14786 9739 14789
rect 7741 14784 9739 14786
rect 7741 14728 7746 14784
rect 7802 14728 8390 14784
rect 8446 14728 9678 14784
rect 9734 14728 9739 14784
rect 7741 14726 9739 14728
rect 7741 14723 7807 14726
rect 8385 14723 8451 14726
rect 9673 14723 9739 14726
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 10225 14514 10291 14517
rect 7054 14512 10291 14514
rect 7054 14456 10230 14512
rect 10286 14456 10291 14512
rect 7054 14454 10291 14456
rect 2589 14378 2655 14381
rect 6821 14378 6887 14381
rect 7054 14378 7114 14454
rect 10225 14451 10291 14454
rect 2589 14376 7114 14378
rect 2589 14320 2594 14376
rect 2650 14320 6826 14376
rect 6882 14320 7114 14376
rect 2589 14318 7114 14320
rect 7189 14378 7255 14381
rect 10041 14378 10107 14381
rect 7189 14376 10107 14378
rect 7189 14320 7194 14376
rect 7250 14320 10046 14376
rect 10102 14320 10107 14376
rect 7189 14318 10107 14320
rect 2589 14315 2655 14318
rect 6821 14315 6887 14318
rect 7189 14315 7255 14318
rect 10041 14315 10107 14318
rect 9581 14242 9647 14245
rect 12341 14242 12407 14245
rect 9581 14240 12407 14242
rect 9581 14184 9586 14240
rect 9642 14184 12346 14240
rect 12402 14184 12407 14240
rect 9581 14182 12407 14184
rect 9581 14179 9647 14182
rect 12341 14179 12407 14182
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 1761 13970 1827 13973
rect 1761 13968 6746 13970
rect 1761 13912 1766 13968
rect 1822 13912 6746 13968
rect 1761 13910 6746 13912
rect 1761 13907 1827 13910
rect 6686 13698 6746 13910
rect 8017 13834 8083 13837
rect 11278 13834 11284 13836
rect 8017 13832 11284 13834
rect 8017 13776 8022 13832
rect 8078 13776 11284 13832
rect 8017 13774 11284 13776
rect 8017 13771 8083 13774
rect 11278 13772 11284 13774
rect 11348 13772 11354 13836
rect 9673 13698 9739 13701
rect 6686 13696 9739 13698
rect 6686 13640 9678 13696
rect 9734 13640 9739 13696
rect 6686 13638 9739 13640
rect 9673 13635 9739 13638
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 4521 13426 4587 13429
rect 10777 13426 10843 13429
rect 4521 13424 10843 13426
rect 4521 13368 4526 13424
rect 4582 13368 10782 13424
rect 10838 13368 10843 13424
rect 4521 13366 10843 13368
rect 4521 13363 4587 13366
rect 10777 13363 10843 13366
rect 2589 13290 2655 13293
rect 4429 13290 4495 13293
rect 7833 13290 7899 13293
rect 10225 13290 10291 13293
rect 2589 13288 10291 13290
rect 2589 13232 2594 13288
rect 2650 13232 4434 13288
rect 4490 13232 7838 13288
rect 7894 13232 10230 13288
rect 10286 13232 10291 13288
rect 2589 13230 10291 13232
rect 2589 13227 2655 13230
rect 4429 13227 4495 13230
rect 7833 13227 7899 13230
rect 10225 13227 10291 13230
rect 11145 13154 11211 13157
rect 13077 13154 13143 13157
rect 11145 13152 13143 13154
rect 11145 13096 11150 13152
rect 11206 13096 13082 13152
rect 13138 13096 13143 13152
rect 11145 13094 13143 13096
rect 11145 13091 11211 13094
rect 13077 13091 13143 13094
rect 3610 13088 3930 13089
rect 0 13018 480 13048
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 480 12958
rect 1577 12955 1643 12958
rect 8661 12746 8727 12749
rect 12525 12746 12591 12749
rect 8661 12744 12591 12746
rect 8661 12688 8666 12744
rect 8722 12688 12530 12744
rect 12586 12688 12591 12744
rect 8661 12686 12591 12688
rect 8661 12683 8727 12686
rect 12525 12683 12591 12686
rect 10041 12612 10107 12613
rect 9990 12548 9996 12612
rect 10060 12610 10107 12612
rect 10060 12608 10152 12610
rect 10102 12552 10152 12608
rect 10060 12550 10152 12552
rect 10060 12548 10107 12550
rect 10041 12547 10107 12548
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 4705 12474 4771 12477
rect 9622 12474 9628 12476
rect 4705 12472 6194 12474
rect 4705 12416 4710 12472
rect 4766 12416 6194 12472
rect 4705 12414 6194 12416
rect 4705 12411 4771 12414
rect 1393 12338 1459 12341
rect 2037 12338 2103 12341
rect 5809 12338 5875 12341
rect 1393 12336 5875 12338
rect 1393 12280 1398 12336
rect 1454 12280 2042 12336
rect 2098 12280 5814 12336
rect 5870 12280 5875 12336
rect 1393 12278 5875 12280
rect 6134 12338 6194 12414
rect 6686 12414 9628 12474
rect 6686 12338 6746 12414
rect 9622 12412 9628 12414
rect 9692 12474 9698 12476
rect 10409 12474 10475 12477
rect 10777 12474 10843 12477
rect 9692 12414 10196 12474
rect 9692 12412 9698 12414
rect 10136 12341 10196 12414
rect 10409 12472 10843 12474
rect 10409 12416 10414 12472
rect 10470 12416 10782 12472
rect 10838 12416 10843 12472
rect 10409 12414 10843 12416
rect 10409 12411 10475 12414
rect 10777 12411 10843 12414
rect 6134 12278 6746 12338
rect 9673 12338 9739 12341
rect 9990 12338 9996 12340
rect 9673 12336 9996 12338
rect 9673 12280 9678 12336
rect 9734 12280 9996 12336
rect 9673 12278 9996 12280
rect 1393 12275 1459 12278
rect 2037 12275 2103 12278
rect 5809 12275 5875 12278
rect 9673 12275 9739 12278
rect 9990 12276 9996 12278
rect 10060 12276 10066 12340
rect 10133 12336 10199 12341
rect 10133 12280 10138 12336
rect 10194 12280 10199 12336
rect 10133 12275 10199 12280
rect 11278 12276 11284 12340
rect 11348 12338 11354 12340
rect 11973 12338 12039 12341
rect 11348 12336 12039 12338
rect 11348 12280 11978 12336
rect 12034 12280 12039 12336
rect 11348 12278 12039 12280
rect 11348 12276 11354 12278
rect 11973 12275 12039 12278
rect 10777 12066 10843 12069
rect 11329 12066 11395 12069
rect 10777 12064 11395 12066
rect 10777 12008 10782 12064
rect 10838 12008 11334 12064
rect 11390 12008 11395 12064
rect 10777 12006 11395 12008
rect 10777 12003 10843 12006
rect 11329 12003 11395 12006
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 3601 11794 3667 11797
rect 9489 11794 9555 11797
rect 10317 11794 10383 11797
rect 3601 11792 10383 11794
rect 3601 11736 3606 11792
rect 3662 11736 9494 11792
rect 9550 11736 10322 11792
rect 10378 11736 10383 11792
rect 3601 11734 10383 11736
rect 3601 11731 3667 11734
rect 9489 11731 9555 11734
rect 10317 11731 10383 11734
rect 10501 11796 10567 11797
rect 10501 11792 10548 11796
rect 10612 11794 10618 11796
rect 10501 11736 10506 11792
rect 10501 11732 10548 11736
rect 10612 11734 10658 11794
rect 10612 11732 10618 11734
rect 10501 11731 10567 11732
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3141 11386 3207 11389
rect 5901 11386 5967 11389
rect 3141 11384 5967 11386
rect 3141 11328 3146 11384
rect 3202 11328 5906 11384
rect 5962 11328 5967 11384
rect 3141 11326 5967 11328
rect 3141 11323 3207 11326
rect 5901 11323 5967 11326
rect 3509 11250 3575 11253
rect 5165 11252 5231 11253
rect 5165 11250 5212 11252
rect 3509 11248 5212 11250
rect 3509 11192 3514 11248
rect 3570 11192 5170 11248
rect 3509 11190 5212 11192
rect 3509 11187 3575 11190
rect 5165 11188 5212 11190
rect 5276 11188 5282 11252
rect 5993 11250 6059 11253
rect 12709 11250 12775 11253
rect 5993 11248 12775 11250
rect 5993 11192 5998 11248
rect 6054 11192 12714 11248
rect 12770 11192 12775 11248
rect 5993 11190 12775 11192
rect 5165 11187 5231 11188
rect 5993 11187 6059 11190
rect 12709 11187 12775 11190
rect 0 10978 480 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 480 10918
rect 1577 10915 1643 10918
rect 9397 10978 9463 10981
rect 13445 10978 13511 10981
rect 9397 10976 13511 10978
rect 9397 10920 9402 10976
rect 9458 10920 13450 10976
rect 13506 10920 13511 10976
rect 9397 10918 13511 10920
rect 9397 10915 9463 10918
rect 13445 10915 13511 10918
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 13445 10706 13511 10709
rect 15377 10706 15443 10709
rect 13445 10704 15443 10706
rect 13445 10648 13450 10704
rect 13506 10648 15382 10704
rect 15438 10648 15443 10704
rect 13445 10646 15443 10648
rect 13445 10643 13511 10646
rect 15377 10643 15443 10646
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 4153 10162 4219 10165
rect 8477 10162 8543 10165
rect 4153 10160 8543 10162
rect 4153 10104 4158 10160
rect 4214 10104 8482 10160
rect 8538 10104 8543 10160
rect 4153 10102 8543 10104
rect 4153 10099 4219 10102
rect 8477 10099 8543 10102
rect 12157 10026 12223 10029
rect 15520 10026 16000 10056
rect 12157 10024 16000 10026
rect 12157 9968 12162 10024
rect 12218 9968 16000 10024
rect 12157 9966 16000 9968
rect 12157 9963 12223 9966
rect 15520 9936 16000 9966
rect 9397 9890 9463 9893
rect 11237 9890 11303 9893
rect 9397 9888 11303 9890
rect 9397 9832 9402 9888
rect 9458 9832 11242 9888
rect 11298 9832 11303 9888
rect 9397 9830 11303 9832
rect 9397 9827 9463 9830
rect 11237 9827 11303 9830
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 9397 9754 9463 9757
rect 11053 9754 11119 9757
rect 9397 9752 11119 9754
rect 9397 9696 9402 9752
rect 9458 9696 11058 9752
rect 11114 9696 11119 9752
rect 9397 9694 11119 9696
rect 9397 9691 9463 9694
rect 11053 9691 11119 9694
rect 6453 9618 6519 9621
rect 10041 9618 10107 9621
rect 6453 9616 10107 9618
rect 6453 9560 6458 9616
rect 6514 9560 10046 9616
rect 10102 9560 10107 9616
rect 6453 9558 10107 9560
rect 6453 9555 6519 9558
rect 10041 9555 10107 9558
rect 5901 9346 5967 9349
rect 6085 9346 6151 9349
rect 5901 9344 6151 9346
rect 5901 9288 5906 9344
rect 5962 9288 6090 9344
rect 6146 9288 6151 9344
rect 5901 9286 6151 9288
rect 5901 9283 5967 9286
rect 6085 9283 6151 9286
rect 8201 9346 8267 9349
rect 9857 9346 9923 9349
rect 8201 9344 9923 9346
rect 8201 9288 8206 9344
rect 8262 9288 9862 9344
rect 9918 9288 9923 9344
rect 8201 9286 9923 9288
rect 8201 9283 8267 9286
rect 9857 9283 9923 9286
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 5165 9210 5231 9213
rect 5165 9208 5274 9210
rect 5165 9152 5170 9208
rect 5226 9152 5274 9208
rect 5165 9147 5274 9152
rect 5214 9074 5274 9147
rect 13721 9074 13787 9077
rect 5214 9072 13787 9074
rect 5214 9016 13726 9072
rect 13782 9016 13787 9072
rect 5214 9014 13787 9016
rect 13721 9011 13787 9014
rect 0 8938 480 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 480 8878
rect 1577 8875 1643 8878
rect 12341 8938 12407 8941
rect 15745 8938 15811 8941
rect 12341 8936 15811 8938
rect 12341 8880 12346 8936
rect 12402 8880 15750 8936
rect 15806 8880 15811 8936
rect 12341 8878 15811 8880
rect 12341 8875 12407 8878
rect 15745 8875 15811 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 3049 8394 3115 8397
rect 9673 8394 9739 8397
rect 3049 8392 9739 8394
rect 3049 8336 3054 8392
rect 3110 8336 9678 8392
rect 9734 8336 9739 8392
rect 3049 8334 9739 8336
rect 3049 8331 3115 8334
rect 9673 8331 9739 8334
rect 11973 8396 12039 8397
rect 11973 8392 12020 8396
rect 12084 8394 12090 8396
rect 11973 8336 11978 8392
rect 11973 8332 12020 8336
rect 12084 8334 12130 8394
rect 12084 8332 12090 8334
rect 11973 8331 12039 8332
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 7465 7850 7531 7853
rect 13169 7850 13235 7853
rect 13629 7850 13695 7853
rect 7465 7848 13695 7850
rect 7465 7792 7470 7848
rect 7526 7792 13174 7848
rect 13230 7792 13634 7848
rect 13690 7792 13695 7848
rect 7465 7790 13695 7792
rect 7465 7787 7531 7790
rect 13169 7787 13235 7790
rect 13629 7787 13695 7790
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 4337 7442 4403 7445
rect 8661 7442 8727 7445
rect 9213 7442 9279 7445
rect 4337 7440 9279 7442
rect 4337 7384 4342 7440
rect 4398 7384 8666 7440
rect 8722 7384 9218 7440
rect 9274 7384 9279 7440
rect 4337 7382 9279 7384
rect 4337 7379 4403 7382
rect 8661 7379 8727 7382
rect 9213 7379 9279 7382
rect 3325 7306 3391 7309
rect 10501 7306 10567 7309
rect 3325 7304 10567 7306
rect 3325 7248 3330 7304
rect 3386 7248 10506 7304
rect 10562 7248 10567 7304
rect 3325 7246 10567 7248
rect 3325 7243 3391 7246
rect 10501 7243 10567 7246
rect 10777 7306 10843 7309
rect 12893 7306 12959 7309
rect 10777 7304 12959 7306
rect 10777 7248 10782 7304
rect 10838 7248 12898 7304
rect 12954 7248 12959 7304
rect 10777 7246 12959 7248
rect 10777 7243 10843 7246
rect 12893 7243 12959 7246
rect 2957 7170 3023 7173
rect 5625 7170 5691 7173
rect 2957 7168 5691 7170
rect 2957 7112 2962 7168
rect 3018 7112 5630 7168
rect 5686 7112 5691 7168
rect 2957 7110 5691 7112
rect 2957 7107 3023 7110
rect 5625 7107 5691 7110
rect 8385 7170 8451 7173
rect 9673 7170 9739 7173
rect 8385 7168 9739 7170
rect 8385 7112 8390 7168
rect 8446 7112 9678 7168
rect 9734 7112 9739 7168
rect 8385 7110 9739 7112
rect 8385 7107 8451 7110
rect 6277 7104 6597 7105
rect 0 7034 480 7064
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 9400 7037 9460 7110
rect 9673 7107 9739 7110
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 2313 7034 2379 7037
rect 8293 7034 8359 7037
rect 0 7032 2379 7034
rect 0 6976 2318 7032
rect 2374 6976 2379 7032
rect 0 6974 2379 6976
rect 0 6944 480 6974
rect 2313 6971 2379 6974
rect 7790 7032 8359 7034
rect 7790 6976 8298 7032
rect 8354 6976 8359 7032
rect 7790 6974 8359 6976
rect 2773 6898 2839 6901
rect 5901 6898 5967 6901
rect 7790 6898 7850 6974
rect 8293 6971 8359 6974
rect 9397 7032 9463 7037
rect 11421 7036 11487 7037
rect 11421 7034 11468 7036
rect 9397 6976 9402 7032
rect 9458 6976 9463 7032
rect 9397 6971 9463 6976
rect 11376 7032 11468 7034
rect 11376 6976 11426 7032
rect 11376 6974 11468 6976
rect 11421 6972 11468 6974
rect 11532 6972 11538 7036
rect 11421 6971 11487 6972
rect 2773 6896 7850 6898
rect 2773 6840 2778 6896
rect 2834 6840 5906 6896
rect 5962 6840 7850 6896
rect 2773 6838 7850 6840
rect 2773 6835 2839 6838
rect 5901 6835 5967 6838
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 3601 6354 3667 6357
rect 7005 6354 7071 6357
rect 3601 6352 7071 6354
rect 3601 6296 3606 6352
rect 3662 6296 7010 6352
rect 7066 6296 7071 6352
rect 3601 6294 7071 6296
rect 3601 6291 3667 6294
rect 7005 6291 7071 6294
rect 4705 6218 4771 6221
rect 7741 6218 7807 6221
rect 4705 6216 7807 6218
rect 4705 6160 4710 6216
rect 4766 6160 7746 6216
rect 7802 6160 7807 6216
rect 4705 6158 7807 6160
rect 4705 6155 4771 6158
rect 7741 6155 7807 6158
rect 2497 6082 2563 6085
rect 6085 6082 6151 6085
rect 2497 6080 6151 6082
rect 2497 6024 2502 6080
rect 2558 6024 6090 6080
rect 6146 6024 6151 6080
rect 2497 6022 6151 6024
rect 2497 6019 2563 6022
rect 6085 6019 6151 6022
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 7005 5946 7071 5949
rect 7557 5946 7623 5949
rect 10685 5946 10751 5949
rect 7005 5944 10751 5946
rect 7005 5888 7010 5944
rect 7066 5888 7562 5944
rect 7618 5888 10690 5944
rect 10746 5888 10751 5944
rect 7005 5886 10751 5888
rect 7005 5883 7071 5886
rect 7557 5883 7623 5886
rect 10685 5883 10751 5886
rect 9397 5810 9463 5813
rect 10409 5810 10475 5813
rect 12525 5810 12591 5813
rect 9397 5808 12591 5810
rect 9397 5752 9402 5808
rect 9458 5752 10414 5808
rect 10470 5752 12530 5808
rect 12586 5752 12591 5808
rect 9397 5750 12591 5752
rect 9397 5747 9463 5750
rect 10409 5747 10475 5750
rect 12525 5747 12591 5750
rect 565 5674 631 5677
rect 4245 5674 4311 5677
rect 565 5672 4311 5674
rect 565 5616 570 5672
rect 626 5616 4250 5672
rect 4306 5616 4311 5672
rect 565 5614 4311 5616
rect 565 5611 631 5614
rect 4245 5611 4311 5614
rect 5257 5674 5323 5677
rect 7189 5674 7255 5677
rect 5257 5672 7255 5674
rect 5257 5616 5262 5672
rect 5318 5616 7194 5672
rect 7250 5616 7255 5672
rect 5257 5614 7255 5616
rect 5257 5611 5323 5614
rect 7189 5611 7255 5614
rect 7925 5674 7991 5677
rect 12433 5674 12499 5677
rect 7925 5672 12499 5674
rect 7925 5616 7930 5672
rect 7986 5616 12438 5672
rect 12494 5616 12499 5672
rect 7925 5614 12499 5616
rect 7925 5611 7991 5614
rect 12433 5611 12499 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 7373 5266 7439 5269
rect 10777 5266 10843 5269
rect 7373 5264 10843 5266
rect 7373 5208 7378 5264
rect 7434 5208 10782 5264
rect 10838 5208 10843 5264
rect 7373 5206 10843 5208
rect 7373 5203 7439 5206
rect 10777 5203 10843 5206
rect 5717 5130 5783 5133
rect 5901 5130 5967 5133
rect 10409 5130 10475 5133
rect 5717 5128 10475 5130
rect 5717 5072 5722 5128
rect 5778 5072 5906 5128
rect 5962 5072 10414 5128
rect 10470 5072 10475 5128
rect 5717 5070 10475 5072
rect 5717 5067 5783 5070
rect 5901 5067 5967 5070
rect 10409 5067 10475 5070
rect 0 4994 480 5024
rect 1577 4994 1643 4997
rect 0 4992 1643 4994
rect 0 4936 1582 4992
rect 1638 4936 1643 4992
rect 0 4934 1643 4936
rect 0 4904 480 4934
rect 1577 4931 1643 4934
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 6085 4722 6151 4725
rect 9857 4722 9923 4725
rect 6085 4720 9923 4722
rect 6085 4664 6090 4720
rect 6146 4664 9862 4720
rect 9918 4664 9923 4720
rect 6085 4662 9923 4664
rect 6085 4659 6151 4662
rect 9857 4659 9923 4662
rect 2865 4586 2931 4589
rect 7465 4586 7531 4589
rect 10225 4586 10291 4589
rect 2865 4584 7531 4586
rect 2865 4528 2870 4584
rect 2926 4528 7470 4584
rect 7526 4528 7531 4584
rect 2865 4526 7531 4528
rect 2865 4523 2931 4526
rect 7465 4523 7531 4526
rect 7606 4584 10291 4586
rect 7606 4528 10230 4584
rect 10286 4528 10291 4584
rect 7606 4526 10291 4528
rect 5349 4450 5415 4453
rect 7281 4450 7347 4453
rect 5349 4448 7347 4450
rect 5349 4392 5354 4448
rect 5410 4392 7286 4448
rect 7342 4392 7347 4448
rect 5349 4390 7347 4392
rect 5349 4387 5415 4390
rect 7281 4387 7347 4390
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 5625 4314 5691 4317
rect 7606 4314 7666 4526
rect 10225 4523 10291 4526
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 5625 4312 7666 4314
rect 5625 4256 5630 4312
rect 5686 4256 7666 4312
rect 5625 4254 7666 4256
rect 11881 4314 11947 4317
rect 12014 4314 12020 4316
rect 11881 4312 12020 4314
rect 11881 4256 11886 4312
rect 11942 4256 12020 4312
rect 11881 4254 12020 4256
rect 5625 4251 5691 4254
rect 11881 4251 11947 4254
rect 12014 4252 12020 4254
rect 12084 4252 12090 4316
rect 197 4178 263 4181
rect 3141 4178 3207 4181
rect 197 4176 3207 4178
rect 197 4120 202 4176
rect 258 4120 3146 4176
rect 3202 4120 3207 4176
rect 197 4118 3207 4120
rect 197 4115 263 4118
rect 3141 4115 3207 4118
rect 3325 4178 3391 4181
rect 6361 4178 6427 4181
rect 3325 4176 6427 4178
rect 3325 4120 3330 4176
rect 3386 4120 6366 4176
rect 6422 4120 6427 4176
rect 3325 4118 6427 4120
rect 3325 4115 3391 4118
rect 6361 4115 6427 4118
rect 7741 4178 7807 4181
rect 13537 4178 13603 4181
rect 7741 4176 13603 4178
rect 7741 4120 7746 4176
rect 7802 4120 13542 4176
rect 13598 4120 13603 4176
rect 7741 4118 13603 4120
rect 7741 4115 7807 4118
rect 13537 4115 13603 4118
rect 6269 4042 6335 4045
rect 8017 4042 8083 4045
rect 11513 4042 11579 4045
rect 6269 4040 7298 4042
rect 6269 3984 6274 4040
rect 6330 3984 7298 4040
rect 6269 3982 7298 3984
rect 6269 3979 6335 3982
rect 7238 3906 7298 3982
rect 8017 4040 11579 4042
rect 8017 3984 8022 4040
rect 8078 3984 11518 4040
rect 11574 3984 11579 4040
rect 8017 3982 11579 3984
rect 8017 3979 8083 3982
rect 11513 3979 11579 3982
rect 13721 4042 13787 4045
rect 14641 4042 14707 4045
rect 13721 4040 14707 4042
rect 13721 3984 13726 4040
rect 13782 3984 14646 4040
rect 14702 3984 14707 4040
rect 13721 3982 14707 3984
rect 13721 3979 13787 3982
rect 14641 3979 14707 3982
rect 10317 3906 10383 3909
rect 7238 3904 10383 3906
rect 7238 3848 10322 3904
rect 10378 3848 10383 3904
rect 7238 3846 10383 3848
rect 10317 3843 10383 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 1761 3770 1827 3773
rect 5717 3770 5783 3773
rect 1761 3768 5783 3770
rect 1761 3712 1766 3768
rect 1822 3712 5722 3768
rect 5778 3712 5783 3768
rect 1761 3710 5783 3712
rect 1761 3707 1827 3710
rect 5717 3707 5783 3710
rect 1669 3634 1735 3637
rect 9305 3634 9371 3637
rect 1669 3632 9371 3634
rect 1669 3576 1674 3632
rect 1730 3576 9310 3632
rect 9366 3576 9371 3632
rect 1669 3574 9371 3576
rect 1669 3571 1735 3574
rect 9305 3571 9371 3574
rect 4521 3498 4587 3501
rect 11053 3498 11119 3501
rect 4521 3496 11119 3498
rect 4521 3440 4526 3496
rect 4582 3440 11058 3496
rect 11114 3440 11119 3496
rect 4521 3438 11119 3440
rect 4521 3435 4587 3438
rect 11053 3435 11119 3438
rect 12249 3498 12315 3501
rect 12249 3496 14842 3498
rect 12249 3440 12254 3496
rect 12310 3440 14842 3496
rect 12249 3438 14842 3440
rect 12249 3435 12315 3438
rect 4705 3362 4771 3365
rect 8477 3362 8543 3365
rect 4705 3360 8543 3362
rect 4705 3304 4710 3360
rect 4766 3304 8482 3360
rect 8538 3304 8543 3360
rect 4705 3302 8543 3304
rect 14782 3362 14842 3438
rect 15520 3362 16000 3392
rect 14782 3302 16000 3362
rect 4705 3299 4771 3302
rect 8477 3299 8543 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 15520 3272 16000 3302
rect 14277 3231 14597 3232
rect 4245 3226 4311 3229
rect 11605 3226 11671 3229
rect 13813 3226 13879 3229
rect 4245 3224 8540 3226
rect 4245 3168 4250 3224
rect 4306 3168 8540 3224
rect 4245 3166 8540 3168
rect 4245 3163 4311 3166
rect 3969 3090 4035 3093
rect 8293 3090 8359 3093
rect 3969 3088 8359 3090
rect 3969 3032 3974 3088
rect 4030 3032 8298 3088
rect 8354 3032 8359 3088
rect 3969 3030 8359 3032
rect 8480 3090 8540 3166
rect 11286 3224 13879 3226
rect 11286 3168 11610 3224
rect 11666 3168 13818 3224
rect 13874 3168 13879 3224
rect 11286 3166 13879 3168
rect 11053 3090 11119 3093
rect 8480 3088 11119 3090
rect 8480 3032 11058 3088
rect 11114 3032 11119 3088
rect 8480 3030 11119 3032
rect 3969 3027 4035 3030
rect 8293 3027 8359 3030
rect 11053 3027 11119 3030
rect 0 2954 480 2984
rect 1945 2954 2011 2957
rect 0 2952 2011 2954
rect 0 2896 1950 2952
rect 2006 2896 2011 2952
rect 0 2894 2011 2896
rect 0 2864 480 2894
rect 1945 2891 2011 2894
rect 3509 2954 3575 2957
rect 9121 2954 9187 2957
rect 3509 2952 9187 2954
rect 3509 2896 3514 2952
rect 3570 2896 9126 2952
rect 9182 2896 9187 2952
rect 3509 2894 9187 2896
rect 3509 2891 3575 2894
rect 9121 2891 9187 2894
rect 9673 2954 9739 2957
rect 10041 2954 10107 2957
rect 11286 2954 11346 3166
rect 11605 3163 11671 3166
rect 13813 3163 13879 3166
rect 9673 2952 11346 2954
rect 9673 2896 9678 2952
rect 9734 2896 10046 2952
rect 10102 2896 11346 2952
rect 9673 2894 11346 2896
rect 9673 2891 9739 2894
rect 10041 2891 10107 2894
rect 2681 2818 2747 2821
rect 4337 2818 4403 2821
rect 2681 2816 4403 2818
rect 2681 2760 2686 2816
rect 2742 2760 4342 2816
rect 4398 2760 4403 2816
rect 2681 2758 4403 2760
rect 2681 2755 2747 2758
rect 4337 2755 4403 2758
rect 7649 2818 7715 2821
rect 7925 2818 7991 2821
rect 7649 2816 7991 2818
rect 7649 2760 7654 2816
rect 7710 2760 7930 2816
rect 7986 2760 7991 2816
rect 7649 2758 7991 2760
rect 7649 2755 7715 2758
rect 7925 2755 7991 2758
rect 8477 2818 8543 2821
rect 8845 2818 8911 2821
rect 9489 2818 9555 2821
rect 10409 2818 10475 2821
rect 8477 2816 10475 2818
rect 8477 2760 8482 2816
rect 8538 2760 8850 2816
rect 8906 2760 9494 2816
rect 9550 2760 10414 2816
rect 10470 2760 10475 2816
rect 8477 2758 10475 2760
rect 8477 2755 8543 2758
rect 8845 2755 8911 2758
rect 9489 2755 9555 2758
rect 10409 2755 10475 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 2405 2682 2471 2685
rect 5073 2682 5139 2685
rect 2405 2680 5139 2682
rect 2405 2624 2410 2680
rect 2466 2624 5078 2680
rect 5134 2624 5139 2680
rect 2405 2622 5139 2624
rect 2405 2619 2471 2622
rect 5073 2619 5139 2622
rect 11462 2484 11468 2548
rect 11532 2546 11538 2548
rect 11789 2546 11855 2549
rect 11532 2544 11855 2546
rect 11532 2488 11794 2544
rect 11850 2488 11855 2544
rect 11532 2486 11855 2488
rect 11532 2484 11538 2486
rect 11789 2483 11855 2486
rect 8477 2410 8543 2413
rect 14917 2410 14983 2413
rect 8477 2408 14983 2410
rect 8477 2352 8482 2408
rect 8538 2352 14922 2408
rect 14978 2352 14983 2408
rect 8477 2350 14983 2352
rect 8477 2347 8543 2350
rect 14917 2347 14983 2350
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 5257 2002 5323 2005
rect 13721 2002 13787 2005
rect 5257 2000 13787 2002
rect 5257 1944 5262 2000
rect 5318 1944 13726 2000
rect 13782 1944 13787 2000
rect 5257 1942 13787 1944
rect 5257 1939 5323 1942
rect 13721 1939 13787 1942
rect 2589 1458 2655 1461
rect 7097 1458 7163 1461
rect 2589 1456 7163 1458
rect 2589 1400 2594 1456
rect 2650 1400 7102 1456
rect 7158 1400 7163 1456
rect 2589 1398 7163 1400
rect 2589 1395 2655 1398
rect 7097 1395 7163 1398
rect 0 1050 480 1080
rect 2497 1050 2563 1053
rect 0 1048 2563 1050
rect 0 992 2502 1048
rect 2558 992 2563 1048
rect 0 990 2563 992
rect 0 960 480 990
rect 2497 987 2563 990
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 8156 34308 8220 34372
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 9996 32056 10060 32060
rect 9996 32000 10046 32056
rect 10046 32000 10060 32056
rect 9996 31996 10060 32000
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 8156 29820 8220 29884
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 9996 29004 10060 29068
rect 9996 28868 10060 28932
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 6132 28596 6196 28660
rect 9444 28460 9508 28524
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 9444 24652 9508 24716
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 9996 20224 10060 20228
rect 9996 20168 10010 20224
rect 10010 20168 10060 20224
rect 9996 20164 10060 20168
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 6132 19892 6196 19956
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 9628 18940 9692 19004
rect 10548 18532 10612 18596
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 10548 17988 10612 18052
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 5212 15132 5276 15196
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 11284 13772 11348 13836
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 9996 12608 10060 12612
rect 9996 12552 10046 12608
rect 10046 12552 10060 12608
rect 9996 12548 10060 12552
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 9628 12412 9692 12476
rect 9996 12276 10060 12340
rect 11284 12276 11348 12340
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 10548 11792 10612 11796
rect 10548 11736 10562 11792
rect 10562 11736 10612 11792
rect 10548 11732 10612 11736
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 5212 11248 5276 11252
rect 5212 11192 5226 11248
rect 5226 11192 5276 11248
rect 5212 11188 5276 11192
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 12020 8392 12084 8396
rect 12020 8336 12034 8392
rect 12034 8336 12084 8392
rect 12020 8332 12084 8336
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 11468 7032 11532 7036
rect 11468 6976 11482 7032
rect 11482 6976 11532 7032
rect 11468 6972 11532 6976
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 12020 4252 12084 4316
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 11468 2484 11532 2548
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8155 34372 8221 34373
rect 8155 34308 8156 34372
rect 8220 34308 8221 34372
rect 8155 34307 8221 34308
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 8158 29885 8218 34307
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 9995 32060 10061 32061
rect 9995 31996 9996 32060
rect 10060 31996 10061 32060
rect 9995 31995 10061 31996
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8155 29884 8221 29885
rect 8155 29820 8156 29884
rect 8220 29820 8221 29884
rect 8155 29819 8221 29820
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6131 28660 6197 28661
rect 6131 28596 6132 28660
rect 6196 28596 6197 28660
rect 6131 28595 6197 28596
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 6134 19957 6194 28595
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6131 19956 6197 19957
rect 6131 19892 6132 19956
rect 6196 19892 6197 19956
rect 6131 19891 6197 19892
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 5211 15196 5277 15197
rect 5211 15132 5212 15196
rect 5276 15132 5277 15196
rect 5211 15131 5277 15132
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 5214 11253 5274 15131
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 5211 11252 5277 11253
rect 5211 11188 5212 11252
rect 5276 11188 5277 11252
rect 5211 11187 5277 11188
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 9998 29069 10058 31995
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 9995 29068 10061 29069
rect 9995 29004 9996 29068
rect 10060 29004 10061 29068
rect 9995 29003 10061 29004
rect 9995 28932 10061 28933
rect 9995 28868 9996 28932
rect 10060 28868 10061 28932
rect 9995 28867 10061 28868
rect 9443 28524 9509 28525
rect 9443 28460 9444 28524
rect 9508 28460 9509 28524
rect 9443 28459 9509 28460
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 9446 24717 9506 28459
rect 9443 24716 9509 24717
rect 9443 24652 9444 24716
rect 9508 24652 9509 24716
rect 9443 24651 9509 24652
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 9998 20229 10058 28867
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 9995 20228 10061 20229
rect 9995 20164 9996 20228
rect 10060 20164 10061 20228
rect 9995 20163 10061 20164
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 9627 19004 9693 19005
rect 9627 18940 9628 19004
rect 9692 18940 9693 19004
rect 9627 18939 9693 18940
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 9630 12477 9690 18939
rect 10547 18596 10613 18597
rect 10547 18532 10548 18596
rect 10612 18532 10613 18596
rect 10547 18531 10613 18532
rect 10550 18053 10610 18531
rect 10547 18052 10613 18053
rect 10547 17988 10548 18052
rect 10612 17988 10613 18052
rect 10547 17987 10613 17988
rect 9995 12612 10061 12613
rect 9995 12548 9996 12612
rect 10060 12548 10061 12612
rect 9995 12547 10061 12548
rect 9627 12476 9693 12477
rect 9627 12412 9628 12476
rect 9692 12412 9693 12476
rect 9627 12411 9693 12412
rect 9998 12341 10058 12547
rect 9995 12340 10061 12341
rect 9995 12276 9996 12340
rect 10060 12276 10061 12340
rect 9995 12275 10061 12276
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 10550 11797 10610 17987
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11283 13836 11349 13837
rect 11283 13772 11284 13836
rect 11348 13772 11349 13836
rect 11283 13771 11349 13772
rect 11286 12341 11346 13771
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11283 12340 11349 12341
rect 11283 12276 11284 12340
rect 11348 12276 11349 12340
rect 11283 12275 11349 12276
rect 10547 11796 10613 11797
rect 10547 11732 10548 11796
rect 10612 11732 10613 11796
rect 10547 11731 10613 11732
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 12019 8396 12085 8397
rect 12019 8332 12020 8396
rect 12084 8332 12085 8396
rect 12019 8331 12085 8332
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11467 7036 11533 7037
rect 11467 6972 11468 7036
rect 11532 6972 11533 7036
rect 11467 6971 11533 6972
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 11470 2549 11530 6971
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 12022 4317 12082 8331
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 12019 4316 12085 4317
rect 12019 4252 12020 4316
rect 12084 4252 12085 4316
rect 12019 4251 12085 4252
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11467 2548 11533 2549
rect 11467 2484 11468 2548
rect 11532 2484 11533 2548
rect 11467 2483 11533 2484
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 2128 11930 2688
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_34 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4232 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37
timestamp 1604681595
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4876 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_50
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50
timestamp 1604681595
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_54
timestamp 1604681595
transform 1 0 6072 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58
timestamp 1604681595
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1604681595
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10028 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_140 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13984 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_142
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_6
timestamp 1604681595
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1604681595
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_38
timestamp 1604681595
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 8096 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1604681595
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10028 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1604681595
transform 1 0 8924 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1604681595
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11592 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_110
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_133 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_13
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_16
timestamp 1604681595
transform 1 0 2576 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_3_40
timestamp 1604681595
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_52
timestamp 1604681595
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 5520 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_56
timestamp 1604681595
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_85
timestamp 1604681595
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_136 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4968 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_4_61
timestamp 1604681595
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_65
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_78
timestamp 1604681595
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1604681595
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10212 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_86
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1604681595
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1604681595
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11776 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 13340 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_137
timestamp 1604681595
transform 1 0 13708 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1604681595
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3404 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1604681595
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1604681595
transform 1 0 5520 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_55
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_108
timestamp 1604681595
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_116
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_136
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1604681595
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 1840 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp 1604681595
transform 1 0 2576 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_12
timestamp 1604681595
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 2944 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 2300 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_17
timestamp 1604681595
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_28
timestamp 1604681595
transform 1 0 3680 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1604681595
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_34
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_41
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_46
timestamp 1604681595
transform 1 0 5336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 5612 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp 1604681595
transform 1 0 7728 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_68
timestamp 1604681595
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_71
timestamp 1604681595
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_64
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 6992 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_77
timestamp 1604681595
transform 1 0 8188 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_99
timestamp 1604681595
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_95
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1604681595
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_132
timestamp 1604681595
transform 1 0 13248 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_126
timestamp 1604681595
transform 1 0 12696 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_138
timestamp 1604681595
transform 1 0 13800 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 2024 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_14
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_18
timestamp 1604681595
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1604681595
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_48
timestamp 1604681595
transform 1 0 5520 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1604681595
transform 1 0 6992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1604681595
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_108
timestamp 1604681595
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_131
timestamp 1604681595
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_17
timestamp 1604681595
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_25
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_30
timestamp 1604681595
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_42
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_46
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_58
timestamp 1604681595
transform 1 0 6440 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_70
timestamp 1604681595
transform 1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1604681595
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_140
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1604681595
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 1604681595
transform 1 0 5612 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_53
timestamp 1604681595
transform 1 0 5980 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_60
timestamp 1604681595
transform 1 0 6624 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11684 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_106
timestamp 1604681595
transform 1 0 10856 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_112
timestamp 1604681595
transform 1 0 11408 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_134
timestamp 1604681595
transform 1 0 13432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_103
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_115
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 1472 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_38
timestamp 1604681595
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_42
timestamp 1604681595
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_69
timestamp 1604681595
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_82
timestamp 1604681595
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2852 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1604681595
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_49
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_49
timestamp 1604681595
transform 1 0 5612 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 5336 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6072 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_69
timestamp 1604681595
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_80
timestamp 1604681595
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_76
timestamp 1604681595
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_87
timestamp 1604681595
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 8832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1604681595
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_102
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_111
timestamp 1604681595
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_108
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11500 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1604681595
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_122
timestamp 1604681595
transform 1 0 12328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_134
timestamp 1604681595
transform 1 0 13432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_13
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4508 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_29
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_33
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1604681595
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_50
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_56
timestamp 1604681595
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1604681595
transform 1 0 7084 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_92
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1604681595
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1604681595
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_112
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_126
timestamp 1604681595
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_130
timestamp 1604681595
transform 1 0 13064 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_142
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_24
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1604681595
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_39
timestamp 1604681595
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5428 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_66
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_78
timestamp 1604681595
transform 1 0 8280 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12144 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1604681595
transform 1 0 11776 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_133
timestamp 1604681595
transform 1 0 13340 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_13
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_17
timestamp 1604681595
transform 1 0 2668 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 3128 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_48
timestamp 1604681595
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_52
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_58
timestamp 1604681595
transform 1 0 6440 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_73
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1604681595
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_81
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 11132 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_116
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_136
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_9
timestamp 1604681595
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_13
timestamp 1604681595
transform 1 0 2300 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1604681595
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_24
timestamp 1604681595
transform 1 0 3312 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1604681595
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_63
timestamp 1604681595
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_67
timestamp 1604681595
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1604681595
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11592 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_133
timestamp 1604681595
transform 1 0 13340 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1604681595
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_8
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_13
timestamp 1604681595
transform 1 0 2300 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2208 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1604681595
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_35
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_31
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_51
timestamp 1604681595
transform 1 0 5796 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1604681595
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_59
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_55
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_70
timestamp 1604681595
transform 1 0 7544 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_79
timestamp 1604681595
transform 1 0 8372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1604681595
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_109
timestamp 1604681595
transform 1 0 11132 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_111
timestamp 1604681595
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1604681595
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1604681595
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11684 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_139
timestamp 1604681595
transform 1 0 13892 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_134
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2116 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1604681595
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1604681595
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6900 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1604681595
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1604681595
transform 1 0 13156 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_134
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_13
timestamp 1604681595
transform 1 0 2300 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5612 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_62
timestamp 1604681595
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7176 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_65
timestamp 1604681595
transform 1 0 7084 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_86
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_96
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_100
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_103
timestamp 1604681595
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1604681595
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1604681595
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 1604681595
transform 1 0 13156 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_138
timestamp 1604681595
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_9
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_13
timestamp 1604681595
transform 1 0 2300 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_16
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_40
timestamp 1604681595
transform 1 0 4784 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 1604681595
transform 1 0 5520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_70
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1604681595
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_116
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_143
timestamp 1604681595
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_46
timestamp 1604681595
transform 1 0 5336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_58
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_70
timestamp 1604681595
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_74
timestamp 1604681595
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10028 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11592 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_133
timestamp 1604681595
transform 1 0 13340 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1604681595
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_20
timestamp 1604681595
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_24
timestamp 1604681595
transform 1 0 3312 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_32
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_35
timestamp 1604681595
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp 1604681595
transform 1 0 5060 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7728 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_91
timestamp 1604681595
transform 1 0 9476 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1604681595
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_139
timestamp 1604681595
transform 1 0 13892 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_145
timestamp 1604681595
transform 1 0 14444 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_13
timestamp 1604681595
transform 1 0 2300 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1604681595
transform 1 0 2116 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_21
timestamp 1604681595
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 3404 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1604681595
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_34
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4140 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_46
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_42
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5704 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1604681595
transform 1 0 7452 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1604681595
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_69
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_78
timestamp 1604681595
transform 1 0 8280 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_74
timestamp 1604681595
transform 1 0 7912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8096 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8096 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_95
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_114
timestamp 1604681595
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_110
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11408 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11960 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_137
timestamp 1604681595
transform 1 0 13708 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1604681595
transform 1 0 13616 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4140 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_52
timestamp 1604681595
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_81
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1604681595
transform 1 0 8924 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_106
timestamp 1604681595
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_123
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1604681595
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_131
timestamp 1604681595
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_143
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_34
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8648 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7084 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1604681595
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_99
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_140
timestamp 1604681595
transform 1 0 13984 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_9
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_17
timestamp 1604681595
transform 1 0 2668 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5796 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_46
timestamp 1604681595
transform 1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_50
timestamp 1604681595
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_60
timestamp 1604681595
transform 1 0 6624 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11500 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_110
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_132
timestamp 1604681595
transform 1 0 13248 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_144
timestamp 1604681595
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_35
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_50
timestamp 1604681595
transform 1 0 5704 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1604681595
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1604681595
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7544 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10304 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_99
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1604681595
transform 1 0 11500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1604681595
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_18
timestamp 1604681595
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604681595
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_39
timestamp 1604681595
transform 1 0 4692 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5888 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_43
timestamp 1604681595
transform 1 0 5060 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_51
timestamp 1604681595
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_61
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1604681595
transform 1 0 7084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_77
timestamp 1604681595
transform 1 0 8188 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_81
timestamp 1604681595
transform 1 0 8556 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 10488 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1604681595
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_132
timestamp 1604681595
transform 1 0 13248 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1604681595
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_13
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_17
timestamp 1604681595
transform 1 0 2668 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_25
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_21
timestamp 1604681595
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_29
timestamp 1604681595
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_25
timestamp 1604681595
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_21
timestamp 1604681595
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_33
timestamp 1604681595
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4508 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_41
timestamp 1604681595
transform 1 0 4876 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_49
timestamp 1604681595
transform 1 0 5612 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_50
timestamp 1604681595
transform 1 0 5704 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_46
timestamp 1604681595
transform 1 0 5336 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5796 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 8280 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_70
timestamp 1604681595
transform 1 0 7544 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_75
timestamp 1604681595
transform 1 0 8004 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_81
timestamp 1604681595
transform 1 0 8556 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10212 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604681595
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_116
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_118
timestamp 1604681595
transform 1 0 11960 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_143
timestamp 1604681595
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_130
timestamp 1604681595
transform 1 0 13064 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_142
timestamp 1604681595
transform 1 0 14168 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2392 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1604681595
transform 1 0 1748 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_10
timestamp 1604681595
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_23
timestamp 1604681595
transform 1 0 3220 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_40
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5336 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 5520 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1604681595
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7820 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 7268 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_66
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1604681595
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_82
timestamp 1604681595
transform 1 0 8648 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_90
timestamp 1604681595
transform 1 0 9384 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_95
timestamp 1604681595
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_99
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_103
timestamp 1604681595
transform 1 0 10580 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12052 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1604681595
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1604681595
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_127
timestamp 1604681595
transform 1 0 12788 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_133
timestamp 1604681595
transform 1 0 13340 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_138
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1604681595
transform 1 0 14168 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_51
timestamp 1604681595
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_55
timestamp 1604681595
transform 1 0 6164 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7084 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_36_63
timestamp 1604681595
transform 1 0 6900 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9292 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1604681595
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_102
timestamp 1604681595
transform 1 0 10488 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12052 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_36_114
timestamp 1604681595
transform 1 0 11592 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_118
timestamp 1604681595
transform 1 0 11960 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_138
timestamp 1604681595
transform 1 0 13800 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_11
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_34
timestamp 1604681595
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_38
timestamp 1604681595
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_42
timestamp 1604681595
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7544 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7360 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_66
timestamp 1604681595
transform 1 0 7176 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_79
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9292 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_104
timestamp 1604681595
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_108
timestamp 1604681595
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_112
timestamp 1604681595
transform 1 0 11408 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1604681595
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 12052 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_139
timestamp 1604681595
transform 1 0 13892 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_145
timestamp 1604681595
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_17
timestamp 1604681595
transform 1 0 2668 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4784 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5796 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_49
timestamp 1604681595
transform 1 0 5612 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1604681595
transform 1 0 5980 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_69
timestamp 1604681595
transform 1 0 7452 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_72
timestamp 1604681595
transform 1 0 7728 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9292 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1604681595
transform 1 0 8924 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1604681595
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_99
timestamp 1604681595
transform 1 0 10212 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12052 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_111
timestamp 1604681595
transform 1 0 11316 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_116
timestamp 1604681595
transform 1 0 11776 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_138
timestamp 1604681595
transform 1 0 13800 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_46
timestamp 1604681595
transform 1 0 5336 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_47
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5612 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_55
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5612 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_80
timestamp 1604681595
transform 1 0 8464 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_72
timestamp 1604681595
transform 1 0 7728 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_102
timestamp 1604681595
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_89
timestamp 1604681595
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1604681595
transform 1 0 11224 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_106
timestamp 1604681595
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_106
timestamp 1604681595
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11408 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_116
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11592 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_132
timestamp 1604681595
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_136
timestamp 1604681595
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_140
timestamp 1604681595
transform 1 0 13984 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_133
timestamp 1604681595
transform 1 0 13340 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_30
timestamp 1604681595
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_34
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_40
timestamp 1604681595
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_71
timestamp 1604681595
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_75
timestamp 1604681595
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_79
timestamp 1604681595
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_83
timestamp 1604681595
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_96
timestamp 1604681595
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_100
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1604681595
transform 1 0 11500 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_136
timestamp 1604681595
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_140
timestamp 1604681595
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_144
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 6532 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5980 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_51
timestamp 1604681595
transform 1 0 5796 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_55
timestamp 1604681595
transform 1 0 6164 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_62
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_42_82
timestamp 1604681595
transform 1 0 8648 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10396 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10212 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_86
timestamp 1604681595
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_89
timestamp 1604681595
transform 1 0 9292 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_97
timestamp 1604681595
transform 1 0 10028 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12328 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_110
timestamp 1604681595
transform 1 0 11224 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_114
timestamp 1604681595
transform 1 0 11592 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_131
timestamp 1604681595
transform 1 0 13156 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_143
timestamp 1604681595
transform 1 0 14260 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604681595
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_9
timestamp 1604681595
transform 1 0 1932 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_13
timestamp 1604681595
transform 1 0 2300 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3864 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3496 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_25
timestamp 1604681595
transform 1 0 3404 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_28
timestamp 1604681595
transform 1 0 3680 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1604681595
transform 1 0 5796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1604681595
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8740 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_71
timestamp 1604681595
transform 1 0 7636 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_77
timestamp 1604681595
transform 1 0 8188 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_81
timestamp 1604681595
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 10304 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10120 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9752 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_92
timestamp 1604681595
transform 1 0 9568 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_96
timestamp 1604681595
transform 1 0 9936 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 12512 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11960 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_112
timestamp 1604681595
transform 1 0 11408 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_116
timestamp 1604681595
transform 1 0 11776 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_120
timestamp 1604681595
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_123
timestamp 1604681595
transform 1 0 12420 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1604681595
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_139
timestamp 1604681595
transform 1 0 13892 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_145
timestamp 1604681595
transform 1 0 14444 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604681595
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604681595
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604681595
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1604681595
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604681595
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_32
timestamp 1604681595
transform 1 0 4048 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_36
timestamp 1604681595
transform 1 0 4416 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_40
timestamp 1604681595
transform 1 0 4784 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5244 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7176 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 7544 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_64
timestamp 1604681595
transform 1 0 6992 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_68
timestamp 1604681595
transform 1 0 7360 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_72
timestamp 1604681595
transform 1 0 7728 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_93
timestamp 1604681595
transform 1 0 9660 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_88
timestamp 1604681595
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_84
timestamp 1604681595
transform 1 0 8832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_101
timestamp 1604681595
transform 1 0 10396 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_97
timestamp 1604681595
transform 1 0 10028 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10488 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11500 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_111
timestamp 1604681595
transform 1 0 11316 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_115
timestamp 1604681595
transform 1 0 11684 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_119
timestamp 1604681595
transform 1 0 12052 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_131
timestamp 1604681595
transform 1 0 13156 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_143
timestamp 1604681595
transform 1 0 14260 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604681595
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604681595
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1604681595
transform 1 0 1380 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1604681595
transform 1 0 1748 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_19
timestamp 1604681595
transform 1 0 2852 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3956 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_23
timestamp 1604681595
transform 1 0 3220 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_27
timestamp 1604681595
transform 1 0 3588 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_40
timestamp 1604681595
transform 1 0 4784 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_44
timestamp 1604681595
transform 1 0 5152 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 5520 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 5704 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1604681595
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_53
timestamp 1604681595
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8740 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8372 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_71
timestamp 1604681595
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_75
timestamp 1604681595
transform 1 0 8004 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_81
timestamp 1604681595
transform 1 0 8556 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8924 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_94
timestamp 1604681595
transform 1 0 9752 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_98
timestamp 1604681595
transform 1 0 10120 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11684 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 12052 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_111
timestamp 1604681595
transform 1 0 11316 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_117
timestamp 1604681595
transform 1 0 11868 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_121
timestamp 1604681595
transform 1 0 12236 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1604681595
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1604681595
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_143
timestamp 1604681595
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604681595
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_7
timestamp 1604681595
transform 1 0 1748 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 1932 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604681595
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604681595
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_11
timestamp 1604681595
transform 1 0 2116 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 2300 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1604681595
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_9
timestamp 1604681595
transform 1 0 1932 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_21
timestamp 1604681595
transform 1 0 3036 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1604681595
transform 1 0 3772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1604681595
transform 1 0 4876 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1604681595
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_39
timestamp 1604681595
transform 1 0 4692 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_45
timestamp 1604681595
transform 1 0 5244 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_48
timestamp 1604681595
transform 1 0 5520 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5336 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_52
timestamp 1604681595
transform 1 0 5888 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5704 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_56
timestamp 1604681595
transform 1 0 6256 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_55
timestamp 1604681595
transform 1 0 6164 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6348 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6072 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 6532 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_62
timestamp 1604681595
transform 1 0 6808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_62
timestamp 1604681595
transform 1 0 6808 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 7084 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8372 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_73
timestamp 1604681595
transform 1 0 7820 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_77
timestamp 1604681595
transform 1 0 8188 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_88
timestamp 1604681595
transform 1 0 9200 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_84
timestamp 1604681595
transform 1 0 8832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_100
timestamp 1604681595
transform 1 0 10304 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_102
timestamp 1604681595
transform 1 0 10488 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 10488 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_104
timestamp 1604681595
transform 1 0 10672 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_112
timestamp 1604681595
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1604681595
transform 1 0 11500 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_106
timestamp 1604681595
transform 1 0 10856 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11224 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 11224 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_116
timestamp 1604681595
transform 1 0 11776 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1604681595
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11684 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_46_134
timestamp 1604681595
transform 1 0 13432 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1604681595
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_143
timestamp 1604681595
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604681595
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604681595
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604681595
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_7
timestamp 1604681595
transform 1 0 1748 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_13
timestamp 1604681595
transform 1 0 2300 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_16
timestamp 1604681595
transform 1 0 2576 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_20
timestamp 1604681595
transform 1 0 2944 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 4692 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4232 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_25
timestamp 1604681595
transform 1 0 3404 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_32
timestamp 1604681595
transform 1 0 4048 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_36
timestamp 1604681595
transform 1 0 4416 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5704 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5152 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5520 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6808 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_42
timestamp 1604681595
transform 1 0 4968 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_46
timestamp 1604681595
transform 1 0 5336 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_59
timestamp 1604681595
transform 1 0 6532 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 8280 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 7176 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7544 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_64
timestamp 1604681595
transform 1 0 6992 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_68
timestamp 1604681595
transform 1 0 7360 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_72
timestamp 1604681595
transform 1 0 7728 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_81
timestamp 1604681595
transform 1 0 8556 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1604681595
transform 1 0 8924 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_89
timestamp 1604681595
transform 1 0 9292 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1604681595
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_97
timestamp 1604681595
transform 1 0 10028 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_104
timestamp 1604681595
transform 1 0 10672 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11224 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1604681595
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1604681595
transform 1 0 14076 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1604681595
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604681595
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604681595
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_9
timestamp 1604681595
transform 1 0 1932 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_13
timestamp 1604681595
transform 1 0 2300 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_16
timestamp 1604681595
transform 1 0 2576 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_20
timestamp 1604681595
transform 1 0 2944 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4784 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3220 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4600 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_32
timestamp 1604681595
transform 1 0 4048 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_36
timestamp 1604681595
transform 1 0 4416 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5796 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_49
timestamp 1604681595
transform 1 0 5612 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_53
timestamp 1604681595
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1604681595
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8740 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_71
timestamp 1604681595
transform 1 0 7636 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_75
timestamp 1604681595
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_79
timestamp 1604681595
transform 1 0 8372 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9476 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10672 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_85
timestamp 1604681595
transform 1 0 8924 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1604681595
transform 1 0 9292 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_102
timestamp 1604681595
transform 1 0 10488 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_106
timestamp 1604681595
transform 1 0 10856 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_118
timestamp 1604681595
transform 1 0 11960 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1604681595
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1604681595
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_143
timestamp 1604681595
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604681595
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604681595
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1604681595
transform 1 0 1380 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_7
timestamp 1604681595
transform 1 0 1748 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_13
timestamp 1604681595
transform 1 0 2300 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_23
timestamp 1604681595
transform 1 0 3220 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_27
timestamp 1604681595
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_41
timestamp 1604681595
transform 1 0 4876 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5060 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6624 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_45
timestamp 1604681595
transform 1 0 5244 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_58
timestamp 1604681595
transform 1 0 6440 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_62
timestamp 1604681595
transform 1 0 6808 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7176 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8188 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6992 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_75
timestamp 1604681595
transform 1 0 8004 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_79
timestamp 1604681595
transform 1 0 8372 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_83
timestamp 1604681595
transform 1 0 8740 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 1604681595
transform 1 0 9476 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_112
timestamp 1604681595
transform 1 0 11408 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_124
timestamp 1604681595
transform 1 0 12512 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_136
timestamp 1604681595
transform 1 0 13616 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_144
timestamp 1604681595
transform 1 0 14352 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604681595
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604681595
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2944 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_9
timestamp 1604681595
transform 1 0 1932 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_13
timestamp 1604681595
transform 1 0 2300 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_19
timestamp 1604681595
transform 1 0 2852 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 3496 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3312 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_22
timestamp 1604681595
transform 1 0 3128 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5428 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6072 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_45
timestamp 1604681595
transform 1 0 5244 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_49
timestamp 1604681595
transform 1 0 5612 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_53
timestamp 1604681595
transform 1 0 5980 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_59
timestamp 1604681595
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_62
timestamp 1604681595
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7636 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7452 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7084 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_67
timestamp 1604681595
transform 1 0 7268 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_90
timestamp 1604681595
transform 1 0 9384 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_95
timestamp 1604681595
transform 1 0 9844 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_99
timestamp 1604681595
transform 1 0 10212 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_103
timestamp 1604681595
transform 1 0 10580 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1604681595
transform 1 0 11500 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_107
timestamp 1604681595
transform 1 0 10948 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11316 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_121
timestamp 1604681595
transform 1 0 12236 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_117
timestamp 1604681595
transform 1 0 11868 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12052 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11684 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1604681595
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1604681595
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_143
timestamp 1604681595
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604681595
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604681595
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604681595
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1604681595
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1604681595
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1604681595
transform 1 0 1380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_7
timestamp 1604681595
transform 1 0 1748 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_19
timestamp 1604681595
transform 1 0 2852 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4140 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_27
timestamp 1604681595
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_32
timestamp 1604681595
transform 1 0 4048 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_31
timestamp 1604681595
transform 1 0 3956 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_39
timestamp 1604681595
transform 1 0 4692 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_48
timestamp 1604681595
transform 1 0 5520 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_44
timestamp 1604681595
transform 1 0 5152 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_50
timestamp 1604681595
transform 1 0 5704 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_42
timestamp 1604681595
transform 1 0 4968 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5336 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5796 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4968 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1604681595
transform 1 0 6348 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_53
timestamp 1604681595
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_54
timestamp 1604681595
transform 1 0 6072 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 5888 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_62
timestamp 1604681595
transform 1 0 6808 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_66
timestamp 1604681595
transform 1 0 7176 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_72
timestamp 1604681595
transform 1 0 7728 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_67
timestamp 1604681595
transform 1 0 7268 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7544 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7544 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_79
timestamp 1604681595
transform 1 0 8372 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8556 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_83
timestamp 1604681595
transform 1 0 8740 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1604681595
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_87
timestamp 1604681595
transform 1 0 9108 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_84
timestamp 1604681595
transform 1 0 8832 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9200 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 9384 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_97
timestamp 1604681595
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_102
timestamp 1604681595
transform 1 0 10488 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_114
timestamp 1604681595
transform 1 0 11592 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1604681595
transform 1 0 11224 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_110
timestamp 1604681595
transform 1 0 11224 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_106
timestamp 1604681595
transform 1 0 10856 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11408 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11316 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_123
timestamp 1604681595
transform 1 0 12420 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_119
timestamp 1604681595
transform 1 0 12052 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12604 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11868 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_120
timestamp 1604681595
transform 1 0 12144 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_132
timestamp 1604681595
transform 1 0 13248 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_144
timestamp 1604681595
transform 1 0 14352 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_127
timestamp 1604681595
transform 1 0 12788 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_139
timestamp 1604681595
transform 1 0 13892 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_145
timestamp 1604681595
transform 1 0 14444 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604681595
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604681595
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604681595
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_9
timestamp 1604681595
transform 1 0 1932 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_21
timestamp 1604681595
transform 1 0 3036 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1604681595
transform 1 0 3772 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_32
timestamp 1604681595
transform 1 0 4048 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_40
timestamp 1604681595
transform 1 0 4784 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4968 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_54_61
timestamp 1604681595
transform 1 0 6716 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6900 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7268 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8464 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_65
timestamp 1604681595
transform 1 0 7084 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_78
timestamp 1604681595
transform 1 0 8280 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1604681595
transform 1 0 8648 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_86
timestamp 1604681595
transform 1 0 9016 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_102
timestamp 1604681595
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11408 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11040 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_106
timestamp 1604681595
transform 1 0 10856 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_110
timestamp 1604681595
transform 1 0 11224 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_131
timestamp 1604681595
transform 1 0 13156 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_143
timestamp 1604681595
transform 1 0 14260 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604681595
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604681595
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1604681595
transform 1 0 1380 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1604681595
transform 1 0 1748 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_19
timestamp 1604681595
transform 1 0 2852 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 3956 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3772 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3404 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_27
timestamp 1604681595
transform 1 0 3588 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_50
timestamp 1604681595
transform 1 0 5704 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_56
timestamp 1604681595
transform 1 0 6256 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_60
timestamp 1604681595
transform 1 0 6624 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8648 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_71
timestamp 1604681595
transform 1 0 7636 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_75
timestamp 1604681595
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_79
timestamp 1604681595
transform 1 0 8372 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8832 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10488 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10304 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9936 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_93
timestamp 1604681595
transform 1 0 9660 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_98
timestamp 1604681595
transform 1 0 10120 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_111
timestamp 1604681595
transform 1 0 11316 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_115
timestamp 1604681595
transform 1 0 11684 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_118
timestamp 1604681595
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_132
timestamp 1604681595
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_136
timestamp 1604681595
transform 1 0 13616 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_144
timestamp 1604681595
transform 1 0 14352 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604681595
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604681595
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 2760 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_9
timestamp 1604681595
transform 1 0 1932 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_17
timestamp 1604681595
transform 1 0 2668 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1604681595
transform 1 0 2944 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_28
timestamp 1604681595
transform 1 0 3680 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1604681595
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1604681595
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_56
timestamp 1604681595
transform 1 0 6256 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 7820 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7452 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_67
timestamp 1604681595
transform 1 0 7268 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_71
timestamp 1604681595
transform 1 0 7636 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10304 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10120 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_84
timestamp 1604681595
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_88
timestamp 1604681595
transform 1 0 9200 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_93
timestamp 1604681595
transform 1 0 9660 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_97
timestamp 1604681595
transform 1 0 10028 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11868 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11684 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_109
timestamp 1604681595
transform 1 0 11132 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12880 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_126
timestamp 1604681595
transform 1 0 12696 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_130
timestamp 1604681595
transform 1 0 13064 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_142
timestamp 1604681595
transform 1 0 14168 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604681595
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 2760 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604681595
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 1932 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 2300 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_7
timestamp 1604681595
transform 1 0 1748 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_11
timestamp 1604681595
transform 1 0 2116 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_15
timestamp 1604681595
transform 1 0 2484 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 3312 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 4048 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_22
timestamp 1604681595
transform 1 0 3128 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_26
timestamp 1604681595
transform 1 0 3496 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_34
timestamp 1604681595
transform 1 0 4232 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 5244 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_42
timestamp 1604681595
transform 1 0 4968 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1604681595
transform 1 0 5428 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1604681595
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_81
timestamp 1604681595
transform 1 0 8556 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9568 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_89
timestamp 1604681595
transform 1 0 9292 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_94
timestamp 1604681595
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 12420 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11132 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11500 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_107
timestamp 1604681595
transform 1 0 10948 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_111
timestamp 1604681595
transform 1 0 11316 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_115
timestamp 1604681595
transform 1 0 11684 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_121
timestamp 1604681595
transform 1 0 12236 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_126
timestamp 1604681595
transform 1 0 12696 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_138
timestamp 1604681595
transform 1 0 13800 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604681595
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 2484 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 1380 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604681595
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_7
timestamp 1604681595
transform 1 0 1748 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_19
timestamp 1604681595
transform 1 0 2852 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 4048 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_36
timestamp 1604681595
transform 1 0 4416 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 6716 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 5244 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_44
timestamp 1604681595
transform 1 0 5152 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_49
timestamp 1604681595
transform 1 0 5612 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 7820 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_65
timestamp 1604681595
transform 1 0 7084 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_69
timestamp 1604681595
transform 1 0 7452 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_77
timestamp 1604681595
transform 1 0 8188 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_81
timestamp 1604681595
transform 1 0 8556 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10488 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9844 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_89
timestamp 1604681595
transform 1 0 9292 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1604681595
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_97
timestamp 1604681595
transform 1 0 10028 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_101
timestamp 1604681595
transform 1 0 10396 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1604681595
transform 1 0 12236 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_133
timestamp 1604681595
transform 1 0 13340 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_145
timestamp 1604681595
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604681595
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_3
timestamp 1604681595
transform 1 0 1380 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_7
timestamp 1604681595
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604681595
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604681595
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_19
timestamp 1604681595
transform 1 0 2852 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_11
timestamp 1604681595
transform 1 0 2116 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 2300 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 2484 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 2116 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1604681595
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1604681595
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_23
timestamp 1604681595
transform 1 0 3220 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 3036 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 3588 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_36
timestamp 1604681595
transform 1 0 4416 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_35
timestamp 1604681595
transform 1 0 4324 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_31
timestamp 1604681595
transform 1 0 3956 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 4508 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 4140 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 4048 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_39
timestamp 1604681595
transform 1 0 4692 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_48
timestamp 1604681595
transform 1 0 5520 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_46
timestamp 1604681595
transform 1 0 5336 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_43
timestamp 1604681595
transform 1 0 5060 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 5704 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 5152 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 5152 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 5520 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_56
timestamp 1604681595
transform 1 0 6256 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_52
timestamp 1604681595
transform 1 0 5888 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_59
timestamp 1604681595
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_56
timestamp 1604681595
transform 1 0 6256 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1604681595
transform 1 0 5888 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 6348 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_61
timestamp 1604681595
transform 1 0 6716 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 6808 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_70
timestamp 1604681595
transform 1 0 7544 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_66
timestamp 1604681595
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 7728 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 7360 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 7452 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_73
timestamp 1604681595
transform 1 0 7820 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_74
timestamp 1604681595
transform 1 0 7912 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 8004 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_77
timestamp 1604681595
transform 1 0 8188 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8004 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_94
timestamp 1604681595
transform 1 0 9752 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_98
timestamp 1604681595
transform 1 0 10120 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_89
timestamp 1604681595
transform 1 0 9292 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11500 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_111
timestamp 1604681595
transform 1 0 11316 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_115
timestamp 1604681595
transform 1 0 11684 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_121
timestamp 1604681595
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_123
timestamp 1604681595
transform 1 0 12420 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_112
timestamp 1604681595
transform 1 0 11408 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_124
timestamp 1604681595
transform 1 0 12512 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 13432 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_131
timestamp 1604681595
transform 1 0 13156 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_138
timestamp 1604681595
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_142
timestamp 1604681595
transform 1 0 14168 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_136
timestamp 1604681595
transform 1 0 13616 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_144
timestamp 1604681595
transform 1 0 14352 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604681595
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604681595
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604681595
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604681595
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604681595
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1604681595
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1604681595
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_51
timestamp 1604681595
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1604681595
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_62
timestamp 1604681595
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 7176 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 8280 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 7728 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_70
timestamp 1604681595
transform 1 0 7544 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_74
timestamp 1604681595
transform 1 0 7912 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_82
timestamp 1604681595
transform 1 0 8648 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 8832 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1604681595
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1604681595
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11500 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11868 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_110
timestamp 1604681595
transform 1 0 11224 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_115
timestamp 1604681595
transform 1 0 11684 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_119
timestamp 1604681595
transform 1 0 12052 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604681595
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1604681595
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_143
timestamp 1604681595
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604681595
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604681595
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604681595
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604681595
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604681595
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1604681595
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1604681595
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1604681595
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1604681595
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_80
timestamp 1604681595
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604681595
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11500 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_62_105
timestamp 1604681595
transform 1 0 10764 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_132
timestamp 1604681595
transform 1 0 13248 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_144
timestamp 1604681595
transform 1 0 14352 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604681595
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604681595
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604681595
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604681595
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604681595
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604681595
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604681595
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604681595
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604681595
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604681595
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604681595
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604681595
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604681595
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604681595
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1604681595
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_143
timestamp 1604681595
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604681595
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604681595
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604681595
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604681595
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604681595
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604681595
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604681595
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604681595
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604681595
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604681595
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604681595
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604681595
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604681595
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604681595
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604681595
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_137
timestamp 1604681595
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1604681595
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604681595
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 2864 480 2984 6 ccff_head
port 0 nsew default input
rlabel metal3 s 15520 9936 16000 10056 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 15520 23264 16000 23384 6 gfpga_pad_EMBEDDED_IO_SOC_DIR
port 82 nsew default tristate
rlabel metal3 s 15520 29928 16000 30048 6 gfpga_pad_EMBEDDED_IO_SOC_IN
port 83 nsew default input
rlabel metal3 s 15520 36592 16000 36712 6 gfpga_pad_EMBEDDED_IO_SOC_OUT
port 84 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 left_grid_pin_16_
port 85 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 left_grid_pin_17_
port 86 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 left_grid_pin_18_
port 87 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 left_grid_pin_19_
port 88 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 left_grid_pin_20_
port 89 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 left_grid_pin_21_
port 90 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 left_grid_pin_22_
port 91 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 left_grid_pin_23_
port 92 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 left_grid_pin_24_
port 93 nsew default tristate
rlabel metal3 s 0 22856 480 22976 6 left_grid_pin_25_
port 94 nsew default tristate
rlabel metal3 s 0 24896 480 25016 6 left_grid_pin_26_
port 95 nsew default tristate
rlabel metal3 s 0 26936 480 27056 6 left_grid_pin_27_
port 96 nsew default tristate
rlabel metal3 s 0 28840 480 28960 6 left_grid_pin_28_
port 97 nsew default tristate
rlabel metal3 s 0 30880 480 31000 6 left_grid_pin_29_
port 98 nsew default tristate
rlabel metal3 s 0 32920 480 33040 6 left_grid_pin_30_
port 99 nsew default tristate
rlabel metal3 s 0 34824 480 34944 6 left_grid_pin_31_
port 100 nsew default tristate
rlabel metal3 s 0 36864 480 36984 6 left_width_0_height_0__pin_0_
port 101 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_width_0_height_0__pin_1_lower
port 102 nsew default tristate
rlabel metal3 s 0 38904 480 39024 6 left_width_0_height_0__pin_1_upper
port 103 nsew default tristate
rlabel metal3 s 15520 3272 16000 3392 6 prog_clk
port 104 nsew default input
rlabel metal3 s 15520 16600 16000 16720 6 right_grid_pin_0_
port 105 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 VPWR
port 106 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 VGND
port 107 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
