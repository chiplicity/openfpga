magic
tech EFS8A
magscale 1 2
timestamp 1602874268
<< locali >>
rect 4899 5015 4933 5083
rect 4899 4981 4905 5015
rect 35627 4777 35633 4811
rect 57247 4777 57253 4811
rect 66171 4777 66177 4811
rect 79235 4777 79241 4811
rect 35627 4709 35661 4777
rect 57247 4709 57281 4777
rect 66171 4709 66205 4777
rect 79235 4709 79269 4777
<< viali >>
rect 37933 6613 37967 6647
rect 37105 6273 37139 6307
rect 37841 6205 37875 6239
rect 38301 6205 38335 6239
rect 38577 6205 38611 6239
rect 38945 6205 38979 6239
rect 77309 6205 77343 6239
rect 77769 6205 77803 6239
rect 37473 6137 37507 6171
rect 36737 6069 36771 6103
rect 37657 6069 37691 6103
rect 77493 6069 77527 6103
rect 37841 5865 37875 5899
rect 60473 5865 60507 5899
rect 63141 5865 63175 5899
rect 77493 5865 77527 5899
rect 51825 5797 51859 5831
rect 60565 5797 60599 5831
rect 63233 5797 63267 5831
rect 38025 5729 38059 5763
rect 38393 5729 38427 5763
rect 38577 5729 38611 5763
rect 39129 5729 39163 5763
rect 51273 5729 51307 5763
rect 60381 5729 60415 5763
rect 63049 5729 63083 5763
rect 68845 5729 68879 5763
rect 37565 5661 37599 5695
rect 60197 5661 60231 5695
rect 60933 5661 60967 5695
rect 62865 5661 62899 5695
rect 63601 5661 63635 5695
rect 68753 5661 68787 5695
rect 87889 5525 87923 5559
rect 37841 5321 37875 5355
rect 39773 5321 39807 5355
rect 59829 5321 59863 5355
rect 60933 5321 60967 5355
rect 63509 5321 63543 5355
rect 76849 5321 76883 5355
rect 60289 5253 60323 5287
rect 18061 5185 18095 5219
rect 51181 5185 51215 5219
rect 62773 5185 62807 5219
rect 77401 5185 77435 5219
rect 2237 5117 2271 5151
rect 4537 5117 4571 5151
rect 38209 5117 38243 5151
rect 38485 5117 38519 5151
rect 38761 5117 38795 5151
rect 39129 5117 39163 5151
rect 77677 5117 77711 5151
rect 87613 5117 87647 5151
rect 88073 5117 88107 5151
rect 2145 5049 2179 5083
rect 2599 5049 2633 5083
rect 18382 5049 18416 5083
rect 37105 5049 37139 5083
rect 37473 5049 37507 5083
rect 63233 5049 63267 5083
rect 77217 5049 77251 5083
rect 77769 5049 77803 5083
rect 78137 5049 78171 5083
rect 87797 5049 87831 5083
rect 88165 5049 88199 5083
rect 88533 5049 88567 5083
rect 3157 4981 3191 5015
rect 4445 4981 4479 5015
rect 4905 4981 4939 5015
rect 5457 4981 5491 5015
rect 17785 4981 17819 5015
rect 18981 4981 19015 5015
rect 36737 4981 36771 5015
rect 38025 4981 38059 5015
rect 60565 4981 60599 5015
rect 68845 4981 68879 5015
rect 77585 4981 77619 5015
rect 87245 4981 87279 5015
rect 87981 4981 88015 5015
rect 1685 4777 1719 4811
rect 4537 4777 4571 4811
rect 18061 4777 18095 4811
rect 35633 4777 35667 4811
rect 37565 4777 37599 4811
rect 37841 4777 37875 4811
rect 57253 4777 57287 4811
rect 62865 4777 62899 4811
rect 66177 4777 66211 4811
rect 77401 4777 77435 4811
rect 79241 4777 79275 4811
rect 87889 4777 87923 4811
rect 37197 4709 37231 4743
rect 49893 4709 49927 4743
rect 88619 4709 88653 4743
rect 38025 4641 38059 4675
rect 38393 4641 38427 4675
rect 38577 4641 38611 4675
rect 39129 4641 39163 4675
rect 49985 4641 50019 4675
rect 65809 4641 65843 4675
rect 78873 4641 78907 4675
rect 35265 4573 35299 4607
rect 56885 4573 56919 4607
rect 88257 4573 88291 4607
rect 2329 4437 2363 4471
rect 36185 4437 36219 4471
rect 57805 4437 57839 4471
rect 66729 4437 66763 4471
rect 79793 4437 79827 4471
rect 89177 4437 89211 4471
rect 2053 4233 2087 4267
rect 35725 4233 35759 4267
rect 38209 4233 38243 4267
rect 57621 4233 57655 4267
rect 66177 4233 66211 4267
rect 79241 4233 79275 4267
rect 88625 4233 88659 4267
rect 37473 4165 37507 4199
rect 37841 4165 37875 4199
rect 38577 4165 38611 4199
rect 88349 4165 88383 4199
rect 1593 4097 1627 4131
rect 7021 4097 7055 4131
rect 20177 4097 20211 4131
rect 20913 4097 20947 4131
rect 1409 4029 1443 4063
rect 6653 4029 6687 4063
rect 6837 4029 6871 4063
rect 20729 4029 20763 4063
rect 7481 3893 7515 3927
rect 20637 3893 20671 3927
rect 21373 3893 21407 3927
rect 35265 3893 35299 3927
rect 49985 3893 50019 3927
rect 56885 3893 56919 3927
rect 65809 3893 65843 3927
rect 78965 3893 78999 3927
rect 6929 3689 6963 3723
rect 53021 3689 53055 3723
rect 36277 3553 36311 3587
rect 52561 3553 52595 3587
rect 64429 3553 64463 3587
rect 78229 3553 78263 3587
rect 88257 3553 88291 3587
rect 36093 3485 36127 3519
rect 52377 3485 52411 3519
rect 64245 3485 64279 3519
rect 78045 3485 78079 3519
rect 88441 3485 88475 3519
rect 1685 3349 1719 3383
rect 36737 3349 36771 3383
rect 64889 3349 64923 3383
rect 78689 3349 78723 3383
rect 88901 3349 88935 3383
rect 2053 3145 2087 3179
rect 36461 3145 36495 3179
rect 52745 3145 52779 3179
rect 64705 3145 64739 3179
rect 78505 3145 78539 3179
rect 80713 3145 80747 3179
rect 87981 3145 88015 3179
rect 89085 3145 89119 3179
rect 1409 2941 1443 2975
rect 12449 2941 12483 2975
rect 13001 2941 13035 2975
rect 25513 2941 25547 2975
rect 80069 2941 80103 2975
rect 88073 2941 88107 2975
rect 78137 2873 78171 2907
rect 1593 2805 1627 2839
rect 12633 2805 12667 2839
rect 25697 2805 25731 2839
rect 26157 2805 26191 2839
rect 36185 2805 36219 2839
rect 52469 2805 52503 2839
rect 64337 2805 64371 2839
rect 80253 2805 80287 2839
rect 88257 2805 88291 2839
rect 88717 2805 88751 2839
rect 53941 2601 53975 2635
rect 67005 2601 67039 2635
rect 67465 2601 67499 2635
rect 39313 2465 39347 2499
rect 39865 2465 39899 2499
rect 53297 2465 53331 2499
rect 66821 2465 66855 2499
rect 39497 2261 39531 2295
rect 53481 2261 53515 2295
<< metal1 >>
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 20162 13512 20168 13524
rect 19392 13484 20168 13512
rect 19392 13472 19398 13484
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 33134 13472 33140 13524
rect 33192 13512 33198 13524
rect 33686 13512 33692 13524
rect 33192 13484 33692 13512
rect 33192 13472 33198 13484
rect 33686 13472 33692 13484
rect 33744 13472 33750 13524
rect 86954 13472 86960 13524
rect 87012 13512 87018 13524
rect 87690 13512 87696 13524
rect 87012 13484 87696 13512
rect 87012 13472 87018 13484
rect 87690 13472 87696 13484
rect 87748 13472 87754 13524
rect 1104 11450 106812 11472
rect 1104 11398 36982 11450
rect 37034 11398 37046 11450
rect 37098 11398 37110 11450
rect 37162 11398 37174 11450
rect 37226 11398 72982 11450
rect 73034 11398 73046 11450
rect 73098 11398 73110 11450
rect 73162 11398 73174 11450
rect 73226 11398 106812 11450
rect 1104 11376 106812 11398
rect 1104 10906 106812 10928
rect 1104 10854 18982 10906
rect 19034 10854 19046 10906
rect 19098 10854 19110 10906
rect 19162 10854 19174 10906
rect 19226 10854 54982 10906
rect 55034 10854 55046 10906
rect 55098 10854 55110 10906
rect 55162 10854 55174 10906
rect 55226 10854 90982 10906
rect 91034 10854 91046 10906
rect 91098 10854 91110 10906
rect 91162 10854 91174 10906
rect 91226 10854 106812 10906
rect 1104 10832 106812 10854
rect 1104 10362 106812 10384
rect 1104 10310 36982 10362
rect 37034 10310 37046 10362
rect 37098 10310 37110 10362
rect 37162 10310 37174 10362
rect 37226 10310 72982 10362
rect 73034 10310 73046 10362
rect 73098 10310 73110 10362
rect 73162 10310 73174 10362
rect 73226 10310 106812 10362
rect 1104 10288 106812 10310
rect 1104 9818 106812 9840
rect 1104 9766 18982 9818
rect 19034 9766 19046 9818
rect 19098 9766 19110 9818
rect 19162 9766 19174 9818
rect 19226 9766 54982 9818
rect 55034 9766 55046 9818
rect 55098 9766 55110 9818
rect 55162 9766 55174 9818
rect 55226 9766 90982 9818
rect 91034 9766 91046 9818
rect 91098 9766 91110 9818
rect 91162 9766 91174 9818
rect 91226 9766 106812 9818
rect 1104 9744 106812 9766
rect 73338 9324 73344 9376
rect 73396 9364 73402 9376
rect 74166 9364 74172 9376
rect 73396 9336 74172 9364
rect 73396 9324 73402 9336
rect 74166 9324 74172 9336
rect 74224 9324 74230 9376
rect 1104 9274 106812 9296
rect 1104 9222 36982 9274
rect 37034 9222 37046 9274
rect 37098 9222 37110 9274
rect 37162 9222 37174 9274
rect 37226 9222 72982 9274
rect 73034 9222 73046 9274
rect 73098 9222 73110 9274
rect 73162 9222 73174 9274
rect 73226 9222 106812 9274
rect 1104 9200 106812 9222
rect 1104 8730 106812 8752
rect 1104 8678 18982 8730
rect 19034 8678 19046 8730
rect 19098 8678 19110 8730
rect 19162 8678 19174 8730
rect 19226 8678 54982 8730
rect 55034 8678 55046 8730
rect 55098 8678 55110 8730
rect 55162 8678 55174 8730
rect 55226 8678 90982 8730
rect 91034 8678 91046 8730
rect 91098 8678 91110 8730
rect 91162 8678 91174 8730
rect 91226 8678 106812 8730
rect 1104 8656 106812 8678
rect 1104 8186 106812 8208
rect 1104 8134 36982 8186
rect 37034 8134 37046 8186
rect 37098 8134 37110 8186
rect 37162 8134 37174 8186
rect 37226 8134 72982 8186
rect 73034 8134 73046 8186
rect 73098 8134 73110 8186
rect 73162 8134 73174 8186
rect 73226 8134 106812 8186
rect 1104 8112 106812 8134
rect 1104 7642 106812 7664
rect 1104 7590 18982 7642
rect 19034 7590 19046 7642
rect 19098 7590 19110 7642
rect 19162 7590 19174 7642
rect 19226 7590 54982 7642
rect 55034 7590 55046 7642
rect 55098 7590 55110 7642
rect 55162 7590 55174 7642
rect 55226 7590 90982 7642
rect 91034 7590 91046 7642
rect 91098 7590 91110 7642
rect 91162 7590 91174 7642
rect 91226 7590 106812 7642
rect 1104 7568 106812 7590
rect 1104 7098 106812 7120
rect 1104 7046 36982 7098
rect 37034 7046 37046 7098
rect 37098 7046 37110 7098
rect 37162 7046 37174 7098
rect 37226 7046 72982 7098
rect 73034 7046 73046 7098
rect 73098 7046 73110 7098
rect 73162 7046 73174 7098
rect 73226 7046 106812 7098
rect 1104 7024 106812 7046
rect 37918 6644 37924 6656
rect 37879 6616 37924 6644
rect 37918 6604 37924 6616
rect 37976 6604 37982 6656
rect 1104 6554 106812 6576
rect 1104 6502 18982 6554
rect 19034 6502 19046 6554
rect 19098 6502 19110 6554
rect 19162 6502 19174 6554
rect 19226 6502 54982 6554
rect 55034 6502 55046 6554
rect 55098 6502 55110 6554
rect 55162 6502 55174 6554
rect 55226 6502 90982 6554
rect 91034 6502 91046 6554
rect 91098 6502 91110 6554
rect 91162 6502 91174 6554
rect 91226 6502 106812 6554
rect 1104 6480 106812 6502
rect 37093 6307 37151 6313
rect 37093 6273 37105 6307
rect 37139 6304 37151 6307
rect 37139 6276 38608 6304
rect 37139 6273 37151 6276
rect 37093 6267 37151 6273
rect 38580 6248 38608 6276
rect 37829 6239 37887 6245
rect 37829 6205 37841 6239
rect 37875 6236 37887 6239
rect 37918 6236 37924 6248
rect 37875 6208 37924 6236
rect 37875 6205 37887 6208
rect 37829 6199 37887 6205
rect 37918 6196 37924 6208
rect 37976 6196 37982 6248
rect 38289 6239 38347 6245
rect 38289 6205 38301 6239
rect 38335 6236 38347 6239
rect 38378 6236 38384 6248
rect 38335 6208 38384 6236
rect 38335 6205 38347 6208
rect 38289 6199 38347 6205
rect 38378 6196 38384 6208
rect 38436 6196 38442 6248
rect 38562 6236 38568 6248
rect 38523 6208 38568 6236
rect 38562 6196 38568 6208
rect 38620 6196 38626 6248
rect 38933 6239 38991 6245
rect 38933 6205 38945 6239
rect 38979 6236 38991 6239
rect 39206 6236 39212 6248
rect 38979 6208 39212 6236
rect 38979 6205 38991 6208
rect 38933 6199 38991 6205
rect 37461 6171 37519 6177
rect 37461 6137 37473 6171
rect 37507 6168 37519 6171
rect 38948 6168 38976 6199
rect 39206 6196 39212 6208
rect 39264 6196 39270 6248
rect 63126 6196 63132 6248
rect 63184 6236 63190 6248
rect 77297 6239 77355 6245
rect 77297 6236 77309 6239
rect 63184 6208 77309 6236
rect 63184 6196 63190 6208
rect 77297 6205 77309 6208
rect 77343 6236 77355 6239
rect 77754 6236 77760 6248
rect 77343 6208 77760 6236
rect 77343 6205 77355 6208
rect 77297 6199 77355 6205
rect 77754 6196 77760 6208
rect 77812 6196 77818 6248
rect 37507 6140 38976 6168
rect 37507 6137 37519 6140
rect 37461 6131 37519 6137
rect 36722 6100 36728 6112
rect 36683 6072 36728 6100
rect 36722 6060 36728 6072
rect 36780 6060 36786 6112
rect 37642 6100 37648 6112
rect 37603 6072 37648 6100
rect 37642 6060 37648 6072
rect 37700 6060 37706 6112
rect 77478 6100 77484 6112
rect 77439 6072 77484 6100
rect 77478 6060 77484 6072
rect 77536 6060 77542 6112
rect 1104 6010 106812 6032
rect 1104 5958 36982 6010
rect 37034 5958 37046 6010
rect 37098 5958 37110 6010
rect 37162 5958 37174 6010
rect 37226 5958 72982 6010
rect 73034 5958 73046 6010
rect 73098 5958 73110 6010
rect 73162 5958 73174 6010
rect 73226 5958 106812 6010
rect 1104 5936 106812 5958
rect 37826 5896 37832 5908
rect 37787 5868 37832 5896
rect 37826 5856 37832 5868
rect 37884 5856 37890 5908
rect 38102 5896 38108 5908
rect 38028 5868 38108 5896
rect 38028 5769 38056 5868
rect 38102 5856 38108 5868
rect 38160 5856 38166 5908
rect 60274 5856 60280 5908
rect 60332 5896 60338 5908
rect 60461 5899 60519 5905
rect 60461 5896 60473 5899
rect 60332 5868 60473 5896
rect 60332 5856 60338 5868
rect 60461 5865 60473 5868
rect 60507 5896 60519 5899
rect 63126 5896 63132 5908
rect 60507 5868 63132 5896
rect 60507 5865 60519 5868
rect 60461 5859 60519 5865
rect 63126 5856 63132 5868
rect 63184 5856 63190 5908
rect 77478 5896 77484 5908
rect 77439 5868 77484 5896
rect 77478 5856 77484 5868
rect 77536 5856 77542 5908
rect 51810 5828 51816 5840
rect 51771 5800 51816 5828
rect 51810 5788 51816 5800
rect 51868 5788 51874 5840
rect 59814 5788 59820 5840
rect 59872 5828 59878 5840
rect 60553 5831 60611 5837
rect 60553 5828 60565 5831
rect 59872 5800 60565 5828
rect 59872 5788 59878 5800
rect 60553 5797 60565 5800
rect 60599 5828 60611 5831
rect 62850 5828 62856 5840
rect 60599 5800 62856 5828
rect 60599 5797 60611 5800
rect 60553 5791 60611 5797
rect 62850 5788 62856 5800
rect 62908 5828 62914 5840
rect 63221 5831 63279 5837
rect 63221 5828 63233 5831
rect 62908 5800 63233 5828
rect 62908 5788 62914 5800
rect 63221 5797 63233 5800
rect 63267 5797 63279 5831
rect 63221 5791 63279 5797
rect 38013 5763 38071 5769
rect 38013 5729 38025 5763
rect 38059 5729 38071 5763
rect 38378 5760 38384 5772
rect 38339 5732 38384 5760
rect 38013 5723 38071 5729
rect 38378 5720 38384 5732
rect 38436 5720 38442 5772
rect 38562 5760 38568 5772
rect 38523 5732 38568 5760
rect 38562 5720 38568 5732
rect 38620 5720 38626 5772
rect 39114 5760 39120 5772
rect 39075 5732 39120 5760
rect 39114 5720 39120 5732
rect 39172 5720 39178 5772
rect 51261 5763 51319 5769
rect 51261 5729 51273 5763
rect 51307 5729 51319 5763
rect 60366 5760 60372 5772
rect 60327 5732 60372 5760
rect 51261 5723 51319 5729
rect 37550 5692 37556 5704
rect 37463 5664 37556 5692
rect 37550 5652 37556 5664
rect 37608 5692 37614 5704
rect 39132 5692 39160 5720
rect 37608 5664 39160 5692
rect 37608 5652 37614 5664
rect 51166 5652 51172 5704
rect 51224 5692 51230 5704
rect 51276 5692 51304 5723
rect 60366 5720 60372 5732
rect 60424 5720 60430 5772
rect 62758 5720 62764 5772
rect 62816 5760 62822 5772
rect 63037 5763 63095 5769
rect 63037 5760 63049 5763
rect 62816 5732 63049 5760
rect 62816 5720 62822 5732
rect 63037 5729 63049 5732
rect 63083 5729 63095 5763
rect 68830 5760 68836 5772
rect 68791 5732 68836 5760
rect 63037 5723 63095 5729
rect 68830 5720 68836 5732
rect 68888 5720 68894 5772
rect 60182 5692 60188 5704
rect 51224 5664 51304 5692
rect 60143 5664 60188 5692
rect 51224 5652 51230 5664
rect 60182 5652 60188 5664
rect 60240 5652 60246 5704
rect 60918 5692 60924 5704
rect 60879 5664 60924 5692
rect 60918 5652 60924 5664
rect 60976 5652 60982 5704
rect 62853 5695 62911 5701
rect 62853 5661 62865 5695
rect 62899 5692 62911 5695
rect 63218 5692 63224 5704
rect 62899 5664 63224 5692
rect 62899 5661 62911 5664
rect 62853 5655 62911 5661
rect 63218 5652 63224 5664
rect 63276 5652 63282 5704
rect 63586 5692 63592 5704
rect 63547 5664 63592 5692
rect 63586 5652 63592 5664
rect 63644 5652 63650 5704
rect 68738 5692 68744 5704
rect 68699 5664 68744 5692
rect 68738 5652 68744 5664
rect 68796 5652 68802 5704
rect 87877 5559 87935 5565
rect 87877 5525 87889 5559
rect 87923 5556 87935 5559
rect 88150 5556 88156 5568
rect 87923 5528 88156 5556
rect 87923 5525 87935 5528
rect 87877 5519 87935 5525
rect 88150 5516 88156 5528
rect 88208 5516 88214 5568
rect 1104 5466 106812 5488
rect 1104 5414 18982 5466
rect 19034 5414 19046 5466
rect 19098 5414 19110 5466
rect 19162 5414 19174 5466
rect 19226 5414 54982 5466
rect 55034 5414 55046 5466
rect 55098 5414 55110 5466
rect 55162 5414 55174 5466
rect 55226 5414 90982 5466
rect 91034 5414 91046 5466
rect 91098 5414 91110 5466
rect 91162 5414 91174 5466
rect 91226 5414 106812 5466
rect 1104 5392 106812 5414
rect 37829 5355 37887 5361
rect 37829 5321 37841 5355
rect 37875 5352 37887 5355
rect 38102 5352 38108 5364
rect 37875 5324 38108 5352
rect 37875 5321 37887 5324
rect 37829 5315 37887 5321
rect 38102 5312 38108 5324
rect 38160 5312 38166 5364
rect 39758 5352 39764 5364
rect 39719 5324 39764 5352
rect 39758 5312 39764 5324
rect 39816 5312 39822 5364
rect 59814 5352 59820 5364
rect 59775 5324 59820 5352
rect 59814 5312 59820 5324
rect 59872 5312 59878 5364
rect 60182 5312 60188 5364
rect 60240 5352 60246 5364
rect 60921 5355 60979 5361
rect 60921 5352 60933 5355
rect 60240 5324 60933 5352
rect 60240 5312 60246 5324
rect 60921 5321 60933 5324
rect 60967 5352 60979 5355
rect 61010 5352 61016 5364
rect 60967 5324 61016 5352
rect 60967 5321 60979 5324
rect 60921 5315 60979 5321
rect 61010 5312 61016 5324
rect 61068 5312 61074 5364
rect 63126 5312 63132 5364
rect 63184 5352 63190 5364
rect 63497 5355 63555 5361
rect 63497 5352 63509 5355
rect 63184 5324 63509 5352
rect 63184 5312 63190 5324
rect 63497 5321 63509 5324
rect 63543 5321 63555 5355
rect 63497 5315 63555 5321
rect 68738 5312 68744 5364
rect 68796 5352 68802 5364
rect 76837 5355 76895 5361
rect 76837 5352 76849 5355
rect 68796 5324 76849 5352
rect 68796 5312 68802 5324
rect 76837 5321 76849 5324
rect 76883 5321 76895 5355
rect 76837 5315 76895 5321
rect 60274 5284 60280 5296
rect 60235 5256 60280 5284
rect 60274 5244 60280 5256
rect 60332 5244 60338 5296
rect 18046 5216 18052 5228
rect 18007 5188 18052 5216
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 37918 5176 37924 5228
rect 37976 5216 37982 5228
rect 39758 5216 39764 5228
rect 37976 5188 39764 5216
rect 37976 5176 37982 5188
rect 2225 5151 2283 5157
rect 2225 5117 2237 5151
rect 2271 5148 2283 5151
rect 2314 5148 2320 5160
rect 2271 5120 2320 5148
rect 2271 5117 2283 5120
rect 2225 5111 2283 5117
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 4522 5148 4528 5160
rect 4483 5120 4528 5148
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 38212 5157 38240 5188
rect 39758 5176 39764 5188
rect 39816 5176 39822 5228
rect 51166 5216 51172 5228
rect 51127 5188 51172 5216
rect 51166 5176 51172 5188
rect 51224 5176 51230 5228
rect 62758 5216 62764 5228
rect 62086 5188 62764 5216
rect 38197 5151 38255 5157
rect 38197 5117 38209 5151
rect 38243 5117 38255 5151
rect 38470 5148 38476 5160
rect 38431 5120 38476 5148
rect 38197 5111 38255 5117
rect 38470 5108 38476 5120
rect 38528 5108 38534 5160
rect 38562 5108 38568 5160
rect 38620 5148 38626 5160
rect 38749 5151 38807 5157
rect 38749 5148 38761 5151
rect 38620 5120 38761 5148
rect 38620 5108 38626 5120
rect 38749 5117 38761 5120
rect 38795 5117 38807 5151
rect 39114 5148 39120 5160
rect 39075 5120 39120 5148
rect 38749 5111 38807 5117
rect 39114 5108 39120 5120
rect 39172 5108 39178 5160
rect 62086 5148 62114 5188
rect 62758 5176 62764 5188
rect 62816 5176 62822 5228
rect 60568 5120 62114 5148
rect 76852 5148 76880 5315
rect 77389 5219 77447 5225
rect 77389 5185 77401 5219
rect 77435 5216 77447 5219
rect 77478 5216 77484 5228
rect 77435 5188 77484 5216
rect 77435 5185 77447 5188
rect 77389 5179 77447 5185
rect 77478 5176 77484 5188
rect 77536 5216 77542 5228
rect 79410 5216 79416 5228
rect 77536 5188 79416 5216
rect 77536 5176 77542 5188
rect 79410 5176 79416 5188
rect 79468 5176 79474 5228
rect 77665 5151 77723 5157
rect 77665 5148 77677 5151
rect 76852 5120 77677 5148
rect 2133 5083 2191 5089
rect 2133 5049 2145 5083
rect 2179 5080 2191 5083
rect 2587 5083 2645 5089
rect 2587 5080 2599 5083
rect 2179 5052 2599 5080
rect 2179 5049 2191 5052
rect 2133 5043 2191 5049
rect 2587 5049 2599 5052
rect 2633 5080 2645 5083
rect 18370 5083 18428 5089
rect 2633 5052 4476 5080
rect 2633 5049 2645 5052
rect 2587 5043 2645 5049
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 4448 5021 4476 5052
rect 18370 5049 18382 5083
rect 18416 5049 18428 5083
rect 18370 5043 18428 5049
rect 37093 5083 37151 5089
rect 37093 5049 37105 5083
rect 37139 5080 37151 5083
rect 37461 5083 37519 5089
rect 37461 5080 37473 5083
rect 37139 5052 37473 5080
rect 37139 5049 37151 5052
rect 37093 5043 37151 5049
rect 37461 5049 37473 5052
rect 37507 5080 37519 5083
rect 38580 5080 38608 5108
rect 37507 5052 38608 5080
rect 37507 5049 37519 5052
rect 37461 5043 37519 5049
rect 3145 5015 3203 5021
rect 3145 5012 3157 5015
rect 1728 4984 3157 5012
rect 1728 4972 1734 4984
rect 3145 4981 3157 4984
rect 3191 4981 3203 5015
rect 3145 4975 3203 4981
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 4890 5012 4896 5024
rect 4479 4984 4896 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5442 5012 5448 5024
rect 5403 4984 5448 5012
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 5012 17834 5024
rect 18385 5012 18413 5043
rect 17828 4984 18413 5012
rect 17828 4972 17834 4984
rect 18874 4972 18880 5024
rect 18932 5012 18938 5024
rect 18969 5015 19027 5021
rect 18969 5012 18981 5015
rect 18932 4984 18981 5012
rect 18932 4972 18938 4984
rect 18969 4981 18981 4984
rect 19015 4981 19027 5015
rect 36722 5012 36728 5024
rect 36683 4984 36728 5012
rect 18969 4975 19027 4981
rect 36722 4972 36728 4984
rect 36780 4972 36786 5024
rect 38010 5012 38016 5024
rect 37971 4984 38016 5012
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 60366 4972 60372 5024
rect 60424 5012 60430 5024
rect 60568 5021 60596 5120
rect 77665 5117 77677 5120
rect 77711 5117 77723 5151
rect 77665 5111 77723 5117
rect 77846 5108 77852 5160
rect 77904 5148 77910 5160
rect 87601 5151 87659 5157
rect 87601 5148 87613 5151
rect 77904 5120 87613 5148
rect 77904 5108 77910 5120
rect 87601 5117 87613 5120
rect 87647 5148 87659 5151
rect 88058 5148 88064 5160
rect 87647 5120 88064 5148
rect 87647 5117 87659 5120
rect 87601 5111 87659 5117
rect 88058 5108 88064 5120
rect 88116 5108 88122 5160
rect 63218 5080 63224 5092
rect 63131 5052 63224 5080
rect 63218 5040 63224 5052
rect 63276 5080 63282 5092
rect 63276 5052 68876 5080
rect 63276 5040 63282 5052
rect 68848 5024 68876 5052
rect 72786 5040 72792 5092
rect 72844 5080 72850 5092
rect 77205 5083 77263 5089
rect 77205 5080 77217 5083
rect 72844 5052 77217 5080
rect 72844 5040 72850 5052
rect 77205 5049 77217 5052
rect 77251 5049 77263 5083
rect 77205 5043 77263 5049
rect 60553 5015 60611 5021
rect 60553 5012 60565 5015
rect 60424 4984 60565 5012
rect 60424 4972 60430 4984
rect 60553 4981 60565 4984
rect 60599 4981 60611 5015
rect 68830 5012 68836 5024
rect 68791 4984 68836 5012
rect 60553 4975 60611 4981
rect 68830 4972 68836 4984
rect 68888 4972 68894 5024
rect 77220 5012 77248 5043
rect 77478 5040 77484 5092
rect 77536 5080 77542 5092
rect 77757 5083 77815 5089
rect 77757 5080 77769 5083
rect 77536 5052 77769 5080
rect 77536 5040 77542 5052
rect 77757 5049 77769 5052
rect 77803 5049 77815 5083
rect 78122 5080 78128 5092
rect 78083 5052 78128 5080
rect 77757 5043 77815 5049
rect 78122 5040 78128 5052
rect 78180 5040 78186 5092
rect 87138 5080 87144 5092
rect 78232 5052 87144 5080
rect 77573 5015 77631 5021
rect 77573 5012 77585 5015
rect 77220 4984 77585 5012
rect 77573 4981 77585 4984
rect 77619 5012 77631 5015
rect 78232 5012 78260 5052
rect 87138 5040 87144 5052
rect 87196 5040 87202 5092
rect 87785 5083 87843 5089
rect 87785 5080 87797 5083
rect 87248 5052 87797 5080
rect 77619 4984 78260 5012
rect 77619 4981 77631 4984
rect 77573 4975 77631 4981
rect 79410 4972 79416 5024
rect 79468 5012 79474 5024
rect 87248 5021 87276 5052
rect 87785 5049 87797 5052
rect 87831 5049 87843 5083
rect 88150 5080 88156 5092
rect 88111 5052 88156 5080
rect 87785 5043 87843 5049
rect 88150 5040 88156 5052
rect 88208 5040 88214 5092
rect 88521 5083 88579 5089
rect 88521 5049 88533 5083
rect 88567 5080 88579 5083
rect 88610 5080 88616 5092
rect 88567 5052 88616 5080
rect 88567 5049 88579 5052
rect 88521 5043 88579 5049
rect 88610 5040 88616 5052
rect 88668 5040 88674 5092
rect 87233 5015 87291 5021
rect 87233 5012 87245 5015
rect 79468 4984 87245 5012
rect 79468 4972 79474 4984
rect 87233 4981 87245 4984
rect 87279 4981 87291 5015
rect 87966 5012 87972 5024
rect 87927 4984 87972 5012
rect 87233 4975 87291 4981
rect 87966 4972 87972 4984
rect 88024 4972 88030 5024
rect 1104 4922 106812 4944
rect 1104 4870 36982 4922
rect 37034 4870 37046 4922
rect 37098 4870 37110 4922
rect 37162 4870 37174 4922
rect 37226 4870 72982 4922
rect 73034 4870 73046 4922
rect 73098 4870 73110 4922
rect 73162 4870 73174 4922
rect 73226 4870 106812 4922
rect 1104 4848 106812 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 18046 4808 18052 4820
rect 18007 4780 18052 4808
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 35250 4768 35256 4820
rect 35308 4808 35314 4820
rect 35621 4811 35679 4817
rect 35621 4808 35633 4811
rect 35308 4780 35633 4808
rect 35308 4768 35314 4780
rect 35621 4777 35633 4780
rect 35667 4777 35679 4811
rect 37550 4808 37556 4820
rect 37511 4780 37556 4808
rect 35621 4771 35679 4777
rect 37550 4768 37556 4780
rect 37608 4768 37614 4820
rect 37826 4808 37832 4820
rect 37787 4780 37832 4808
rect 37826 4768 37832 4780
rect 37884 4768 37890 4820
rect 56870 4768 56876 4820
rect 56928 4808 56934 4820
rect 57241 4811 57299 4817
rect 57241 4808 57253 4811
rect 56928 4780 57253 4808
rect 56928 4768 56934 4780
rect 57241 4777 57253 4780
rect 57287 4777 57299 4811
rect 62850 4808 62856 4820
rect 62811 4780 62856 4808
rect 57241 4771 57299 4777
rect 62850 4768 62856 4780
rect 62908 4768 62914 4820
rect 65794 4768 65800 4820
rect 65852 4808 65858 4820
rect 66165 4811 66223 4817
rect 66165 4808 66177 4811
rect 65852 4780 66177 4808
rect 65852 4768 65858 4780
rect 66165 4777 66177 4780
rect 66211 4777 66223 4811
rect 77386 4808 77392 4820
rect 77347 4780 77392 4808
rect 66165 4771 66223 4777
rect 77386 4768 77392 4780
rect 77444 4768 77450 4820
rect 78950 4768 78956 4820
rect 79008 4808 79014 4820
rect 79229 4811 79287 4817
rect 79229 4808 79241 4811
rect 79008 4780 79241 4808
rect 79008 4768 79014 4780
rect 79229 4777 79241 4780
rect 79275 4777 79287 4811
rect 79229 4771 79287 4777
rect 87138 4768 87144 4820
rect 87196 4808 87202 4820
rect 87877 4811 87935 4817
rect 87877 4808 87889 4811
rect 87196 4780 87889 4808
rect 87196 4768 87202 4780
rect 87877 4777 87889 4780
rect 87923 4808 87935 4811
rect 87966 4808 87972 4820
rect 87923 4780 87972 4808
rect 87923 4777 87935 4780
rect 87877 4771 87935 4777
rect 87966 4768 87972 4780
rect 88024 4768 88030 4820
rect 36722 4700 36728 4752
rect 36780 4740 36786 4752
rect 37185 4743 37243 4749
rect 37185 4740 37197 4743
rect 36780 4712 37197 4740
rect 36780 4700 36786 4712
rect 37185 4709 37197 4712
rect 37231 4740 37243 4743
rect 37458 4740 37464 4752
rect 37231 4712 37464 4740
rect 37231 4709 37243 4712
rect 37185 4703 37243 4709
rect 37458 4700 37464 4712
rect 37516 4740 37522 4752
rect 38470 4740 38476 4752
rect 37516 4712 38476 4740
rect 37516 4700 37522 4712
rect 37918 4632 37924 4684
rect 37976 4672 37982 4684
rect 38013 4675 38071 4681
rect 38013 4672 38025 4675
rect 37976 4644 38025 4672
rect 37976 4632 37982 4644
rect 38013 4641 38025 4644
rect 38059 4672 38071 4675
rect 38102 4672 38108 4684
rect 38059 4644 38108 4672
rect 38059 4641 38071 4644
rect 38013 4635 38071 4641
rect 38102 4632 38108 4644
rect 38160 4632 38166 4684
rect 38396 4681 38424 4712
rect 38470 4700 38476 4712
rect 38528 4700 38534 4752
rect 49878 4740 49884 4752
rect 49839 4712 49884 4740
rect 49878 4700 49884 4712
rect 49936 4700 49942 4752
rect 88607 4743 88665 4749
rect 88607 4709 88619 4743
rect 88653 4740 88665 4743
rect 88702 4740 88708 4752
rect 88653 4712 88708 4740
rect 88653 4709 88665 4712
rect 88607 4703 88665 4709
rect 88702 4700 88708 4712
rect 88760 4700 88766 4752
rect 38381 4675 38439 4681
rect 38381 4641 38393 4675
rect 38427 4641 38439 4675
rect 38562 4672 38568 4684
rect 38523 4644 38568 4672
rect 38381 4635 38439 4641
rect 38562 4632 38568 4644
rect 38620 4632 38626 4684
rect 39117 4675 39175 4681
rect 39117 4641 39129 4675
rect 39163 4641 39175 4675
rect 49970 4672 49976 4684
rect 49931 4644 49976 4672
rect 39117 4635 39175 4641
rect 35253 4607 35311 4613
rect 35253 4573 35265 4607
rect 35299 4604 35311 4607
rect 35710 4604 35716 4616
rect 35299 4576 35716 4604
rect 35299 4573 35311 4576
rect 35253 4567 35311 4573
rect 35710 4564 35716 4576
rect 35768 4564 35774 4616
rect 39132 4604 39160 4635
rect 49970 4632 49976 4644
rect 50028 4632 50034 4684
rect 63586 4632 63592 4684
rect 63644 4672 63650 4684
rect 65797 4675 65855 4681
rect 65797 4672 65809 4675
rect 63644 4644 65809 4672
rect 63644 4632 63650 4644
rect 65797 4641 65809 4644
rect 65843 4672 65855 4675
rect 66162 4672 66168 4684
rect 65843 4644 66168 4672
rect 65843 4641 65855 4644
rect 65797 4635 65855 4641
rect 66162 4632 66168 4644
rect 66220 4632 66226 4684
rect 78122 4632 78128 4684
rect 78180 4672 78186 4684
rect 78861 4675 78919 4681
rect 78861 4672 78873 4675
rect 78180 4644 78873 4672
rect 78180 4632 78186 4644
rect 78861 4641 78873 4644
rect 78907 4672 78919 4675
rect 79226 4672 79232 4684
rect 78907 4644 79232 4672
rect 78907 4641 78919 4644
rect 78861 4635 78919 4641
rect 79226 4632 79232 4644
rect 79284 4632 79290 4684
rect 39206 4604 39212 4616
rect 39132 4576 39212 4604
rect 39206 4564 39212 4576
rect 39264 4564 39270 4616
rect 56873 4607 56931 4613
rect 56873 4573 56885 4607
rect 56919 4604 56931 4607
rect 57606 4604 57612 4616
rect 56919 4576 57612 4604
rect 56919 4573 56931 4576
rect 56873 4567 56931 4573
rect 57606 4564 57612 4576
rect 57664 4564 57670 4616
rect 88245 4607 88303 4613
rect 88245 4573 88257 4607
rect 88291 4604 88303 4607
rect 88610 4604 88616 4616
rect 88291 4576 88616 4604
rect 88291 4573 88303 4576
rect 88245 4567 88303 4573
rect 88610 4564 88616 4576
rect 88668 4564 88674 4616
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 36170 4468 36176 4480
rect 36131 4440 36176 4468
rect 36170 4428 36176 4440
rect 36228 4428 36234 4480
rect 52546 4428 52552 4480
rect 52604 4468 52610 4480
rect 57793 4471 57851 4477
rect 57793 4468 57805 4471
rect 52604 4440 57805 4468
rect 52604 4428 52610 4440
rect 57793 4437 57805 4440
rect 57839 4437 57851 4471
rect 66714 4468 66720 4480
rect 66675 4440 66720 4468
rect 57793 4431 57851 4437
rect 66714 4428 66720 4440
rect 66772 4428 66778 4480
rect 79778 4468 79784 4480
rect 79739 4440 79784 4468
rect 79778 4428 79784 4440
rect 79836 4428 79842 4480
rect 89162 4468 89168 4480
rect 89123 4440 89168 4468
rect 89162 4428 89168 4440
rect 89220 4428 89226 4480
rect 1104 4378 106812 4400
rect 1104 4326 18982 4378
rect 19034 4326 19046 4378
rect 19098 4326 19110 4378
rect 19162 4326 19174 4378
rect 19226 4326 54982 4378
rect 55034 4326 55046 4378
rect 55098 4326 55110 4378
rect 55162 4326 55174 4378
rect 55226 4326 90982 4378
rect 91034 4326 91046 4378
rect 91098 4326 91110 4378
rect 91162 4326 91174 4378
rect 91226 4326 106812 4378
rect 1104 4304 106812 4326
rect 2038 4264 2044 4276
rect 1951 4236 2044 4264
rect 2038 4224 2044 4236
rect 2096 4264 2102 4276
rect 6730 4264 6736 4276
rect 2096 4236 6736 4264
rect 2096 4224 2102 4236
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 35710 4264 35716 4276
rect 35623 4236 35716 4264
rect 35710 4224 35716 4236
rect 35768 4264 35774 4276
rect 38010 4264 38016 4276
rect 35768 4236 38016 4264
rect 35768 4224 35774 4236
rect 38010 4224 38016 4236
rect 38068 4224 38074 4276
rect 38197 4267 38255 4273
rect 38197 4233 38209 4267
rect 38243 4264 38255 4267
rect 39206 4264 39212 4276
rect 38243 4236 39212 4264
rect 38243 4233 38255 4236
rect 38197 4227 38255 4233
rect 39206 4224 39212 4236
rect 39264 4224 39270 4276
rect 57606 4264 57612 4276
rect 57519 4236 57612 4264
rect 57606 4224 57612 4236
rect 57664 4264 57670 4276
rect 60918 4264 60924 4276
rect 57664 4236 60924 4264
rect 57664 4224 57670 4236
rect 60918 4224 60924 4236
rect 60976 4224 60982 4276
rect 66162 4264 66168 4276
rect 66123 4236 66168 4264
rect 66162 4224 66168 4236
rect 66220 4224 66226 4276
rect 79226 4264 79232 4276
rect 79187 4236 79232 4264
rect 79226 4224 79232 4236
rect 79284 4224 79290 4276
rect 88610 4264 88616 4276
rect 88571 4236 88616 4264
rect 88610 4224 88616 4236
rect 88668 4224 88674 4276
rect 37458 4196 37464 4208
rect 37419 4168 37464 4196
rect 37458 4156 37464 4168
rect 37516 4156 37522 4208
rect 37829 4199 37887 4205
rect 37829 4165 37841 4199
rect 37875 4196 37887 4199
rect 37918 4196 37924 4208
rect 37875 4168 37924 4196
rect 37875 4165 37887 4168
rect 37829 4159 37887 4165
rect 37918 4156 37924 4168
rect 37976 4156 37982 4208
rect 38562 4196 38568 4208
rect 38523 4168 38568 4196
rect 38562 4156 38568 4168
rect 38620 4156 38626 4208
rect 88337 4199 88395 4205
rect 88337 4165 88349 4199
rect 88383 4196 88395 4199
rect 88702 4196 88708 4208
rect 88383 4168 88708 4196
rect 88383 4165 88395 4168
rect 88337 4159 88395 4165
rect 88702 4156 88708 4168
rect 88760 4156 88766 4208
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 6914 4128 6920 4140
rect 5500 4100 6920 4128
rect 5500 4088 5506 4100
rect 6914 4088 6920 4100
rect 6972 4128 6978 4140
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6972 4100 7021 4128
rect 6972 4088 6978 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 18932 4100 20177 4128
rect 18932 4088 18938 4100
rect 20165 4097 20177 4100
rect 20211 4128 20223 4131
rect 20901 4131 20959 4137
rect 20901 4128 20913 4131
rect 20211 4100 20913 4128
rect 20211 4097 20223 4100
rect 20165 4091 20223 4097
rect 20901 4097 20913 4100
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 1394 4060 1400 4072
rect 1355 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4020 1458 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 6822 4060 6828 4072
rect 6687 4032 6828 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 12434 3924 12440 3936
rect 7515 3896 12440 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 20622 3924 20628 3936
rect 20583 3896 20628 3924
rect 20622 3884 20628 3896
rect 20680 3924 20686 3936
rect 20732 3924 20760 4023
rect 21358 3924 21364 3936
rect 20680 3896 20760 3924
rect 21319 3896 21364 3924
rect 20680 3884 20686 3896
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 35250 3924 35256 3936
rect 35211 3896 35256 3924
rect 35250 3884 35256 3896
rect 35308 3884 35314 3936
rect 49970 3924 49976 3936
rect 49931 3896 49976 3924
rect 49970 3884 49976 3896
rect 50028 3884 50034 3936
rect 56870 3924 56876 3936
rect 56831 3896 56876 3924
rect 56870 3884 56876 3896
rect 56928 3884 56934 3936
rect 65794 3924 65800 3936
rect 65755 3896 65800 3924
rect 65794 3884 65800 3896
rect 65852 3884 65858 3936
rect 78950 3924 78956 3936
rect 78911 3896 78956 3924
rect 78950 3884 78956 3896
rect 79008 3884 79014 3936
rect 1104 3834 106812 3856
rect 1104 3782 36982 3834
rect 37034 3782 37046 3834
rect 37098 3782 37110 3834
rect 37162 3782 37174 3834
rect 37226 3782 72982 3834
rect 73034 3782 73046 3834
rect 73098 3782 73110 3834
rect 73162 3782 73174 3834
rect 73226 3782 106812 3834
rect 1104 3760 106812 3782
rect 6914 3720 6920 3732
rect 6875 3692 6920 3720
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 53009 3723 53067 3729
rect 53009 3689 53021 3723
rect 53055 3720 53067 3723
rect 53926 3720 53932 3732
rect 53055 3692 53932 3720
rect 53055 3689 53067 3692
rect 53009 3683 53067 3689
rect 53926 3680 53932 3692
rect 53984 3720 53990 3732
rect 60734 3720 60740 3732
rect 53984 3692 60740 3720
rect 53984 3680 53990 3692
rect 60734 3680 60740 3692
rect 60792 3680 60798 3732
rect 36170 3544 36176 3596
rect 36228 3584 36234 3596
rect 36265 3587 36323 3593
rect 36265 3584 36277 3587
rect 36228 3556 36277 3584
rect 36228 3544 36234 3556
rect 36265 3553 36277 3556
rect 36311 3553 36323 3587
rect 52546 3584 52552 3596
rect 52507 3556 52552 3584
rect 36265 3547 36323 3553
rect 52546 3544 52552 3556
rect 52604 3544 52610 3596
rect 64417 3587 64475 3593
rect 64417 3553 64429 3587
rect 64463 3584 64475 3587
rect 64690 3584 64696 3596
rect 64463 3556 64696 3584
rect 64463 3553 64475 3556
rect 64417 3547 64475 3553
rect 64690 3544 64696 3556
rect 64748 3584 64754 3596
rect 66714 3584 66720 3596
rect 64748 3556 66720 3584
rect 64748 3544 64754 3556
rect 66714 3544 66720 3556
rect 66772 3544 66778 3596
rect 78217 3587 78275 3593
rect 78217 3553 78229 3587
rect 78263 3584 78275 3587
rect 78490 3584 78496 3596
rect 78263 3556 78496 3584
rect 78263 3553 78275 3556
rect 78217 3547 78275 3553
rect 78490 3544 78496 3556
rect 78548 3584 78554 3596
rect 79778 3584 79784 3596
rect 78548 3556 79784 3584
rect 78548 3544 78554 3556
rect 79778 3544 79784 3556
rect 79836 3544 79842 3596
rect 88245 3587 88303 3593
rect 88245 3553 88257 3587
rect 88291 3584 88303 3587
rect 88702 3584 88708 3596
rect 88291 3556 88708 3584
rect 88291 3553 88303 3556
rect 88245 3547 88303 3553
rect 88702 3544 88708 3556
rect 88760 3544 88766 3596
rect 36078 3516 36084 3528
rect 36039 3488 36084 3516
rect 36078 3476 36084 3488
rect 36136 3476 36142 3528
rect 52362 3516 52368 3528
rect 52323 3488 52368 3516
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 64230 3516 64236 3528
rect 64191 3488 64236 3516
rect 64230 3476 64236 3488
rect 64288 3476 64294 3528
rect 78030 3516 78036 3528
rect 77991 3488 78036 3516
rect 78030 3476 78036 3488
rect 78088 3476 78094 3528
rect 88429 3519 88487 3525
rect 88429 3485 88441 3519
rect 88475 3516 88487 3519
rect 89162 3516 89168 3528
rect 88475 3488 89168 3516
rect 88475 3485 88487 3488
rect 88429 3479 88487 3485
rect 89162 3476 89168 3488
rect 89220 3476 89226 3528
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1673 3383 1731 3389
rect 1673 3380 1685 3383
rect 1452 3352 1685 3380
rect 1452 3340 1458 3352
rect 1673 3349 1685 3352
rect 1719 3380 1731 3383
rect 2958 3380 2964 3392
rect 1719 3352 2964 3380
rect 1719 3349 1731 3352
rect 1673 3343 1731 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 36722 3380 36728 3392
rect 36683 3352 36728 3380
rect 36722 3340 36728 3352
rect 36780 3340 36786 3392
rect 64877 3383 64935 3389
rect 64877 3349 64889 3383
rect 64923 3380 64935 3383
rect 67450 3380 67456 3392
rect 64923 3352 67456 3380
rect 64923 3349 64935 3352
rect 64877 3343 64935 3349
rect 67450 3340 67456 3352
rect 67508 3340 67514 3392
rect 78677 3383 78735 3389
rect 78677 3349 78689 3383
rect 78723 3380 78735 3383
rect 80698 3380 80704 3392
rect 78723 3352 80704 3380
rect 78723 3349 78735 3352
rect 78677 3343 78735 3349
rect 80698 3340 80704 3352
rect 80756 3340 80762 3392
rect 88886 3380 88892 3392
rect 88847 3352 88892 3380
rect 88886 3340 88892 3352
rect 88944 3340 88950 3392
rect 1104 3290 106812 3312
rect 1104 3238 18982 3290
rect 19034 3238 19046 3290
rect 19098 3238 19110 3290
rect 19162 3238 19174 3290
rect 19226 3238 54982 3290
rect 55034 3238 55046 3290
rect 55098 3238 55110 3290
rect 55162 3238 55174 3290
rect 55226 3238 90982 3290
rect 91034 3238 91046 3290
rect 91098 3238 91110 3290
rect 91162 3238 91174 3290
rect 91226 3238 106812 3290
rect 1104 3216 106812 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 36170 3136 36176 3188
rect 36228 3176 36234 3188
rect 36449 3179 36507 3185
rect 36449 3176 36461 3179
rect 36228 3148 36461 3176
rect 36228 3136 36234 3148
rect 36449 3145 36461 3148
rect 36495 3145 36507 3179
rect 36449 3139 36507 3145
rect 52546 3136 52552 3188
rect 52604 3176 52610 3188
rect 52733 3179 52791 3185
rect 52733 3176 52745 3179
rect 52604 3148 52745 3176
rect 52604 3136 52610 3148
rect 52733 3145 52745 3148
rect 52779 3145 52791 3179
rect 64690 3176 64696 3188
rect 64651 3148 64696 3176
rect 52733 3139 52791 3145
rect 64690 3136 64696 3148
rect 64748 3136 64754 3188
rect 78490 3176 78496 3188
rect 78451 3148 78496 3176
rect 78490 3136 78496 3148
rect 78548 3136 78554 3188
rect 80698 3176 80704 3188
rect 80659 3148 80704 3176
rect 80698 3136 80704 3148
rect 80756 3136 80762 3188
rect 87969 3179 88027 3185
rect 87969 3145 87981 3179
rect 88015 3176 88027 3179
rect 88886 3176 88892 3188
rect 88015 3148 88892 3176
rect 88015 3145 88027 3148
rect 87969 3139 88027 3145
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 12434 2972 12440 2984
rect 12395 2944 12440 2972
rect 12434 2932 12440 2944
rect 12492 2972 12498 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12492 2944 13001 2972
rect 12492 2932 12498 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 21358 2932 21364 2984
rect 21416 2972 21422 2984
rect 25501 2975 25559 2981
rect 25501 2972 25513 2975
rect 21416 2944 25513 2972
rect 21416 2932 21422 2944
rect 25501 2941 25513 2944
rect 25547 2972 25559 2975
rect 26142 2972 26148 2984
rect 25547 2944 26148 2972
rect 25547 2941 25559 2944
rect 25501 2935 25559 2941
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 80057 2975 80115 2981
rect 80057 2941 80069 2975
rect 80103 2972 80115 2975
rect 80698 2972 80704 2984
rect 80103 2944 80704 2972
rect 80103 2941 80115 2944
rect 80057 2935 80115 2941
rect 80698 2932 80704 2944
rect 80756 2932 80762 2984
rect 88076 2981 88104 3148
rect 88886 3136 88892 3148
rect 88944 3136 88950 3188
rect 89073 3179 89131 3185
rect 89073 3145 89085 3179
rect 89119 3176 89131 3179
rect 89162 3176 89168 3188
rect 89119 3148 89168 3176
rect 89119 3145 89131 3148
rect 89073 3139 89131 3145
rect 89162 3136 89168 3148
rect 89220 3136 89226 3188
rect 88061 2975 88119 2981
rect 88061 2941 88073 2975
rect 88107 2941 88119 2975
rect 88061 2935 88119 2941
rect 78030 2864 78036 2916
rect 78088 2904 78094 2916
rect 78125 2907 78183 2913
rect 78125 2904 78137 2907
rect 78088 2876 78137 2904
rect 78088 2864 78094 2876
rect 78125 2873 78137 2876
rect 78171 2904 78183 2907
rect 84378 2904 84384 2916
rect 78171 2876 84384 2904
rect 78171 2873 78183 2876
rect 78125 2867 78183 2873
rect 84378 2864 84384 2876
rect 84436 2864 84442 2916
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 12618 2836 12624 2848
rect 12579 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 25682 2836 25688 2848
rect 25643 2808 25688 2836
rect 25682 2796 25688 2808
rect 25740 2796 25746 2848
rect 26142 2836 26148 2848
rect 26103 2808 26148 2836
rect 26142 2796 26148 2808
rect 26200 2796 26206 2848
rect 36170 2836 36176 2848
rect 36131 2808 36176 2836
rect 36170 2796 36176 2808
rect 36228 2796 36234 2848
rect 52362 2796 52368 2848
rect 52420 2836 52426 2848
rect 52457 2839 52515 2845
rect 52457 2836 52469 2839
rect 52420 2808 52469 2836
rect 52420 2796 52426 2808
rect 52457 2805 52469 2808
rect 52503 2836 52515 2839
rect 57054 2836 57060 2848
rect 52503 2808 57060 2836
rect 52503 2805 52515 2808
rect 52457 2799 52515 2805
rect 57054 2796 57060 2808
rect 57112 2796 57118 2848
rect 64230 2796 64236 2848
rect 64288 2836 64294 2848
rect 64325 2839 64383 2845
rect 64325 2836 64337 2839
rect 64288 2808 64337 2836
rect 64288 2796 64294 2808
rect 64325 2805 64337 2808
rect 64371 2836 64383 2839
rect 70486 2836 70492 2848
rect 64371 2808 70492 2836
rect 64371 2805 64383 2808
rect 64325 2799 64383 2805
rect 70486 2796 70492 2808
rect 70544 2796 70550 2848
rect 80238 2836 80244 2848
rect 80199 2808 80244 2836
rect 80238 2796 80244 2808
rect 80296 2796 80302 2848
rect 88242 2836 88248 2848
rect 88203 2808 88248 2836
rect 88242 2796 88248 2808
rect 88300 2796 88306 2848
rect 88702 2836 88708 2848
rect 88663 2808 88708 2836
rect 88702 2796 88708 2808
rect 88760 2796 88766 2848
rect 1104 2746 106812 2768
rect 1104 2694 36982 2746
rect 37034 2694 37046 2746
rect 37098 2694 37110 2746
rect 37162 2694 37174 2746
rect 37226 2694 72982 2746
rect 73034 2694 73046 2746
rect 73098 2694 73110 2746
rect 73162 2694 73174 2746
rect 73226 2694 106812 2746
rect 1104 2672 106812 2694
rect 46934 2632 46940 2644
rect 39868 2604 46940 2632
rect 36722 2456 36728 2508
rect 36780 2496 36786 2508
rect 39868 2505 39896 2604
rect 46934 2592 46940 2604
rect 46992 2592 46998 2644
rect 53926 2632 53932 2644
rect 53887 2604 53932 2632
rect 53926 2592 53932 2604
rect 53984 2592 53990 2644
rect 66993 2635 67051 2641
rect 66993 2601 67005 2635
rect 67039 2632 67051 2635
rect 67358 2632 67364 2644
rect 67039 2604 67364 2632
rect 67039 2601 67051 2604
rect 66993 2595 67051 2601
rect 67358 2592 67364 2604
rect 67416 2592 67422 2644
rect 67450 2592 67456 2644
rect 67508 2632 67514 2644
rect 67508 2604 67553 2632
rect 67508 2592 67514 2604
rect 39301 2499 39359 2505
rect 39301 2496 39313 2499
rect 36780 2468 39313 2496
rect 36780 2456 36786 2468
rect 39301 2465 39313 2468
rect 39347 2496 39359 2499
rect 39853 2499 39911 2505
rect 39853 2496 39865 2499
rect 39347 2468 39865 2496
rect 39347 2465 39359 2468
rect 39301 2459 39359 2465
rect 39853 2465 39865 2468
rect 39899 2465 39911 2499
rect 39853 2459 39911 2465
rect 53285 2499 53343 2505
rect 53285 2465 53297 2499
rect 53331 2496 53343 2499
rect 53944 2496 53972 2592
rect 53331 2468 53972 2496
rect 66809 2499 66867 2505
rect 53331 2465 53343 2468
rect 53285 2459 53343 2465
rect 66809 2465 66821 2499
rect 66855 2496 66867 2499
rect 67468 2496 67496 2592
rect 66855 2468 67496 2496
rect 66855 2465 66867 2468
rect 66809 2459 66867 2465
rect 39482 2292 39488 2304
rect 39443 2264 39488 2292
rect 39482 2252 39488 2264
rect 39540 2252 39546 2304
rect 53466 2292 53472 2304
rect 53427 2264 53472 2292
rect 53466 2252 53472 2264
rect 53524 2252 53530 2304
rect 1104 2202 106812 2224
rect 1104 2150 18982 2202
rect 19034 2150 19046 2202
rect 19098 2150 19110 2202
rect 19162 2150 19174 2202
rect 19226 2150 54982 2202
rect 55034 2150 55046 2202
rect 55098 2150 55110 2202
rect 55162 2150 55174 2202
rect 55226 2150 90982 2202
rect 91034 2150 91046 2202
rect 91098 2150 91110 2202
rect 91162 2150 91174 2202
rect 91226 2150 106812 2202
rect 1104 2128 106812 2150
<< via1 >>
rect 19340 13472 19392 13524
rect 20168 13472 20220 13524
rect 33140 13472 33192 13524
rect 33692 13472 33744 13524
rect 86960 13472 87012 13524
rect 87696 13472 87748 13524
rect 36982 11398 37034 11450
rect 37046 11398 37098 11450
rect 37110 11398 37162 11450
rect 37174 11398 37226 11450
rect 72982 11398 73034 11450
rect 73046 11398 73098 11450
rect 73110 11398 73162 11450
rect 73174 11398 73226 11450
rect 18982 10854 19034 10906
rect 19046 10854 19098 10906
rect 19110 10854 19162 10906
rect 19174 10854 19226 10906
rect 54982 10854 55034 10906
rect 55046 10854 55098 10906
rect 55110 10854 55162 10906
rect 55174 10854 55226 10906
rect 90982 10854 91034 10906
rect 91046 10854 91098 10906
rect 91110 10854 91162 10906
rect 91174 10854 91226 10906
rect 36982 10310 37034 10362
rect 37046 10310 37098 10362
rect 37110 10310 37162 10362
rect 37174 10310 37226 10362
rect 72982 10310 73034 10362
rect 73046 10310 73098 10362
rect 73110 10310 73162 10362
rect 73174 10310 73226 10362
rect 18982 9766 19034 9818
rect 19046 9766 19098 9818
rect 19110 9766 19162 9818
rect 19174 9766 19226 9818
rect 54982 9766 55034 9818
rect 55046 9766 55098 9818
rect 55110 9766 55162 9818
rect 55174 9766 55226 9818
rect 90982 9766 91034 9818
rect 91046 9766 91098 9818
rect 91110 9766 91162 9818
rect 91174 9766 91226 9818
rect 73344 9324 73396 9376
rect 74172 9324 74224 9376
rect 36982 9222 37034 9274
rect 37046 9222 37098 9274
rect 37110 9222 37162 9274
rect 37174 9222 37226 9274
rect 72982 9222 73034 9274
rect 73046 9222 73098 9274
rect 73110 9222 73162 9274
rect 73174 9222 73226 9274
rect 18982 8678 19034 8730
rect 19046 8678 19098 8730
rect 19110 8678 19162 8730
rect 19174 8678 19226 8730
rect 54982 8678 55034 8730
rect 55046 8678 55098 8730
rect 55110 8678 55162 8730
rect 55174 8678 55226 8730
rect 90982 8678 91034 8730
rect 91046 8678 91098 8730
rect 91110 8678 91162 8730
rect 91174 8678 91226 8730
rect 36982 8134 37034 8186
rect 37046 8134 37098 8186
rect 37110 8134 37162 8186
rect 37174 8134 37226 8186
rect 72982 8134 73034 8186
rect 73046 8134 73098 8186
rect 73110 8134 73162 8186
rect 73174 8134 73226 8186
rect 18982 7590 19034 7642
rect 19046 7590 19098 7642
rect 19110 7590 19162 7642
rect 19174 7590 19226 7642
rect 54982 7590 55034 7642
rect 55046 7590 55098 7642
rect 55110 7590 55162 7642
rect 55174 7590 55226 7642
rect 90982 7590 91034 7642
rect 91046 7590 91098 7642
rect 91110 7590 91162 7642
rect 91174 7590 91226 7642
rect 36982 7046 37034 7098
rect 37046 7046 37098 7098
rect 37110 7046 37162 7098
rect 37174 7046 37226 7098
rect 72982 7046 73034 7098
rect 73046 7046 73098 7098
rect 73110 7046 73162 7098
rect 73174 7046 73226 7098
rect 37924 6647 37976 6656
rect 37924 6613 37933 6647
rect 37933 6613 37967 6647
rect 37967 6613 37976 6647
rect 37924 6604 37976 6613
rect 18982 6502 19034 6554
rect 19046 6502 19098 6554
rect 19110 6502 19162 6554
rect 19174 6502 19226 6554
rect 54982 6502 55034 6554
rect 55046 6502 55098 6554
rect 55110 6502 55162 6554
rect 55174 6502 55226 6554
rect 90982 6502 91034 6554
rect 91046 6502 91098 6554
rect 91110 6502 91162 6554
rect 91174 6502 91226 6554
rect 37924 6196 37976 6248
rect 38384 6196 38436 6248
rect 38568 6239 38620 6248
rect 38568 6205 38577 6239
rect 38577 6205 38611 6239
rect 38611 6205 38620 6239
rect 38568 6196 38620 6205
rect 39212 6196 39264 6248
rect 63132 6196 63184 6248
rect 77760 6239 77812 6248
rect 77760 6205 77769 6239
rect 77769 6205 77803 6239
rect 77803 6205 77812 6239
rect 77760 6196 77812 6205
rect 36728 6103 36780 6112
rect 36728 6069 36737 6103
rect 36737 6069 36771 6103
rect 36771 6069 36780 6103
rect 36728 6060 36780 6069
rect 37648 6103 37700 6112
rect 37648 6069 37657 6103
rect 37657 6069 37691 6103
rect 37691 6069 37700 6103
rect 37648 6060 37700 6069
rect 77484 6103 77536 6112
rect 77484 6069 77493 6103
rect 77493 6069 77527 6103
rect 77527 6069 77536 6103
rect 77484 6060 77536 6069
rect 36982 5958 37034 6010
rect 37046 5958 37098 6010
rect 37110 5958 37162 6010
rect 37174 5958 37226 6010
rect 72982 5958 73034 6010
rect 73046 5958 73098 6010
rect 73110 5958 73162 6010
rect 73174 5958 73226 6010
rect 37832 5899 37884 5908
rect 37832 5865 37841 5899
rect 37841 5865 37875 5899
rect 37875 5865 37884 5899
rect 37832 5856 37884 5865
rect 38108 5856 38160 5908
rect 60280 5856 60332 5908
rect 63132 5899 63184 5908
rect 63132 5865 63141 5899
rect 63141 5865 63175 5899
rect 63175 5865 63184 5899
rect 63132 5856 63184 5865
rect 77484 5899 77536 5908
rect 77484 5865 77493 5899
rect 77493 5865 77527 5899
rect 77527 5865 77536 5899
rect 77484 5856 77536 5865
rect 51816 5831 51868 5840
rect 51816 5797 51825 5831
rect 51825 5797 51859 5831
rect 51859 5797 51868 5831
rect 51816 5788 51868 5797
rect 59820 5788 59872 5840
rect 62856 5788 62908 5840
rect 38384 5763 38436 5772
rect 38384 5729 38393 5763
rect 38393 5729 38427 5763
rect 38427 5729 38436 5763
rect 38384 5720 38436 5729
rect 38568 5763 38620 5772
rect 38568 5729 38577 5763
rect 38577 5729 38611 5763
rect 38611 5729 38620 5763
rect 38568 5720 38620 5729
rect 39120 5763 39172 5772
rect 39120 5729 39129 5763
rect 39129 5729 39163 5763
rect 39163 5729 39172 5763
rect 39120 5720 39172 5729
rect 60372 5763 60424 5772
rect 37556 5695 37608 5704
rect 37556 5661 37565 5695
rect 37565 5661 37599 5695
rect 37599 5661 37608 5695
rect 37556 5652 37608 5661
rect 51172 5652 51224 5704
rect 60372 5729 60381 5763
rect 60381 5729 60415 5763
rect 60415 5729 60424 5763
rect 60372 5720 60424 5729
rect 62764 5720 62816 5772
rect 68836 5763 68888 5772
rect 68836 5729 68845 5763
rect 68845 5729 68879 5763
rect 68879 5729 68888 5763
rect 68836 5720 68888 5729
rect 60188 5695 60240 5704
rect 60188 5661 60197 5695
rect 60197 5661 60231 5695
rect 60231 5661 60240 5695
rect 60188 5652 60240 5661
rect 60924 5695 60976 5704
rect 60924 5661 60933 5695
rect 60933 5661 60967 5695
rect 60967 5661 60976 5695
rect 60924 5652 60976 5661
rect 63224 5652 63276 5704
rect 63592 5695 63644 5704
rect 63592 5661 63601 5695
rect 63601 5661 63635 5695
rect 63635 5661 63644 5695
rect 63592 5652 63644 5661
rect 68744 5695 68796 5704
rect 68744 5661 68753 5695
rect 68753 5661 68787 5695
rect 68787 5661 68796 5695
rect 68744 5652 68796 5661
rect 88156 5516 88208 5568
rect 18982 5414 19034 5466
rect 19046 5414 19098 5466
rect 19110 5414 19162 5466
rect 19174 5414 19226 5466
rect 54982 5414 55034 5466
rect 55046 5414 55098 5466
rect 55110 5414 55162 5466
rect 55174 5414 55226 5466
rect 90982 5414 91034 5466
rect 91046 5414 91098 5466
rect 91110 5414 91162 5466
rect 91174 5414 91226 5466
rect 38108 5312 38160 5364
rect 39764 5355 39816 5364
rect 39764 5321 39773 5355
rect 39773 5321 39807 5355
rect 39807 5321 39816 5355
rect 39764 5312 39816 5321
rect 59820 5355 59872 5364
rect 59820 5321 59829 5355
rect 59829 5321 59863 5355
rect 59863 5321 59872 5355
rect 59820 5312 59872 5321
rect 60188 5312 60240 5364
rect 61016 5312 61068 5364
rect 63132 5312 63184 5364
rect 68744 5312 68796 5364
rect 60280 5287 60332 5296
rect 60280 5253 60289 5287
rect 60289 5253 60323 5287
rect 60323 5253 60332 5287
rect 60280 5244 60332 5253
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 37924 5176 37976 5228
rect 2320 5108 2372 5160
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 39764 5176 39816 5228
rect 51172 5219 51224 5228
rect 51172 5185 51181 5219
rect 51181 5185 51215 5219
rect 51215 5185 51224 5219
rect 51172 5176 51224 5185
rect 62764 5219 62816 5228
rect 38476 5151 38528 5160
rect 38476 5117 38485 5151
rect 38485 5117 38519 5151
rect 38519 5117 38528 5151
rect 38476 5108 38528 5117
rect 38568 5108 38620 5160
rect 39120 5151 39172 5160
rect 39120 5117 39129 5151
rect 39129 5117 39163 5151
rect 39163 5117 39172 5151
rect 39120 5108 39172 5117
rect 62764 5185 62773 5219
rect 62773 5185 62807 5219
rect 62807 5185 62816 5219
rect 62764 5176 62816 5185
rect 77484 5176 77536 5228
rect 79416 5176 79468 5228
rect 1676 4972 1728 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18880 4972 18932 5024
rect 36728 5015 36780 5024
rect 36728 4981 36737 5015
rect 36737 4981 36771 5015
rect 36771 4981 36780 5015
rect 36728 4972 36780 4981
rect 38016 5015 38068 5024
rect 38016 4981 38025 5015
rect 38025 4981 38059 5015
rect 38059 4981 38068 5015
rect 38016 4972 38068 4981
rect 60372 4972 60424 5024
rect 77852 5108 77904 5160
rect 88064 5151 88116 5160
rect 88064 5117 88073 5151
rect 88073 5117 88107 5151
rect 88107 5117 88116 5151
rect 88064 5108 88116 5117
rect 63224 5083 63276 5092
rect 63224 5049 63233 5083
rect 63233 5049 63267 5083
rect 63267 5049 63276 5083
rect 63224 5040 63276 5049
rect 72792 5040 72844 5092
rect 68836 5015 68888 5024
rect 68836 4981 68845 5015
rect 68845 4981 68879 5015
rect 68879 4981 68888 5015
rect 68836 4972 68888 4981
rect 77484 5040 77536 5092
rect 78128 5083 78180 5092
rect 78128 5049 78137 5083
rect 78137 5049 78171 5083
rect 78171 5049 78180 5083
rect 78128 5040 78180 5049
rect 87144 5040 87196 5092
rect 79416 4972 79468 5024
rect 88156 5083 88208 5092
rect 88156 5049 88165 5083
rect 88165 5049 88199 5083
rect 88199 5049 88208 5083
rect 88156 5040 88208 5049
rect 88616 5040 88668 5092
rect 87972 5015 88024 5024
rect 87972 4981 87981 5015
rect 87981 4981 88015 5015
rect 88015 4981 88024 5015
rect 87972 4972 88024 4981
rect 36982 4870 37034 4922
rect 37046 4870 37098 4922
rect 37110 4870 37162 4922
rect 37174 4870 37226 4922
rect 72982 4870 73034 4922
rect 73046 4870 73098 4922
rect 73110 4870 73162 4922
rect 73174 4870 73226 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 35256 4768 35308 4820
rect 37556 4811 37608 4820
rect 37556 4777 37565 4811
rect 37565 4777 37599 4811
rect 37599 4777 37608 4811
rect 37556 4768 37608 4777
rect 37832 4811 37884 4820
rect 37832 4777 37841 4811
rect 37841 4777 37875 4811
rect 37875 4777 37884 4811
rect 37832 4768 37884 4777
rect 56876 4768 56928 4820
rect 62856 4811 62908 4820
rect 62856 4777 62865 4811
rect 62865 4777 62899 4811
rect 62899 4777 62908 4811
rect 62856 4768 62908 4777
rect 65800 4768 65852 4820
rect 77392 4811 77444 4820
rect 77392 4777 77401 4811
rect 77401 4777 77435 4811
rect 77435 4777 77444 4811
rect 77392 4768 77444 4777
rect 78956 4768 79008 4820
rect 87144 4768 87196 4820
rect 87972 4768 88024 4820
rect 36728 4700 36780 4752
rect 37464 4700 37516 4752
rect 37924 4632 37976 4684
rect 38108 4632 38160 4684
rect 38476 4700 38528 4752
rect 49884 4743 49936 4752
rect 49884 4709 49893 4743
rect 49893 4709 49927 4743
rect 49927 4709 49936 4743
rect 49884 4700 49936 4709
rect 88708 4700 88760 4752
rect 38568 4675 38620 4684
rect 38568 4641 38577 4675
rect 38577 4641 38611 4675
rect 38611 4641 38620 4675
rect 38568 4632 38620 4641
rect 49976 4675 50028 4684
rect 35716 4564 35768 4616
rect 49976 4641 49985 4675
rect 49985 4641 50019 4675
rect 50019 4641 50028 4675
rect 49976 4632 50028 4641
rect 63592 4632 63644 4684
rect 66168 4632 66220 4684
rect 78128 4632 78180 4684
rect 79232 4632 79284 4684
rect 39212 4564 39264 4616
rect 57612 4564 57664 4616
rect 88616 4564 88668 4616
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 36176 4471 36228 4480
rect 36176 4437 36185 4471
rect 36185 4437 36219 4471
rect 36219 4437 36228 4471
rect 36176 4428 36228 4437
rect 52552 4428 52604 4480
rect 66720 4471 66772 4480
rect 66720 4437 66729 4471
rect 66729 4437 66763 4471
rect 66763 4437 66772 4471
rect 66720 4428 66772 4437
rect 79784 4471 79836 4480
rect 79784 4437 79793 4471
rect 79793 4437 79827 4471
rect 79827 4437 79836 4471
rect 79784 4428 79836 4437
rect 89168 4471 89220 4480
rect 89168 4437 89177 4471
rect 89177 4437 89211 4471
rect 89211 4437 89220 4471
rect 89168 4428 89220 4437
rect 18982 4326 19034 4378
rect 19046 4326 19098 4378
rect 19110 4326 19162 4378
rect 19174 4326 19226 4378
rect 54982 4326 55034 4378
rect 55046 4326 55098 4378
rect 55110 4326 55162 4378
rect 55174 4326 55226 4378
rect 90982 4326 91034 4378
rect 91046 4326 91098 4378
rect 91110 4326 91162 4378
rect 91174 4326 91226 4378
rect 2044 4267 2096 4276
rect 2044 4233 2053 4267
rect 2053 4233 2087 4267
rect 2087 4233 2096 4267
rect 2044 4224 2096 4233
rect 6736 4224 6788 4276
rect 35716 4267 35768 4276
rect 35716 4233 35725 4267
rect 35725 4233 35759 4267
rect 35759 4233 35768 4267
rect 35716 4224 35768 4233
rect 38016 4224 38068 4276
rect 39212 4224 39264 4276
rect 57612 4267 57664 4276
rect 57612 4233 57621 4267
rect 57621 4233 57655 4267
rect 57655 4233 57664 4267
rect 57612 4224 57664 4233
rect 60924 4224 60976 4276
rect 66168 4267 66220 4276
rect 66168 4233 66177 4267
rect 66177 4233 66211 4267
rect 66211 4233 66220 4267
rect 66168 4224 66220 4233
rect 79232 4267 79284 4276
rect 79232 4233 79241 4267
rect 79241 4233 79275 4267
rect 79275 4233 79284 4267
rect 79232 4224 79284 4233
rect 88616 4267 88668 4276
rect 88616 4233 88625 4267
rect 88625 4233 88659 4267
rect 88659 4233 88668 4267
rect 88616 4224 88668 4233
rect 37464 4199 37516 4208
rect 37464 4165 37473 4199
rect 37473 4165 37507 4199
rect 37507 4165 37516 4199
rect 37464 4156 37516 4165
rect 37924 4156 37976 4208
rect 38568 4199 38620 4208
rect 38568 4165 38577 4199
rect 38577 4165 38611 4199
rect 38611 4165 38620 4199
rect 38568 4156 38620 4165
rect 88708 4156 88760 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 5448 4088 5500 4140
rect 6920 4088 6972 4140
rect 18880 4088 18932 4140
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 12440 3884 12492 3936
rect 20628 3927 20680 3936
rect 20628 3893 20637 3927
rect 20637 3893 20671 3927
rect 20671 3893 20680 3927
rect 21364 3927 21416 3936
rect 20628 3884 20680 3893
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 35256 3927 35308 3936
rect 35256 3893 35265 3927
rect 35265 3893 35299 3927
rect 35299 3893 35308 3927
rect 35256 3884 35308 3893
rect 49976 3927 50028 3936
rect 49976 3893 49985 3927
rect 49985 3893 50019 3927
rect 50019 3893 50028 3927
rect 49976 3884 50028 3893
rect 56876 3927 56928 3936
rect 56876 3893 56885 3927
rect 56885 3893 56919 3927
rect 56919 3893 56928 3927
rect 56876 3884 56928 3893
rect 65800 3927 65852 3936
rect 65800 3893 65809 3927
rect 65809 3893 65843 3927
rect 65843 3893 65852 3927
rect 65800 3884 65852 3893
rect 78956 3927 79008 3936
rect 78956 3893 78965 3927
rect 78965 3893 78999 3927
rect 78999 3893 79008 3927
rect 78956 3884 79008 3893
rect 36982 3782 37034 3834
rect 37046 3782 37098 3834
rect 37110 3782 37162 3834
rect 37174 3782 37226 3834
rect 72982 3782 73034 3834
rect 73046 3782 73098 3834
rect 73110 3782 73162 3834
rect 73174 3782 73226 3834
rect 6920 3723 6972 3732
rect 6920 3689 6929 3723
rect 6929 3689 6963 3723
rect 6963 3689 6972 3723
rect 6920 3680 6972 3689
rect 53932 3680 53984 3732
rect 60740 3680 60792 3732
rect 36176 3544 36228 3596
rect 52552 3587 52604 3596
rect 52552 3553 52561 3587
rect 52561 3553 52595 3587
rect 52595 3553 52604 3587
rect 52552 3544 52604 3553
rect 64696 3544 64748 3596
rect 66720 3544 66772 3596
rect 78496 3544 78548 3596
rect 79784 3544 79836 3596
rect 88708 3544 88760 3596
rect 36084 3519 36136 3528
rect 36084 3485 36093 3519
rect 36093 3485 36127 3519
rect 36127 3485 36136 3519
rect 36084 3476 36136 3485
rect 52368 3519 52420 3528
rect 52368 3485 52377 3519
rect 52377 3485 52411 3519
rect 52411 3485 52420 3519
rect 52368 3476 52420 3485
rect 64236 3519 64288 3528
rect 64236 3485 64245 3519
rect 64245 3485 64279 3519
rect 64279 3485 64288 3519
rect 64236 3476 64288 3485
rect 78036 3519 78088 3528
rect 78036 3485 78045 3519
rect 78045 3485 78079 3519
rect 78079 3485 78088 3519
rect 78036 3476 78088 3485
rect 89168 3476 89220 3528
rect 1400 3340 1452 3392
rect 2964 3340 3016 3392
rect 36728 3383 36780 3392
rect 36728 3349 36737 3383
rect 36737 3349 36771 3383
rect 36771 3349 36780 3383
rect 36728 3340 36780 3349
rect 67456 3340 67508 3392
rect 80704 3340 80756 3392
rect 88892 3383 88944 3392
rect 88892 3349 88901 3383
rect 88901 3349 88935 3383
rect 88935 3349 88944 3383
rect 88892 3340 88944 3349
rect 18982 3238 19034 3290
rect 19046 3238 19098 3290
rect 19110 3238 19162 3290
rect 19174 3238 19226 3290
rect 54982 3238 55034 3290
rect 55046 3238 55098 3290
rect 55110 3238 55162 3290
rect 55174 3238 55226 3290
rect 90982 3238 91034 3290
rect 91046 3238 91098 3290
rect 91110 3238 91162 3290
rect 91174 3238 91226 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 36176 3136 36228 3188
rect 52552 3136 52604 3188
rect 64696 3179 64748 3188
rect 64696 3145 64705 3179
rect 64705 3145 64739 3179
rect 64739 3145 64748 3179
rect 64696 3136 64748 3145
rect 78496 3179 78548 3188
rect 78496 3145 78505 3179
rect 78505 3145 78539 3179
rect 78539 3145 78548 3179
rect 78496 3136 78548 3145
rect 80704 3179 80756 3188
rect 80704 3145 80713 3179
rect 80713 3145 80747 3179
rect 80747 3145 80756 3179
rect 80704 3136 80756 3145
rect 2044 2932 2096 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 21364 2932 21416 2984
rect 26148 2932 26200 2984
rect 80704 2932 80756 2984
rect 88892 3136 88944 3188
rect 89168 3136 89220 3188
rect 78036 2864 78088 2916
rect 84384 2864 84436 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 25688 2839 25740 2848
rect 25688 2805 25697 2839
rect 25697 2805 25731 2839
rect 25731 2805 25740 2839
rect 25688 2796 25740 2805
rect 26148 2839 26200 2848
rect 26148 2805 26157 2839
rect 26157 2805 26191 2839
rect 26191 2805 26200 2839
rect 26148 2796 26200 2805
rect 36176 2839 36228 2848
rect 36176 2805 36185 2839
rect 36185 2805 36219 2839
rect 36219 2805 36228 2839
rect 36176 2796 36228 2805
rect 52368 2796 52420 2848
rect 57060 2796 57112 2848
rect 64236 2796 64288 2848
rect 70492 2796 70544 2848
rect 80244 2839 80296 2848
rect 80244 2805 80253 2839
rect 80253 2805 80287 2839
rect 80287 2805 80296 2839
rect 80244 2796 80296 2805
rect 88248 2839 88300 2848
rect 88248 2805 88257 2839
rect 88257 2805 88291 2839
rect 88291 2805 88300 2839
rect 88248 2796 88300 2805
rect 88708 2839 88760 2848
rect 88708 2805 88717 2839
rect 88717 2805 88751 2839
rect 88751 2805 88760 2839
rect 88708 2796 88760 2805
rect 36982 2694 37034 2746
rect 37046 2694 37098 2746
rect 37110 2694 37162 2746
rect 37174 2694 37226 2746
rect 72982 2694 73034 2746
rect 73046 2694 73098 2746
rect 73110 2694 73162 2746
rect 73174 2694 73226 2746
rect 36728 2456 36780 2508
rect 46940 2592 46992 2644
rect 53932 2635 53984 2644
rect 53932 2601 53941 2635
rect 53941 2601 53975 2635
rect 53975 2601 53984 2635
rect 53932 2592 53984 2601
rect 67364 2592 67416 2644
rect 67456 2635 67508 2644
rect 67456 2601 67465 2635
rect 67465 2601 67499 2635
rect 67499 2601 67508 2635
rect 67456 2592 67508 2601
rect 39488 2295 39540 2304
rect 39488 2261 39497 2295
rect 39497 2261 39531 2295
rect 39531 2261 39540 2295
rect 39488 2252 39540 2261
rect 53472 2295 53524 2304
rect 53472 2261 53481 2295
rect 53481 2261 53515 2295
rect 53515 2261 53524 2295
rect 53472 2252 53524 2261
rect 18982 2150 19034 2202
rect 19046 2150 19098 2202
rect 19110 2150 19162 2202
rect 19174 2150 19226 2202
rect 54982 2150 55034 2202
rect 55046 2150 55098 2202
rect 55110 2150 55162 2202
rect 55174 2150 55226 2202
rect 90982 2150 91034 2202
rect 91046 2150 91098 2202
rect 91110 2150 91162 2202
rect 91174 2150 91226 2202
<< metal2 >>
rect 6734 13520 6790 14000
rect 19340 13524 19392 13530
rect 4526 5264 4582 5273
rect 4526 5199 4582 5208
rect 4540 5166 4568 5199
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4826 1716 4966
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 4154 1716 4762
rect 2332 4486 2360 5102
rect 4540 4826 4568 5102
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 1596 4146 1716 4154
rect 1584 4140 1716 4146
rect 1636 4126 1716 4140
rect 1584 4082 1636 4088
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1412 3398 1440 4014
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 2056 3194 2084 4218
rect 2332 3641 2360 4422
rect 4908 3913 4936 4966
rect 5460 4146 5488 4966
rect 6748 4282 6776 13520
rect 20166 13524 20222 14000
rect 20166 13520 20168 13524
rect 19340 13466 19392 13472
rect 20220 13520 20222 13524
rect 33140 13524 33192 13530
rect 20168 13466 20220 13472
rect 33690 13524 33746 14000
rect 47214 13546 47270 14000
rect 33690 13520 33692 13524
rect 33140 13466 33192 13472
rect 33744 13520 33746 13524
rect 46952 13520 47270 13546
rect 60738 13520 60794 14000
rect 74170 13520 74226 14000
rect 86960 13524 87012 13530
rect 33692 13466 33744 13472
rect 46952 13518 47256 13520
rect 18956 10908 19252 10928
rect 19012 10906 19036 10908
rect 19092 10906 19116 10908
rect 19172 10906 19196 10908
rect 19034 10854 19036 10906
rect 19098 10854 19110 10906
rect 19172 10854 19174 10906
rect 19012 10852 19036 10854
rect 19092 10852 19116 10854
rect 19172 10852 19196 10854
rect 18956 10832 19252 10852
rect 18956 9820 19252 9840
rect 19012 9818 19036 9820
rect 19092 9818 19116 9820
rect 19172 9818 19196 9820
rect 19034 9766 19036 9818
rect 19098 9766 19110 9818
rect 19172 9766 19174 9818
rect 19012 9764 19036 9766
rect 19092 9764 19116 9766
rect 19172 9764 19196 9766
rect 18956 9744 19252 9764
rect 18956 8732 19252 8752
rect 19012 8730 19036 8732
rect 19092 8730 19116 8732
rect 19172 8730 19196 8732
rect 19034 8678 19036 8730
rect 19098 8678 19110 8730
rect 19172 8678 19174 8730
rect 19012 8676 19036 8678
rect 19092 8676 19116 8678
rect 19172 8676 19196 8678
rect 18956 8656 19252 8676
rect 18956 7644 19252 7664
rect 19012 7642 19036 7644
rect 19092 7642 19116 7644
rect 19172 7642 19196 7644
rect 19034 7590 19036 7642
rect 19098 7590 19110 7642
rect 19172 7590 19174 7642
rect 19012 7588 19036 7590
rect 19092 7588 19116 7590
rect 19172 7588 19196 7590
rect 18956 7568 19252 7588
rect 18956 6556 19252 6576
rect 19012 6554 19036 6556
rect 19092 6554 19116 6556
rect 19172 6554 19196 6556
rect 19034 6502 19036 6554
rect 19098 6502 19110 6554
rect 19172 6502 19174 6554
rect 19012 6500 19036 6502
rect 19092 6500 19116 6502
rect 19172 6500 19196 6502
rect 18956 6480 19252 6500
rect 18956 5468 19252 5488
rect 19012 5466 19036 5468
rect 19092 5466 19116 5468
rect 19172 5466 19196 5468
rect 19034 5414 19036 5466
rect 19098 5414 19110 5466
rect 19172 5414 19174 5466
rect 19012 5412 19036 5414
rect 19092 5412 19116 5414
rect 19172 5412 19196 5414
rect 18956 5392 19252 5412
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18064 5137 18092 5170
rect 18050 5128 18106 5137
rect 18050 5063 18106 5072
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 4894 3904 4950 3913
rect 4894 3839 4950 3848
rect 2318 3632 2374 3641
rect 2318 3567 2374 3576
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 1465 1624 2790
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 2976 82 3004 3334
rect 6840 2553 6868 4014
rect 6932 3738 6960 4082
rect 12438 4040 12494 4049
rect 12438 3975 12494 3984
rect 12452 3942 12480 3975
rect 12440 3936 12492 3942
rect 17788 3913 17816 4966
rect 18064 4826 18092 5063
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18892 4146 18920 4966
rect 18956 4380 19252 4400
rect 19012 4378 19036 4380
rect 19092 4378 19116 4380
rect 19172 4378 19196 4380
rect 19034 4326 19036 4378
rect 19098 4326 19110 4378
rect 19172 4326 19174 4378
rect 19012 4324 19036 4326
rect 19092 4324 19116 4326
rect 19172 4324 19196 4326
rect 18956 4304 19252 4324
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 19352 4049 19380 13466
rect 20180 13435 20208 13466
rect 19338 4040 19394 4049
rect 19338 3975 19394 3984
rect 20628 3936 20680 3942
rect 12440 3878 12492 3884
rect 17774 3904 17830 3913
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 12452 2990 12480 3878
rect 20628 3878 20680 3884
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 17774 3839 17830 3848
rect 18956 3292 19252 3312
rect 19012 3290 19036 3292
rect 19092 3290 19116 3292
rect 19172 3290 19196 3292
rect 19034 3238 19036 3290
rect 19098 3238 19110 3290
rect 19172 3238 19174 3290
rect 19012 3236 19036 3238
rect 19092 3236 19116 3238
rect 19172 3236 19196 3238
rect 18956 3216 19252 3236
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 6826 2544 6882 2553
rect 6826 2479 6882 2488
rect 12636 2417 12664 2790
rect 16854 2544 16910 2553
rect 16854 2479 16910 2488
rect 12622 2408 12678 2417
rect 12622 2343 12678 2352
rect 9770 1456 9826 1465
rect 9770 1391 9826 1400
rect 3330 82 3386 480
rect 2976 54 3386 82
rect 9784 82 9812 1391
rect 10046 82 10102 480
rect 9784 54 10102 82
rect 3330 0 3386 54
rect 10046 0 10102 54
rect 16762 82 16818 480
rect 16868 82 16896 2479
rect 18956 2204 19252 2224
rect 19012 2202 19036 2204
rect 19092 2202 19116 2204
rect 19172 2202 19196 2204
rect 19034 2150 19036 2202
rect 19098 2150 19110 2202
rect 19172 2150 19174 2202
rect 19012 2148 19036 2150
rect 19092 2148 19116 2150
rect 19172 2148 19196 2150
rect 18956 2128 19252 2148
rect 20640 1465 20668 3878
rect 21376 2990 21404 3878
rect 21364 2984 21416 2990
rect 26148 2984 26200 2990
rect 21364 2926 21416 2932
rect 26146 2952 26148 2961
rect 33152 2961 33180 13466
rect 33704 13435 33732 13466
rect 36956 11452 37252 11472
rect 37012 11450 37036 11452
rect 37092 11450 37116 11452
rect 37172 11450 37196 11452
rect 37034 11398 37036 11450
rect 37098 11398 37110 11450
rect 37172 11398 37174 11450
rect 37012 11396 37036 11398
rect 37092 11396 37116 11398
rect 37172 11396 37196 11398
rect 36956 11376 37252 11396
rect 36956 10364 37252 10384
rect 37012 10362 37036 10364
rect 37092 10362 37116 10364
rect 37172 10362 37196 10364
rect 37034 10310 37036 10362
rect 37098 10310 37110 10362
rect 37172 10310 37174 10362
rect 37012 10308 37036 10310
rect 37092 10308 37116 10310
rect 37172 10308 37196 10310
rect 36956 10288 37252 10308
rect 36956 9276 37252 9296
rect 37012 9274 37036 9276
rect 37092 9274 37116 9276
rect 37172 9274 37196 9276
rect 37034 9222 37036 9274
rect 37098 9222 37110 9274
rect 37172 9222 37174 9274
rect 37012 9220 37036 9222
rect 37092 9220 37116 9222
rect 37172 9220 37196 9222
rect 36956 9200 37252 9220
rect 36956 8188 37252 8208
rect 37012 8186 37036 8188
rect 37092 8186 37116 8188
rect 37172 8186 37196 8188
rect 37034 8134 37036 8186
rect 37098 8134 37110 8186
rect 37172 8134 37174 8186
rect 37012 8132 37036 8134
rect 37092 8132 37116 8134
rect 37172 8132 37196 8134
rect 36956 8112 37252 8132
rect 36956 7100 37252 7120
rect 37012 7098 37036 7100
rect 37092 7098 37116 7100
rect 37172 7098 37196 7100
rect 37034 7046 37036 7098
rect 37098 7046 37110 7098
rect 37172 7046 37174 7098
rect 37012 7044 37036 7046
rect 37092 7044 37116 7046
rect 37172 7044 37196 7046
rect 36956 7024 37252 7044
rect 37924 6656 37976 6662
rect 37924 6598 37976 6604
rect 37936 6254 37964 6598
rect 38566 6352 38622 6361
rect 38566 6287 38622 6296
rect 38580 6254 38608 6287
rect 37924 6248 37976 6254
rect 37924 6190 37976 6196
rect 38384 6248 38436 6254
rect 38384 6190 38436 6196
rect 38568 6248 38620 6254
rect 38568 6190 38620 6196
rect 39212 6248 39264 6254
rect 39212 6190 39264 6196
rect 36728 6112 36780 6118
rect 36728 6054 36780 6060
rect 37648 6112 37700 6118
rect 37648 6054 37700 6060
rect 36740 5030 36768 6054
rect 36956 6012 37252 6032
rect 37012 6010 37036 6012
rect 37092 6010 37116 6012
rect 37172 6010 37196 6012
rect 37034 5958 37036 6010
rect 37098 5958 37110 6010
rect 37172 5958 37174 6010
rect 37012 5956 37036 5958
rect 37092 5956 37116 5958
rect 37172 5956 37196 5958
rect 36956 5936 37252 5956
rect 37556 5704 37608 5710
rect 37556 5646 37608 5652
rect 36728 5024 36780 5030
rect 36728 4966 36780 4972
rect 35256 4820 35308 4826
rect 35256 4762 35308 4768
rect 35268 3942 35296 4762
rect 36740 4758 36768 4966
rect 36956 4924 37252 4944
rect 37012 4922 37036 4924
rect 37092 4922 37116 4924
rect 37172 4922 37196 4924
rect 37034 4870 37036 4922
rect 37098 4870 37110 4922
rect 37172 4870 37174 4922
rect 37012 4868 37036 4870
rect 37092 4868 37116 4870
rect 37172 4868 37196 4870
rect 36956 4848 37252 4868
rect 37568 4826 37596 5646
rect 37660 5273 37688 6054
rect 37832 5908 37884 5914
rect 37832 5850 37884 5856
rect 37646 5264 37702 5273
rect 37646 5199 37702 5208
rect 37844 5137 37872 5850
rect 37936 5234 37964 6190
rect 38108 5908 38160 5914
rect 38108 5850 38160 5856
rect 38120 5817 38148 5850
rect 38106 5808 38162 5817
rect 38396 5778 38424 6190
rect 38580 5778 38608 6190
rect 38106 5743 38162 5752
rect 38384 5772 38436 5778
rect 38120 5370 38148 5743
rect 38568 5772 38620 5778
rect 38436 5732 38516 5760
rect 38384 5714 38436 5720
rect 38108 5364 38160 5370
rect 38108 5306 38160 5312
rect 37924 5228 37976 5234
rect 37924 5170 37976 5176
rect 37830 5128 37886 5137
rect 37830 5063 37886 5072
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 37556 4820 37608 4826
rect 37556 4762 37608 4768
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 36728 4752 36780 4758
rect 36728 4694 36780 4700
rect 37464 4752 37516 4758
rect 37464 4694 37516 4700
rect 35716 4616 35768 4622
rect 35716 4558 35768 4564
rect 35728 4282 35756 4558
rect 36176 4480 36228 4486
rect 36176 4422 36228 4428
rect 35716 4276 35768 4282
rect 35716 4218 35768 4224
rect 35256 3936 35308 3942
rect 35254 3904 35256 3913
rect 35308 3904 35310 3913
rect 35254 3839 35310 3848
rect 35268 3097 35296 3839
rect 36188 3602 36216 4422
rect 37476 4214 37504 4694
rect 37464 4208 37516 4214
rect 37464 4150 37516 4156
rect 36956 3836 37252 3856
rect 37012 3834 37036 3836
rect 37092 3834 37116 3836
rect 37172 3834 37196 3836
rect 37034 3782 37036 3834
rect 37098 3782 37110 3834
rect 37172 3782 37174 3834
rect 37012 3780 37036 3782
rect 37092 3780 37116 3782
rect 37172 3780 37196 3782
rect 36956 3760 37252 3780
rect 37844 3641 37872 4762
rect 37924 4684 37976 4690
rect 37924 4626 37976 4632
rect 37936 4214 37964 4626
rect 38028 4282 38056 4966
rect 38120 4690 38148 5306
rect 38488 5166 38516 5732
rect 38568 5714 38620 5720
rect 39120 5772 39172 5778
rect 39120 5714 39172 5720
rect 38580 5166 38608 5714
rect 39132 5681 39160 5714
rect 39118 5672 39174 5681
rect 39118 5607 39174 5616
rect 39132 5166 39160 5607
rect 38476 5160 38528 5166
rect 38476 5102 38528 5108
rect 38568 5160 38620 5166
rect 38568 5102 38620 5108
rect 39120 5160 39172 5166
rect 39120 5102 39172 5108
rect 38488 4865 38516 5102
rect 38474 4856 38530 4865
rect 38474 4791 38530 4800
rect 38488 4758 38516 4791
rect 38476 4752 38528 4758
rect 38476 4694 38528 4700
rect 38580 4690 38608 5102
rect 39224 4729 39252 6190
rect 39764 5364 39816 5370
rect 39764 5306 39816 5312
rect 39776 5273 39804 5306
rect 39762 5264 39818 5273
rect 39762 5199 39764 5208
rect 39816 5199 39818 5208
rect 39764 5170 39816 5176
rect 39776 5139 39804 5170
rect 39210 4720 39266 4729
rect 38108 4684 38160 4690
rect 38108 4626 38160 4632
rect 38568 4684 38620 4690
rect 39210 4655 39266 4664
rect 38568 4626 38620 4632
rect 38016 4276 38068 4282
rect 38016 4218 38068 4224
rect 38580 4214 38608 4626
rect 39224 4622 39252 4655
rect 39212 4616 39264 4622
rect 39212 4558 39264 4564
rect 39224 4282 39252 4558
rect 39212 4276 39264 4282
rect 39212 4218 39264 4224
rect 37924 4208 37976 4214
rect 37924 4150 37976 4156
rect 38568 4208 38620 4214
rect 38568 4150 38620 4156
rect 37830 3632 37886 3641
rect 36176 3596 36228 3602
rect 37830 3567 37886 3576
rect 36176 3538 36228 3544
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 35254 3088 35310 3097
rect 35254 3023 35310 3032
rect 26200 2952 26202 2961
rect 26146 2887 26202 2896
rect 33138 2952 33194 2961
rect 33138 2887 33194 2896
rect 26160 2854 26188 2887
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 26148 2848 26200 2854
rect 36096 2836 36124 3470
rect 36188 3194 36216 3538
rect 36728 3392 36780 3398
rect 36728 3334 36780 3340
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 36176 2848 36228 2854
rect 36096 2808 36176 2836
rect 26148 2790 26200 2796
rect 36176 2790 36228 2796
rect 25700 2689 25728 2790
rect 25686 2680 25742 2689
rect 25686 2615 25742 2624
rect 36188 2553 36216 2790
rect 36634 2680 36690 2689
rect 36634 2615 36690 2624
rect 36174 2544 36230 2553
rect 36174 2479 36230 2488
rect 23662 2408 23718 2417
rect 23662 2343 23718 2352
rect 20626 1456 20682 1465
rect 20626 1391 20682 1400
rect 16762 54 16896 82
rect 23570 82 23626 480
rect 23676 82 23704 2343
rect 30010 1456 30066 1465
rect 30010 1391 30066 1400
rect 23570 54 23704 82
rect 30024 82 30052 1391
rect 30286 82 30342 480
rect 30024 54 30342 82
rect 36648 82 36676 2615
rect 36740 2514 36768 3334
rect 36956 2748 37252 2768
rect 37012 2746 37036 2748
rect 37092 2746 37116 2748
rect 37172 2746 37196 2748
rect 37034 2694 37036 2746
rect 37098 2694 37110 2746
rect 37172 2694 37174 2746
rect 37012 2692 37036 2694
rect 37092 2692 37116 2694
rect 37172 2692 37196 2694
rect 36956 2672 37252 2692
rect 46952 2650 46980 13518
rect 54956 10908 55252 10928
rect 55012 10906 55036 10908
rect 55092 10906 55116 10908
rect 55172 10906 55196 10908
rect 55034 10854 55036 10906
rect 55098 10854 55110 10906
rect 55172 10854 55174 10906
rect 55012 10852 55036 10854
rect 55092 10852 55116 10854
rect 55172 10852 55196 10854
rect 54956 10832 55252 10852
rect 54956 9820 55252 9840
rect 55012 9818 55036 9820
rect 55092 9818 55116 9820
rect 55172 9818 55196 9820
rect 55034 9766 55036 9818
rect 55098 9766 55110 9818
rect 55172 9766 55174 9818
rect 55012 9764 55036 9766
rect 55092 9764 55116 9766
rect 55172 9764 55196 9766
rect 54956 9744 55252 9764
rect 54956 8732 55252 8752
rect 55012 8730 55036 8732
rect 55092 8730 55116 8732
rect 55172 8730 55196 8732
rect 55034 8678 55036 8730
rect 55098 8678 55110 8730
rect 55172 8678 55174 8730
rect 55012 8676 55036 8678
rect 55092 8676 55116 8678
rect 55172 8676 55196 8678
rect 54956 8656 55252 8676
rect 54956 7644 55252 7664
rect 55012 7642 55036 7644
rect 55092 7642 55116 7644
rect 55172 7642 55196 7644
rect 55034 7590 55036 7642
rect 55098 7590 55110 7642
rect 55172 7590 55174 7642
rect 55012 7588 55036 7590
rect 55092 7588 55116 7590
rect 55172 7588 55196 7590
rect 54956 7568 55252 7588
rect 54956 6556 55252 6576
rect 55012 6554 55036 6556
rect 55092 6554 55116 6556
rect 55172 6554 55196 6556
rect 55034 6502 55036 6554
rect 55098 6502 55110 6554
rect 55172 6502 55174 6554
rect 55012 6500 55036 6502
rect 55092 6500 55116 6502
rect 55172 6500 55196 6502
rect 54956 6480 55252 6500
rect 51814 5944 51870 5953
rect 51814 5879 51870 5888
rect 59818 5944 59874 5953
rect 59818 5879 59874 5888
rect 60280 5908 60332 5914
rect 51828 5846 51856 5879
rect 59832 5846 59860 5879
rect 60280 5850 60332 5856
rect 51816 5840 51868 5846
rect 51816 5782 51868 5788
rect 59820 5840 59872 5846
rect 59820 5782 59872 5788
rect 51172 5704 51224 5710
rect 51828 5681 51856 5782
rect 51172 5646 51224 5652
rect 51814 5672 51870 5681
rect 51184 5234 51212 5646
rect 51814 5607 51870 5616
rect 54956 5468 55252 5488
rect 55012 5466 55036 5468
rect 55092 5466 55116 5468
rect 55172 5466 55196 5468
rect 55034 5414 55036 5466
rect 55098 5414 55110 5466
rect 55172 5414 55174 5466
rect 55012 5412 55036 5414
rect 55092 5412 55116 5414
rect 55172 5412 55196 5414
rect 54956 5392 55252 5412
rect 59832 5370 59860 5782
rect 60188 5704 60240 5710
rect 60188 5646 60240 5652
rect 60200 5370 60228 5646
rect 59820 5364 59872 5370
rect 59820 5306 59872 5312
rect 60188 5364 60240 5370
rect 60188 5306 60240 5312
rect 60200 5273 60228 5306
rect 60292 5302 60320 5850
rect 60372 5772 60424 5778
rect 60372 5714 60424 5720
rect 60280 5296 60332 5302
rect 60186 5264 60242 5273
rect 51172 5228 51224 5234
rect 60280 5238 60332 5244
rect 60186 5199 60242 5208
rect 51172 5170 51224 5176
rect 51184 5137 51212 5170
rect 51170 5128 51226 5137
rect 51170 5063 51226 5072
rect 49882 4856 49938 4865
rect 49882 4791 49938 4800
rect 49896 4758 49924 4791
rect 49884 4752 49936 4758
rect 51184 4729 51212 5063
rect 60384 5030 60412 5714
rect 60372 5024 60424 5030
rect 60372 4966 60424 4972
rect 56876 4820 56928 4826
rect 56876 4762 56928 4768
rect 49884 4694 49936 4700
rect 51170 4720 51226 4729
rect 49976 4684 50028 4690
rect 51170 4655 51226 4664
rect 49976 4626 50028 4632
rect 49988 3942 50016 4626
rect 52552 4480 52604 4486
rect 52552 4422 52604 4428
rect 49976 3936 50028 3942
rect 49976 3878 50028 3884
rect 49988 3777 50016 3878
rect 49974 3768 50030 3777
rect 49974 3703 50030 3712
rect 52564 3602 52592 4422
rect 54956 4380 55252 4400
rect 55012 4378 55036 4380
rect 55092 4378 55116 4380
rect 55172 4378 55196 4380
rect 55034 4326 55036 4378
rect 55098 4326 55110 4378
rect 55172 4326 55174 4378
rect 55012 4324 55036 4326
rect 55092 4324 55116 4326
rect 55172 4324 55196 4326
rect 54956 4304 55252 4324
rect 56888 3942 56916 4762
rect 57612 4616 57664 4622
rect 57612 4558 57664 4564
rect 57624 4282 57652 4558
rect 57612 4276 57664 4282
rect 57612 4218 57664 4224
rect 56876 3936 56928 3942
rect 56874 3904 56876 3913
rect 56928 3904 56930 3913
rect 56874 3839 56930 3848
rect 53932 3732 53984 3738
rect 53932 3674 53984 3680
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 52380 2854 52408 3470
rect 52564 3194 52592 3538
rect 52552 3188 52604 3194
rect 52552 3130 52604 3136
rect 52368 2848 52420 2854
rect 52368 2790 52420 2796
rect 53944 2650 53972 3674
rect 54956 3292 55252 3312
rect 55012 3290 55036 3292
rect 55092 3290 55116 3292
rect 55172 3290 55196 3292
rect 55034 3238 55036 3290
rect 55098 3238 55110 3290
rect 55172 3238 55174 3290
rect 55012 3236 55036 3238
rect 55092 3236 55116 3238
rect 55172 3236 55196 3238
rect 54956 3216 55252 3236
rect 56888 3097 56916 3839
rect 60384 3777 60412 4966
rect 60370 3768 60426 3777
rect 60752 3738 60780 13520
rect 72956 11452 73252 11472
rect 73012 11450 73036 11452
rect 73092 11450 73116 11452
rect 73172 11450 73196 11452
rect 73034 11398 73036 11450
rect 73098 11398 73110 11450
rect 73172 11398 73174 11450
rect 73012 11396 73036 11398
rect 73092 11396 73116 11398
rect 73172 11396 73196 11398
rect 72956 11376 73252 11396
rect 72956 10364 73252 10384
rect 73012 10362 73036 10364
rect 73092 10362 73116 10364
rect 73172 10362 73196 10364
rect 73034 10310 73036 10362
rect 73098 10310 73110 10362
rect 73172 10310 73174 10362
rect 73012 10308 73036 10310
rect 73092 10308 73116 10310
rect 73172 10308 73196 10310
rect 72956 10288 73252 10308
rect 74184 9382 74212 13520
rect 87694 13524 87750 14000
rect 87694 13520 87696 13524
rect 86960 13466 87012 13472
rect 87748 13520 87750 13524
rect 87696 13466 87748 13472
rect 100772 13518 101168 13546
rect 101218 13520 101274 14000
rect 73344 9376 73396 9382
rect 73344 9318 73396 9324
rect 74172 9376 74224 9382
rect 74172 9318 74224 9324
rect 72956 9276 73252 9296
rect 73012 9274 73036 9276
rect 73092 9274 73116 9276
rect 73172 9274 73196 9276
rect 73034 9222 73036 9274
rect 73098 9222 73110 9274
rect 73172 9222 73174 9274
rect 73012 9220 73036 9222
rect 73092 9220 73116 9222
rect 73172 9220 73196 9222
rect 72956 9200 73252 9220
rect 72956 8188 73252 8208
rect 73012 8186 73036 8188
rect 73092 8186 73116 8188
rect 73172 8186 73196 8188
rect 73034 8134 73036 8186
rect 73098 8134 73110 8186
rect 73172 8134 73174 8186
rect 73012 8132 73036 8134
rect 73092 8132 73116 8134
rect 73172 8132 73196 8134
rect 72956 8112 73252 8132
rect 72956 7100 73252 7120
rect 73012 7098 73036 7100
rect 73092 7098 73116 7100
rect 73172 7098 73196 7100
rect 73034 7046 73036 7098
rect 73098 7046 73110 7098
rect 73172 7046 73174 7098
rect 73012 7044 73036 7046
rect 73092 7044 73116 7046
rect 73172 7044 73196 7046
rect 72956 7024 73252 7044
rect 63132 6248 63184 6254
rect 63132 6190 63184 6196
rect 63144 5914 63172 6190
rect 72956 6012 73252 6032
rect 73012 6010 73036 6012
rect 73092 6010 73116 6012
rect 73172 6010 73196 6012
rect 73034 5958 73036 6010
rect 73098 5958 73110 6010
rect 73172 5958 73174 6010
rect 73012 5956 73036 5958
rect 73092 5956 73116 5958
rect 73172 5956 73196 5958
rect 72956 5936 73252 5956
rect 63132 5908 63184 5914
rect 63132 5850 63184 5856
rect 62856 5840 62908 5846
rect 62856 5782 62908 5788
rect 62764 5772 62816 5778
rect 62764 5714 62816 5720
rect 60924 5704 60976 5710
rect 60924 5646 60976 5652
rect 60936 4282 60964 5646
rect 61014 5536 61070 5545
rect 61014 5471 61070 5480
rect 61028 5370 61056 5471
rect 61016 5364 61068 5370
rect 61016 5306 61068 5312
rect 62776 5234 62804 5714
rect 62764 5228 62816 5234
rect 62764 5170 62816 5176
rect 62776 5137 62804 5170
rect 62762 5128 62818 5137
rect 62762 5063 62818 5072
rect 62868 4826 62896 5782
rect 63144 5370 63172 5850
rect 63222 5808 63278 5817
rect 63222 5743 63278 5752
rect 68836 5772 68888 5778
rect 63236 5710 63264 5743
rect 68836 5714 68888 5720
rect 63224 5704 63276 5710
rect 63224 5646 63276 5652
rect 63592 5704 63644 5710
rect 63592 5646 63644 5652
rect 68744 5704 68796 5710
rect 68744 5646 68796 5652
rect 63132 5364 63184 5370
rect 63132 5306 63184 5312
rect 63236 5098 63264 5646
rect 63224 5092 63276 5098
rect 63224 5034 63276 5040
rect 62856 4820 62908 4826
rect 62856 4762 62908 4768
rect 63604 4690 63632 5646
rect 68756 5545 68784 5646
rect 68742 5536 68798 5545
rect 68742 5471 68798 5480
rect 68756 5370 68784 5471
rect 68744 5364 68796 5370
rect 68744 5306 68796 5312
rect 68848 5030 68876 5714
rect 72792 5092 72844 5098
rect 72792 5034 72844 5040
rect 68836 5024 68888 5030
rect 72804 5001 72832 5034
rect 68836 4966 68888 4972
rect 72790 4992 72846 5001
rect 65800 4820 65852 4826
rect 65800 4762 65852 4768
rect 63592 4684 63644 4690
rect 63592 4626 63644 4632
rect 60924 4276 60976 4282
rect 60924 4218 60976 4224
rect 65812 3942 65840 4762
rect 68848 4729 68876 4966
rect 72790 4927 72846 4936
rect 72956 4924 73252 4944
rect 73012 4922 73036 4924
rect 73092 4922 73116 4924
rect 73172 4922 73196 4924
rect 73034 4870 73036 4922
rect 73098 4870 73110 4922
rect 73172 4870 73174 4922
rect 73012 4868 73036 4870
rect 73092 4868 73116 4870
rect 73172 4868 73196 4870
rect 72956 4848 73252 4868
rect 68834 4720 68890 4729
rect 66168 4684 66220 4690
rect 68834 4655 68890 4664
rect 66168 4626 66220 4632
rect 66180 4282 66208 4626
rect 66720 4480 66772 4486
rect 66720 4422 66772 4428
rect 66168 4276 66220 4282
rect 66168 4218 66220 4224
rect 65800 3936 65852 3942
rect 65798 3904 65800 3913
rect 65852 3904 65854 3913
rect 65798 3839 65854 3848
rect 60370 3703 60426 3712
rect 60740 3732 60792 3738
rect 60740 3674 60792 3680
rect 65812 3641 65840 3839
rect 65798 3632 65854 3641
rect 64696 3596 64748 3602
rect 66732 3602 66760 4422
rect 72956 3836 73252 3856
rect 73012 3834 73036 3836
rect 73092 3834 73116 3836
rect 73172 3834 73196 3836
rect 73034 3782 73036 3834
rect 73098 3782 73110 3834
rect 73172 3782 73174 3834
rect 73012 3780 73036 3782
rect 73092 3780 73116 3782
rect 73172 3780 73196 3782
rect 72956 3760 73252 3780
rect 65798 3567 65854 3576
rect 66720 3596 66772 3602
rect 64696 3538 64748 3544
rect 66720 3538 66772 3544
rect 64236 3528 64288 3534
rect 64236 3470 64288 3476
rect 56874 3088 56930 3097
rect 56874 3023 56930 3032
rect 64248 2854 64276 3470
rect 64708 3194 64736 3538
rect 67456 3392 67508 3398
rect 67456 3334 67508 3340
rect 64696 3188 64748 3194
rect 64696 3130 64748 3136
rect 67468 2961 67496 3334
rect 73356 2961 73384 9318
rect 77758 6352 77814 6361
rect 77758 6287 77814 6296
rect 77772 6254 77800 6287
rect 77760 6248 77812 6254
rect 77482 6216 77538 6225
rect 77760 6190 77812 6196
rect 77482 6151 77538 6160
rect 77496 6118 77524 6151
rect 77484 6112 77536 6118
rect 77484 6054 77536 6060
rect 77496 5914 77524 6054
rect 77484 5908 77536 5914
rect 77484 5850 77536 5856
rect 77496 5234 77524 5850
rect 77484 5228 77536 5234
rect 77484 5170 77536 5176
rect 79416 5228 79468 5234
rect 79416 5170 79468 5176
rect 77852 5160 77904 5166
rect 77390 5128 77446 5137
rect 77852 5102 77904 5108
rect 77484 5092 77536 5098
rect 77446 5072 77484 5080
rect 77390 5063 77484 5072
rect 77404 5052 77484 5063
rect 77404 4826 77432 5052
rect 77484 5034 77536 5040
rect 77392 4820 77444 4826
rect 77392 4762 77444 4768
rect 77864 4729 77892 5102
rect 78128 5092 78180 5098
rect 78128 5034 78180 5040
rect 77850 4720 77906 4729
rect 78140 4690 78168 5034
rect 79428 5030 79456 5170
rect 79416 5024 79468 5030
rect 79416 4966 79468 4972
rect 78956 4820 79008 4826
rect 78956 4762 79008 4768
rect 77850 4655 77906 4664
rect 78128 4684 78180 4690
rect 78128 4626 78180 4632
rect 78968 3942 78996 4762
rect 79232 4684 79284 4690
rect 79232 4626 79284 4632
rect 79244 4282 79272 4626
rect 79784 4480 79836 4486
rect 79784 4422 79836 4428
rect 79232 4276 79284 4282
rect 79232 4218 79284 4224
rect 78956 3936 79008 3942
rect 78954 3904 78956 3913
rect 79008 3904 79010 3913
rect 78954 3839 79010 3848
rect 78968 3641 78996 3839
rect 78954 3632 79010 3641
rect 78496 3596 78548 3602
rect 79796 3602 79824 4422
rect 86972 4049 87000 13466
rect 87708 13435 87736 13466
rect 90956 10908 91252 10928
rect 91012 10906 91036 10908
rect 91092 10906 91116 10908
rect 91172 10906 91196 10908
rect 91034 10854 91036 10906
rect 91098 10854 91110 10906
rect 91172 10854 91174 10906
rect 91012 10852 91036 10854
rect 91092 10852 91116 10854
rect 91172 10852 91196 10854
rect 90956 10832 91252 10852
rect 90956 9820 91252 9840
rect 91012 9818 91036 9820
rect 91092 9818 91116 9820
rect 91172 9818 91196 9820
rect 91034 9766 91036 9818
rect 91098 9766 91110 9818
rect 91172 9766 91174 9818
rect 91012 9764 91036 9766
rect 91092 9764 91116 9766
rect 91172 9764 91196 9766
rect 90956 9744 91252 9764
rect 90956 8732 91252 8752
rect 91012 8730 91036 8732
rect 91092 8730 91116 8732
rect 91172 8730 91196 8732
rect 91034 8678 91036 8730
rect 91098 8678 91110 8730
rect 91172 8678 91174 8730
rect 91012 8676 91036 8678
rect 91092 8676 91116 8678
rect 91172 8676 91196 8678
rect 90956 8656 91252 8676
rect 90956 7644 91252 7664
rect 91012 7642 91036 7644
rect 91092 7642 91116 7644
rect 91172 7642 91196 7644
rect 91034 7590 91036 7642
rect 91098 7590 91110 7642
rect 91172 7590 91174 7642
rect 91012 7588 91036 7590
rect 91092 7588 91116 7590
rect 91172 7588 91196 7590
rect 90956 7568 91252 7588
rect 90956 6556 91252 6576
rect 91012 6554 91036 6556
rect 91092 6554 91116 6556
rect 91172 6554 91196 6556
rect 91034 6502 91036 6554
rect 91098 6502 91110 6554
rect 91172 6502 91174 6554
rect 91012 6500 91036 6502
rect 91092 6500 91116 6502
rect 91172 6500 91196 6502
rect 90956 6480 91252 6500
rect 88062 5672 88118 5681
rect 88062 5607 88118 5616
rect 88076 5166 88104 5607
rect 88156 5568 88208 5574
rect 88156 5510 88208 5516
rect 88064 5160 88116 5166
rect 87970 5128 88026 5137
rect 87144 5092 87196 5098
rect 88064 5102 88116 5108
rect 88168 5098 88196 5510
rect 90956 5468 91252 5488
rect 91012 5466 91036 5468
rect 91092 5466 91116 5468
rect 91172 5466 91196 5468
rect 91034 5414 91036 5466
rect 91098 5414 91110 5466
rect 91172 5414 91174 5466
rect 91012 5412 91036 5414
rect 91092 5412 91116 5414
rect 91172 5412 91196 5414
rect 90956 5392 91252 5412
rect 87970 5063 88026 5072
rect 88156 5092 88208 5098
rect 87144 5034 87196 5040
rect 87156 4826 87184 5034
rect 87984 5030 88012 5063
rect 88156 5034 88208 5040
rect 88616 5092 88668 5098
rect 88616 5034 88668 5040
rect 87972 5024 88024 5030
rect 88168 5001 88196 5034
rect 87972 4966 88024 4972
rect 88154 4992 88210 5001
rect 87984 4826 88012 4966
rect 88154 4927 88210 4936
rect 87144 4820 87196 4826
rect 87144 4762 87196 4768
rect 87972 4820 88024 4826
rect 87972 4762 88024 4768
rect 88628 4622 88656 5034
rect 89810 4992 89866 5001
rect 89810 4927 89866 4936
rect 88706 4856 88762 4865
rect 88706 4791 88762 4800
rect 88720 4758 88748 4791
rect 88708 4752 88760 4758
rect 88708 4694 88760 4700
rect 88616 4616 88668 4622
rect 88616 4558 88668 4564
rect 88628 4282 88656 4558
rect 88616 4276 88668 4282
rect 88616 4218 88668 4224
rect 88720 4214 88748 4694
rect 89168 4480 89220 4486
rect 89168 4422 89220 4428
rect 88708 4208 88760 4214
rect 88708 4150 88760 4156
rect 80702 4040 80758 4049
rect 80702 3975 80758 3984
rect 86958 4040 87014 4049
rect 86958 3975 87014 3984
rect 78954 3567 79010 3576
rect 79784 3596 79836 3602
rect 78496 3538 78548 3544
rect 79784 3538 79836 3544
rect 78036 3528 78088 3534
rect 78036 3470 78088 3476
rect 67454 2952 67510 2961
rect 67454 2887 67510 2896
rect 73342 2952 73398 2961
rect 78048 2922 78076 3470
rect 78508 3194 78536 3538
rect 80716 3398 80744 3975
rect 88720 3913 88748 4150
rect 88706 3904 88762 3913
rect 88706 3839 88762 3848
rect 88708 3596 88760 3602
rect 88708 3538 88760 3544
rect 80704 3392 80756 3398
rect 80704 3334 80756 3340
rect 80716 3194 80744 3334
rect 78496 3188 78548 3194
rect 78496 3130 78548 3136
rect 80704 3188 80756 3194
rect 80704 3130 80756 3136
rect 80716 2990 80744 3130
rect 80704 2984 80756 2990
rect 80704 2926 80756 2932
rect 73342 2887 73398 2896
rect 78036 2916 78088 2922
rect 57060 2848 57112 2854
rect 57060 2790 57112 2796
rect 64236 2848 64288 2854
rect 64236 2790 64288 2796
rect 46940 2644 46992 2650
rect 46940 2586 46992 2592
rect 53932 2644 53984 2650
rect 53932 2586 53984 2592
rect 43902 2544 43958 2553
rect 36728 2508 36780 2514
rect 43902 2479 43958 2488
rect 36728 2450 36780 2456
rect 39488 2304 39540 2310
rect 39488 2246 39540 2252
rect 39500 1329 39528 2246
rect 39486 1320 39542 1329
rect 39486 1255 39542 1264
rect 37002 82 37058 480
rect 36648 54 37058 82
rect 16762 0 16818 54
rect 23570 0 23626 54
rect 30286 0 30342 54
rect 37002 0 37058 54
rect 43810 82 43866 480
rect 43916 82 43944 2479
rect 53472 2304 53524 2310
rect 53472 2246 53524 2252
rect 53484 1329 53512 2246
rect 54956 2204 55252 2224
rect 55012 2202 55036 2204
rect 55092 2202 55116 2204
rect 55172 2202 55196 2204
rect 55034 2150 55036 2202
rect 55098 2150 55110 2202
rect 55172 2150 55174 2202
rect 55012 2148 55036 2150
rect 55092 2148 55116 2150
rect 55172 2148 55196 2150
rect 54956 2128 55252 2148
rect 50250 1320 50306 1329
rect 50250 1255 50306 1264
rect 53470 1320 53526 1329
rect 53470 1255 53526 1264
rect 43810 54 43944 82
rect 50264 82 50292 1255
rect 50526 82 50582 480
rect 50264 54 50582 82
rect 57072 82 57100 2790
rect 67468 2650 67496 2887
rect 78036 2858 78088 2864
rect 84384 2916 84436 2922
rect 84384 2858 84436 2864
rect 70492 2848 70544 2854
rect 70492 2790 70544 2796
rect 80244 2848 80296 2854
rect 80244 2790 80296 2796
rect 67364 2644 67416 2650
rect 67364 2586 67416 2592
rect 67456 2644 67508 2650
rect 67456 2586 67508 2592
rect 67376 2417 67404 2586
rect 67362 2408 67418 2417
rect 67362 2343 67418 2352
rect 64142 1320 64198 1329
rect 64142 1255 64198 1264
rect 57334 82 57390 480
rect 57072 54 57390 82
rect 43810 0 43866 54
rect 50526 0 50582 54
rect 57334 0 57390 54
rect 64050 82 64106 480
rect 64156 82 64184 1255
rect 64050 54 64184 82
rect 70504 82 70532 2790
rect 72956 2748 73252 2768
rect 73012 2746 73036 2748
rect 73092 2746 73116 2748
rect 73172 2746 73196 2748
rect 73034 2694 73036 2746
rect 73098 2694 73110 2746
rect 73172 2694 73174 2746
rect 73012 2692 73036 2694
rect 73092 2692 73116 2694
rect 73172 2692 73196 2694
rect 72956 2672 73252 2692
rect 80256 2689 80284 2790
rect 80242 2680 80298 2689
rect 80242 2615 80298 2624
rect 77298 2408 77354 2417
rect 77298 2343 77354 2352
rect 70766 82 70822 480
rect 70504 54 70822 82
rect 77312 82 77340 2343
rect 77574 82 77630 480
rect 77312 54 77630 82
rect 64050 0 64106 54
rect 70766 0 70822 54
rect 77574 0 77630 54
rect 84290 82 84346 480
rect 84396 82 84424 2858
rect 88720 2854 88748 3538
rect 89180 3534 89208 4422
rect 89168 3528 89220 3534
rect 88890 3496 88946 3505
rect 89168 3470 89220 3476
rect 88890 3431 88946 3440
rect 88904 3398 88932 3431
rect 88892 3392 88944 3398
rect 88892 3334 88944 3340
rect 88904 3194 88932 3334
rect 89180 3194 89208 3470
rect 88892 3188 88944 3194
rect 88892 3130 88944 3136
rect 89168 3188 89220 3194
rect 89168 3130 89220 3136
rect 88248 2848 88300 2854
rect 88248 2790 88300 2796
rect 88708 2848 88760 2854
rect 88708 2790 88760 2796
rect 88260 2417 88288 2790
rect 88246 2408 88302 2417
rect 88246 2343 88302 2352
rect 88720 1465 88748 2790
rect 88706 1456 88762 1465
rect 88706 1391 88762 1400
rect 89824 105 89852 4927
rect 90956 4380 91252 4400
rect 91012 4378 91036 4380
rect 91092 4378 91116 4380
rect 91172 4378 91196 4380
rect 91034 4326 91036 4378
rect 91098 4326 91110 4378
rect 91172 4326 91174 4378
rect 91012 4324 91036 4326
rect 91092 4324 91116 4326
rect 91172 4324 91196 4326
rect 90956 4304 91252 4324
rect 100772 3505 100800 13518
rect 101140 13410 101168 13518
rect 101232 13410 101260 13520
rect 101140 13382 101260 13410
rect 104162 12744 104218 12753
rect 104162 12679 104218 12688
rect 104176 4865 104204 12679
rect 107474 10432 107530 10441
rect 107474 10367 107530 10376
rect 107290 8120 107346 8129
rect 107290 8055 107346 8064
rect 107304 5137 107332 8055
rect 107488 6225 107516 10367
rect 107474 6216 107530 6225
rect 107474 6151 107530 6160
rect 107290 5128 107346 5137
rect 107290 5063 107346 5072
rect 104162 4856 104218 4865
rect 104162 4791 104218 4800
rect 100758 3496 100814 3505
rect 100758 3431 100814 3440
rect 90956 3292 91252 3312
rect 91012 3290 91036 3292
rect 91092 3290 91116 3292
rect 91172 3290 91196 3292
rect 91034 3238 91036 3290
rect 91098 3238 91110 3290
rect 91172 3238 91174 3290
rect 91012 3236 91036 3238
rect 91092 3236 91116 3238
rect 91172 3236 91196 3238
rect 90956 3216 91252 3236
rect 90730 2680 90786 2689
rect 90730 2615 90786 2624
rect 84290 54 84424 82
rect 89810 96 89866 105
rect 84290 0 84346 54
rect 90744 82 90772 2615
rect 104622 2408 104678 2417
rect 104622 2343 104678 2352
rect 90956 2204 91252 2224
rect 91012 2202 91036 2204
rect 91092 2202 91116 2204
rect 91172 2202 91196 2204
rect 91034 2150 91036 2202
rect 91098 2150 91110 2202
rect 91172 2150 91174 2202
rect 91012 2148 91036 2150
rect 91092 2148 91116 2150
rect 91172 2148 91196 2150
rect 90956 2128 91252 2148
rect 97538 1456 97594 1465
rect 97538 1391 97594 1400
rect 91006 82 91062 480
rect 90744 54 91062 82
rect 97552 82 97580 1391
rect 97814 82 97870 480
rect 97552 54 97870 82
rect 89810 31 89866 40
rect 91006 0 91062 54
rect 97814 0 97870 54
rect 104530 82 104586 480
rect 104636 82 104664 2343
rect 105542 1184 105598 1193
rect 105542 1119 105598 1128
rect 105556 105 105584 1119
rect 104530 54 104664 82
rect 105542 96 105598 105
rect 104530 0 104586 54
rect 105542 31 105598 40
<< via2 >>
rect 4526 5208 4582 5264
rect 18956 10906 19012 10908
rect 19036 10906 19092 10908
rect 19116 10906 19172 10908
rect 19196 10906 19252 10908
rect 18956 10854 18982 10906
rect 18982 10854 19012 10906
rect 19036 10854 19046 10906
rect 19046 10854 19092 10906
rect 19116 10854 19162 10906
rect 19162 10854 19172 10906
rect 19196 10854 19226 10906
rect 19226 10854 19252 10906
rect 18956 10852 19012 10854
rect 19036 10852 19092 10854
rect 19116 10852 19172 10854
rect 19196 10852 19252 10854
rect 18956 9818 19012 9820
rect 19036 9818 19092 9820
rect 19116 9818 19172 9820
rect 19196 9818 19252 9820
rect 18956 9766 18982 9818
rect 18982 9766 19012 9818
rect 19036 9766 19046 9818
rect 19046 9766 19092 9818
rect 19116 9766 19162 9818
rect 19162 9766 19172 9818
rect 19196 9766 19226 9818
rect 19226 9766 19252 9818
rect 18956 9764 19012 9766
rect 19036 9764 19092 9766
rect 19116 9764 19172 9766
rect 19196 9764 19252 9766
rect 18956 8730 19012 8732
rect 19036 8730 19092 8732
rect 19116 8730 19172 8732
rect 19196 8730 19252 8732
rect 18956 8678 18982 8730
rect 18982 8678 19012 8730
rect 19036 8678 19046 8730
rect 19046 8678 19092 8730
rect 19116 8678 19162 8730
rect 19162 8678 19172 8730
rect 19196 8678 19226 8730
rect 19226 8678 19252 8730
rect 18956 8676 19012 8678
rect 19036 8676 19092 8678
rect 19116 8676 19172 8678
rect 19196 8676 19252 8678
rect 18956 7642 19012 7644
rect 19036 7642 19092 7644
rect 19116 7642 19172 7644
rect 19196 7642 19252 7644
rect 18956 7590 18982 7642
rect 18982 7590 19012 7642
rect 19036 7590 19046 7642
rect 19046 7590 19092 7642
rect 19116 7590 19162 7642
rect 19162 7590 19172 7642
rect 19196 7590 19226 7642
rect 19226 7590 19252 7642
rect 18956 7588 19012 7590
rect 19036 7588 19092 7590
rect 19116 7588 19172 7590
rect 19196 7588 19252 7590
rect 18956 6554 19012 6556
rect 19036 6554 19092 6556
rect 19116 6554 19172 6556
rect 19196 6554 19252 6556
rect 18956 6502 18982 6554
rect 18982 6502 19012 6554
rect 19036 6502 19046 6554
rect 19046 6502 19092 6554
rect 19116 6502 19162 6554
rect 19162 6502 19172 6554
rect 19196 6502 19226 6554
rect 19226 6502 19252 6554
rect 18956 6500 19012 6502
rect 19036 6500 19092 6502
rect 19116 6500 19172 6502
rect 19196 6500 19252 6502
rect 18956 5466 19012 5468
rect 19036 5466 19092 5468
rect 19116 5466 19172 5468
rect 19196 5466 19252 5468
rect 18956 5414 18982 5466
rect 18982 5414 19012 5466
rect 19036 5414 19046 5466
rect 19046 5414 19092 5466
rect 19116 5414 19162 5466
rect 19162 5414 19172 5466
rect 19196 5414 19226 5466
rect 19226 5414 19252 5466
rect 18956 5412 19012 5414
rect 19036 5412 19092 5414
rect 19116 5412 19172 5414
rect 19196 5412 19252 5414
rect 18050 5072 18106 5128
rect 4894 3848 4950 3904
rect 2318 3576 2374 3632
rect 1582 1400 1638 1456
rect 12438 3984 12494 4040
rect 18956 4378 19012 4380
rect 19036 4378 19092 4380
rect 19116 4378 19172 4380
rect 19196 4378 19252 4380
rect 18956 4326 18982 4378
rect 18982 4326 19012 4378
rect 19036 4326 19046 4378
rect 19046 4326 19092 4378
rect 19116 4326 19162 4378
rect 19162 4326 19172 4378
rect 19196 4326 19226 4378
rect 19226 4326 19252 4378
rect 18956 4324 19012 4326
rect 19036 4324 19092 4326
rect 19116 4324 19172 4326
rect 19196 4324 19252 4326
rect 19338 3984 19394 4040
rect 17774 3848 17830 3904
rect 18956 3290 19012 3292
rect 19036 3290 19092 3292
rect 19116 3290 19172 3292
rect 19196 3290 19252 3292
rect 18956 3238 18982 3290
rect 18982 3238 19012 3290
rect 19036 3238 19046 3290
rect 19046 3238 19092 3290
rect 19116 3238 19162 3290
rect 19162 3238 19172 3290
rect 19196 3238 19226 3290
rect 19226 3238 19252 3290
rect 18956 3236 19012 3238
rect 19036 3236 19092 3238
rect 19116 3236 19172 3238
rect 19196 3236 19252 3238
rect 6826 2488 6882 2544
rect 16854 2488 16910 2544
rect 12622 2352 12678 2408
rect 9770 1400 9826 1456
rect 18956 2202 19012 2204
rect 19036 2202 19092 2204
rect 19116 2202 19172 2204
rect 19196 2202 19252 2204
rect 18956 2150 18982 2202
rect 18982 2150 19012 2202
rect 19036 2150 19046 2202
rect 19046 2150 19092 2202
rect 19116 2150 19162 2202
rect 19162 2150 19172 2202
rect 19196 2150 19226 2202
rect 19226 2150 19252 2202
rect 18956 2148 19012 2150
rect 19036 2148 19092 2150
rect 19116 2148 19172 2150
rect 19196 2148 19252 2150
rect 36956 11450 37012 11452
rect 37036 11450 37092 11452
rect 37116 11450 37172 11452
rect 37196 11450 37252 11452
rect 36956 11398 36982 11450
rect 36982 11398 37012 11450
rect 37036 11398 37046 11450
rect 37046 11398 37092 11450
rect 37116 11398 37162 11450
rect 37162 11398 37172 11450
rect 37196 11398 37226 11450
rect 37226 11398 37252 11450
rect 36956 11396 37012 11398
rect 37036 11396 37092 11398
rect 37116 11396 37172 11398
rect 37196 11396 37252 11398
rect 36956 10362 37012 10364
rect 37036 10362 37092 10364
rect 37116 10362 37172 10364
rect 37196 10362 37252 10364
rect 36956 10310 36982 10362
rect 36982 10310 37012 10362
rect 37036 10310 37046 10362
rect 37046 10310 37092 10362
rect 37116 10310 37162 10362
rect 37162 10310 37172 10362
rect 37196 10310 37226 10362
rect 37226 10310 37252 10362
rect 36956 10308 37012 10310
rect 37036 10308 37092 10310
rect 37116 10308 37172 10310
rect 37196 10308 37252 10310
rect 36956 9274 37012 9276
rect 37036 9274 37092 9276
rect 37116 9274 37172 9276
rect 37196 9274 37252 9276
rect 36956 9222 36982 9274
rect 36982 9222 37012 9274
rect 37036 9222 37046 9274
rect 37046 9222 37092 9274
rect 37116 9222 37162 9274
rect 37162 9222 37172 9274
rect 37196 9222 37226 9274
rect 37226 9222 37252 9274
rect 36956 9220 37012 9222
rect 37036 9220 37092 9222
rect 37116 9220 37172 9222
rect 37196 9220 37252 9222
rect 36956 8186 37012 8188
rect 37036 8186 37092 8188
rect 37116 8186 37172 8188
rect 37196 8186 37252 8188
rect 36956 8134 36982 8186
rect 36982 8134 37012 8186
rect 37036 8134 37046 8186
rect 37046 8134 37092 8186
rect 37116 8134 37162 8186
rect 37162 8134 37172 8186
rect 37196 8134 37226 8186
rect 37226 8134 37252 8186
rect 36956 8132 37012 8134
rect 37036 8132 37092 8134
rect 37116 8132 37172 8134
rect 37196 8132 37252 8134
rect 36956 7098 37012 7100
rect 37036 7098 37092 7100
rect 37116 7098 37172 7100
rect 37196 7098 37252 7100
rect 36956 7046 36982 7098
rect 36982 7046 37012 7098
rect 37036 7046 37046 7098
rect 37046 7046 37092 7098
rect 37116 7046 37162 7098
rect 37162 7046 37172 7098
rect 37196 7046 37226 7098
rect 37226 7046 37252 7098
rect 36956 7044 37012 7046
rect 37036 7044 37092 7046
rect 37116 7044 37172 7046
rect 37196 7044 37252 7046
rect 38566 6296 38622 6352
rect 36956 6010 37012 6012
rect 37036 6010 37092 6012
rect 37116 6010 37172 6012
rect 37196 6010 37252 6012
rect 36956 5958 36982 6010
rect 36982 5958 37012 6010
rect 37036 5958 37046 6010
rect 37046 5958 37092 6010
rect 37116 5958 37162 6010
rect 37162 5958 37172 6010
rect 37196 5958 37226 6010
rect 37226 5958 37252 6010
rect 36956 5956 37012 5958
rect 37036 5956 37092 5958
rect 37116 5956 37172 5958
rect 37196 5956 37252 5958
rect 36956 4922 37012 4924
rect 37036 4922 37092 4924
rect 37116 4922 37172 4924
rect 37196 4922 37252 4924
rect 36956 4870 36982 4922
rect 36982 4870 37012 4922
rect 37036 4870 37046 4922
rect 37046 4870 37092 4922
rect 37116 4870 37162 4922
rect 37162 4870 37172 4922
rect 37196 4870 37226 4922
rect 37226 4870 37252 4922
rect 36956 4868 37012 4870
rect 37036 4868 37092 4870
rect 37116 4868 37172 4870
rect 37196 4868 37252 4870
rect 37646 5208 37702 5264
rect 38106 5752 38162 5808
rect 37830 5072 37886 5128
rect 35254 3884 35256 3904
rect 35256 3884 35308 3904
rect 35308 3884 35310 3904
rect 35254 3848 35310 3884
rect 36956 3834 37012 3836
rect 37036 3834 37092 3836
rect 37116 3834 37172 3836
rect 37196 3834 37252 3836
rect 36956 3782 36982 3834
rect 36982 3782 37012 3834
rect 37036 3782 37046 3834
rect 37046 3782 37092 3834
rect 37116 3782 37162 3834
rect 37162 3782 37172 3834
rect 37196 3782 37226 3834
rect 37226 3782 37252 3834
rect 36956 3780 37012 3782
rect 37036 3780 37092 3782
rect 37116 3780 37172 3782
rect 37196 3780 37252 3782
rect 39118 5616 39174 5672
rect 38474 4800 38530 4856
rect 39762 5228 39818 5264
rect 39762 5208 39764 5228
rect 39764 5208 39816 5228
rect 39816 5208 39818 5228
rect 39210 4664 39266 4720
rect 37830 3576 37886 3632
rect 35254 3032 35310 3088
rect 26146 2932 26148 2952
rect 26148 2932 26200 2952
rect 26200 2932 26202 2952
rect 26146 2896 26202 2932
rect 33138 2896 33194 2952
rect 25686 2624 25742 2680
rect 36634 2624 36690 2680
rect 36174 2488 36230 2544
rect 23662 2352 23718 2408
rect 20626 1400 20682 1456
rect 30010 1400 30066 1456
rect 36956 2746 37012 2748
rect 37036 2746 37092 2748
rect 37116 2746 37172 2748
rect 37196 2746 37252 2748
rect 36956 2694 36982 2746
rect 36982 2694 37012 2746
rect 37036 2694 37046 2746
rect 37046 2694 37092 2746
rect 37116 2694 37162 2746
rect 37162 2694 37172 2746
rect 37196 2694 37226 2746
rect 37226 2694 37252 2746
rect 36956 2692 37012 2694
rect 37036 2692 37092 2694
rect 37116 2692 37172 2694
rect 37196 2692 37252 2694
rect 54956 10906 55012 10908
rect 55036 10906 55092 10908
rect 55116 10906 55172 10908
rect 55196 10906 55252 10908
rect 54956 10854 54982 10906
rect 54982 10854 55012 10906
rect 55036 10854 55046 10906
rect 55046 10854 55092 10906
rect 55116 10854 55162 10906
rect 55162 10854 55172 10906
rect 55196 10854 55226 10906
rect 55226 10854 55252 10906
rect 54956 10852 55012 10854
rect 55036 10852 55092 10854
rect 55116 10852 55172 10854
rect 55196 10852 55252 10854
rect 54956 9818 55012 9820
rect 55036 9818 55092 9820
rect 55116 9818 55172 9820
rect 55196 9818 55252 9820
rect 54956 9766 54982 9818
rect 54982 9766 55012 9818
rect 55036 9766 55046 9818
rect 55046 9766 55092 9818
rect 55116 9766 55162 9818
rect 55162 9766 55172 9818
rect 55196 9766 55226 9818
rect 55226 9766 55252 9818
rect 54956 9764 55012 9766
rect 55036 9764 55092 9766
rect 55116 9764 55172 9766
rect 55196 9764 55252 9766
rect 54956 8730 55012 8732
rect 55036 8730 55092 8732
rect 55116 8730 55172 8732
rect 55196 8730 55252 8732
rect 54956 8678 54982 8730
rect 54982 8678 55012 8730
rect 55036 8678 55046 8730
rect 55046 8678 55092 8730
rect 55116 8678 55162 8730
rect 55162 8678 55172 8730
rect 55196 8678 55226 8730
rect 55226 8678 55252 8730
rect 54956 8676 55012 8678
rect 55036 8676 55092 8678
rect 55116 8676 55172 8678
rect 55196 8676 55252 8678
rect 54956 7642 55012 7644
rect 55036 7642 55092 7644
rect 55116 7642 55172 7644
rect 55196 7642 55252 7644
rect 54956 7590 54982 7642
rect 54982 7590 55012 7642
rect 55036 7590 55046 7642
rect 55046 7590 55092 7642
rect 55116 7590 55162 7642
rect 55162 7590 55172 7642
rect 55196 7590 55226 7642
rect 55226 7590 55252 7642
rect 54956 7588 55012 7590
rect 55036 7588 55092 7590
rect 55116 7588 55172 7590
rect 55196 7588 55252 7590
rect 54956 6554 55012 6556
rect 55036 6554 55092 6556
rect 55116 6554 55172 6556
rect 55196 6554 55252 6556
rect 54956 6502 54982 6554
rect 54982 6502 55012 6554
rect 55036 6502 55046 6554
rect 55046 6502 55092 6554
rect 55116 6502 55162 6554
rect 55162 6502 55172 6554
rect 55196 6502 55226 6554
rect 55226 6502 55252 6554
rect 54956 6500 55012 6502
rect 55036 6500 55092 6502
rect 55116 6500 55172 6502
rect 55196 6500 55252 6502
rect 51814 5888 51870 5944
rect 59818 5888 59874 5944
rect 51814 5616 51870 5672
rect 54956 5466 55012 5468
rect 55036 5466 55092 5468
rect 55116 5466 55172 5468
rect 55196 5466 55252 5468
rect 54956 5414 54982 5466
rect 54982 5414 55012 5466
rect 55036 5414 55046 5466
rect 55046 5414 55092 5466
rect 55116 5414 55162 5466
rect 55162 5414 55172 5466
rect 55196 5414 55226 5466
rect 55226 5414 55252 5466
rect 54956 5412 55012 5414
rect 55036 5412 55092 5414
rect 55116 5412 55172 5414
rect 55196 5412 55252 5414
rect 60186 5208 60242 5264
rect 51170 5072 51226 5128
rect 49882 4800 49938 4856
rect 51170 4664 51226 4720
rect 49974 3712 50030 3768
rect 54956 4378 55012 4380
rect 55036 4378 55092 4380
rect 55116 4378 55172 4380
rect 55196 4378 55252 4380
rect 54956 4326 54982 4378
rect 54982 4326 55012 4378
rect 55036 4326 55046 4378
rect 55046 4326 55092 4378
rect 55116 4326 55162 4378
rect 55162 4326 55172 4378
rect 55196 4326 55226 4378
rect 55226 4326 55252 4378
rect 54956 4324 55012 4326
rect 55036 4324 55092 4326
rect 55116 4324 55172 4326
rect 55196 4324 55252 4326
rect 56874 3884 56876 3904
rect 56876 3884 56928 3904
rect 56928 3884 56930 3904
rect 56874 3848 56930 3884
rect 54956 3290 55012 3292
rect 55036 3290 55092 3292
rect 55116 3290 55172 3292
rect 55196 3290 55252 3292
rect 54956 3238 54982 3290
rect 54982 3238 55012 3290
rect 55036 3238 55046 3290
rect 55046 3238 55092 3290
rect 55116 3238 55162 3290
rect 55162 3238 55172 3290
rect 55196 3238 55226 3290
rect 55226 3238 55252 3290
rect 54956 3236 55012 3238
rect 55036 3236 55092 3238
rect 55116 3236 55172 3238
rect 55196 3236 55252 3238
rect 60370 3712 60426 3768
rect 72956 11450 73012 11452
rect 73036 11450 73092 11452
rect 73116 11450 73172 11452
rect 73196 11450 73252 11452
rect 72956 11398 72982 11450
rect 72982 11398 73012 11450
rect 73036 11398 73046 11450
rect 73046 11398 73092 11450
rect 73116 11398 73162 11450
rect 73162 11398 73172 11450
rect 73196 11398 73226 11450
rect 73226 11398 73252 11450
rect 72956 11396 73012 11398
rect 73036 11396 73092 11398
rect 73116 11396 73172 11398
rect 73196 11396 73252 11398
rect 72956 10362 73012 10364
rect 73036 10362 73092 10364
rect 73116 10362 73172 10364
rect 73196 10362 73252 10364
rect 72956 10310 72982 10362
rect 72982 10310 73012 10362
rect 73036 10310 73046 10362
rect 73046 10310 73092 10362
rect 73116 10310 73162 10362
rect 73162 10310 73172 10362
rect 73196 10310 73226 10362
rect 73226 10310 73252 10362
rect 72956 10308 73012 10310
rect 73036 10308 73092 10310
rect 73116 10308 73172 10310
rect 73196 10308 73252 10310
rect 72956 9274 73012 9276
rect 73036 9274 73092 9276
rect 73116 9274 73172 9276
rect 73196 9274 73252 9276
rect 72956 9222 72982 9274
rect 72982 9222 73012 9274
rect 73036 9222 73046 9274
rect 73046 9222 73092 9274
rect 73116 9222 73162 9274
rect 73162 9222 73172 9274
rect 73196 9222 73226 9274
rect 73226 9222 73252 9274
rect 72956 9220 73012 9222
rect 73036 9220 73092 9222
rect 73116 9220 73172 9222
rect 73196 9220 73252 9222
rect 72956 8186 73012 8188
rect 73036 8186 73092 8188
rect 73116 8186 73172 8188
rect 73196 8186 73252 8188
rect 72956 8134 72982 8186
rect 72982 8134 73012 8186
rect 73036 8134 73046 8186
rect 73046 8134 73092 8186
rect 73116 8134 73162 8186
rect 73162 8134 73172 8186
rect 73196 8134 73226 8186
rect 73226 8134 73252 8186
rect 72956 8132 73012 8134
rect 73036 8132 73092 8134
rect 73116 8132 73172 8134
rect 73196 8132 73252 8134
rect 72956 7098 73012 7100
rect 73036 7098 73092 7100
rect 73116 7098 73172 7100
rect 73196 7098 73252 7100
rect 72956 7046 72982 7098
rect 72982 7046 73012 7098
rect 73036 7046 73046 7098
rect 73046 7046 73092 7098
rect 73116 7046 73162 7098
rect 73162 7046 73172 7098
rect 73196 7046 73226 7098
rect 73226 7046 73252 7098
rect 72956 7044 73012 7046
rect 73036 7044 73092 7046
rect 73116 7044 73172 7046
rect 73196 7044 73252 7046
rect 72956 6010 73012 6012
rect 73036 6010 73092 6012
rect 73116 6010 73172 6012
rect 73196 6010 73252 6012
rect 72956 5958 72982 6010
rect 72982 5958 73012 6010
rect 73036 5958 73046 6010
rect 73046 5958 73092 6010
rect 73116 5958 73162 6010
rect 73162 5958 73172 6010
rect 73196 5958 73226 6010
rect 73226 5958 73252 6010
rect 72956 5956 73012 5958
rect 73036 5956 73092 5958
rect 73116 5956 73172 5958
rect 73196 5956 73252 5958
rect 61014 5480 61070 5536
rect 62762 5072 62818 5128
rect 63222 5752 63278 5808
rect 68742 5480 68798 5536
rect 72790 4936 72846 4992
rect 72956 4922 73012 4924
rect 73036 4922 73092 4924
rect 73116 4922 73172 4924
rect 73196 4922 73252 4924
rect 72956 4870 72982 4922
rect 72982 4870 73012 4922
rect 73036 4870 73046 4922
rect 73046 4870 73092 4922
rect 73116 4870 73162 4922
rect 73162 4870 73172 4922
rect 73196 4870 73226 4922
rect 73226 4870 73252 4922
rect 72956 4868 73012 4870
rect 73036 4868 73092 4870
rect 73116 4868 73172 4870
rect 73196 4868 73252 4870
rect 68834 4664 68890 4720
rect 65798 3884 65800 3904
rect 65800 3884 65852 3904
rect 65852 3884 65854 3904
rect 65798 3848 65854 3884
rect 65798 3576 65854 3632
rect 72956 3834 73012 3836
rect 73036 3834 73092 3836
rect 73116 3834 73172 3836
rect 73196 3834 73252 3836
rect 72956 3782 72982 3834
rect 72982 3782 73012 3834
rect 73036 3782 73046 3834
rect 73046 3782 73092 3834
rect 73116 3782 73162 3834
rect 73162 3782 73172 3834
rect 73196 3782 73226 3834
rect 73226 3782 73252 3834
rect 72956 3780 73012 3782
rect 73036 3780 73092 3782
rect 73116 3780 73172 3782
rect 73196 3780 73252 3782
rect 56874 3032 56930 3088
rect 77758 6296 77814 6352
rect 77482 6160 77538 6216
rect 77390 5072 77446 5128
rect 77850 4664 77906 4720
rect 78954 3884 78956 3904
rect 78956 3884 79008 3904
rect 79008 3884 79010 3904
rect 78954 3848 79010 3884
rect 78954 3576 79010 3632
rect 90956 10906 91012 10908
rect 91036 10906 91092 10908
rect 91116 10906 91172 10908
rect 91196 10906 91252 10908
rect 90956 10854 90982 10906
rect 90982 10854 91012 10906
rect 91036 10854 91046 10906
rect 91046 10854 91092 10906
rect 91116 10854 91162 10906
rect 91162 10854 91172 10906
rect 91196 10854 91226 10906
rect 91226 10854 91252 10906
rect 90956 10852 91012 10854
rect 91036 10852 91092 10854
rect 91116 10852 91172 10854
rect 91196 10852 91252 10854
rect 90956 9818 91012 9820
rect 91036 9818 91092 9820
rect 91116 9818 91172 9820
rect 91196 9818 91252 9820
rect 90956 9766 90982 9818
rect 90982 9766 91012 9818
rect 91036 9766 91046 9818
rect 91046 9766 91092 9818
rect 91116 9766 91162 9818
rect 91162 9766 91172 9818
rect 91196 9766 91226 9818
rect 91226 9766 91252 9818
rect 90956 9764 91012 9766
rect 91036 9764 91092 9766
rect 91116 9764 91172 9766
rect 91196 9764 91252 9766
rect 90956 8730 91012 8732
rect 91036 8730 91092 8732
rect 91116 8730 91172 8732
rect 91196 8730 91252 8732
rect 90956 8678 90982 8730
rect 90982 8678 91012 8730
rect 91036 8678 91046 8730
rect 91046 8678 91092 8730
rect 91116 8678 91162 8730
rect 91162 8678 91172 8730
rect 91196 8678 91226 8730
rect 91226 8678 91252 8730
rect 90956 8676 91012 8678
rect 91036 8676 91092 8678
rect 91116 8676 91172 8678
rect 91196 8676 91252 8678
rect 90956 7642 91012 7644
rect 91036 7642 91092 7644
rect 91116 7642 91172 7644
rect 91196 7642 91252 7644
rect 90956 7590 90982 7642
rect 90982 7590 91012 7642
rect 91036 7590 91046 7642
rect 91046 7590 91092 7642
rect 91116 7590 91162 7642
rect 91162 7590 91172 7642
rect 91196 7590 91226 7642
rect 91226 7590 91252 7642
rect 90956 7588 91012 7590
rect 91036 7588 91092 7590
rect 91116 7588 91172 7590
rect 91196 7588 91252 7590
rect 90956 6554 91012 6556
rect 91036 6554 91092 6556
rect 91116 6554 91172 6556
rect 91196 6554 91252 6556
rect 90956 6502 90982 6554
rect 90982 6502 91012 6554
rect 91036 6502 91046 6554
rect 91046 6502 91092 6554
rect 91116 6502 91162 6554
rect 91162 6502 91172 6554
rect 91196 6502 91226 6554
rect 91226 6502 91252 6554
rect 90956 6500 91012 6502
rect 91036 6500 91092 6502
rect 91116 6500 91172 6502
rect 91196 6500 91252 6502
rect 88062 5616 88118 5672
rect 87970 5072 88026 5128
rect 90956 5466 91012 5468
rect 91036 5466 91092 5468
rect 91116 5466 91172 5468
rect 91196 5466 91252 5468
rect 90956 5414 90982 5466
rect 90982 5414 91012 5466
rect 91036 5414 91046 5466
rect 91046 5414 91092 5466
rect 91116 5414 91162 5466
rect 91162 5414 91172 5466
rect 91196 5414 91226 5466
rect 91226 5414 91252 5466
rect 90956 5412 91012 5414
rect 91036 5412 91092 5414
rect 91116 5412 91172 5414
rect 91196 5412 91252 5414
rect 88154 4936 88210 4992
rect 89810 4936 89866 4992
rect 88706 4800 88762 4856
rect 80702 3984 80758 4040
rect 86958 3984 87014 4040
rect 67454 2896 67510 2952
rect 73342 2896 73398 2952
rect 88706 3848 88762 3904
rect 43902 2488 43958 2544
rect 39486 1264 39542 1320
rect 54956 2202 55012 2204
rect 55036 2202 55092 2204
rect 55116 2202 55172 2204
rect 55196 2202 55252 2204
rect 54956 2150 54982 2202
rect 54982 2150 55012 2202
rect 55036 2150 55046 2202
rect 55046 2150 55092 2202
rect 55116 2150 55162 2202
rect 55162 2150 55172 2202
rect 55196 2150 55226 2202
rect 55226 2150 55252 2202
rect 54956 2148 55012 2150
rect 55036 2148 55092 2150
rect 55116 2148 55172 2150
rect 55196 2148 55252 2150
rect 50250 1264 50306 1320
rect 53470 1264 53526 1320
rect 67362 2352 67418 2408
rect 64142 1264 64198 1320
rect 72956 2746 73012 2748
rect 73036 2746 73092 2748
rect 73116 2746 73172 2748
rect 73196 2746 73252 2748
rect 72956 2694 72982 2746
rect 72982 2694 73012 2746
rect 73036 2694 73046 2746
rect 73046 2694 73092 2746
rect 73116 2694 73162 2746
rect 73162 2694 73172 2746
rect 73196 2694 73226 2746
rect 73226 2694 73252 2746
rect 72956 2692 73012 2694
rect 73036 2692 73092 2694
rect 73116 2692 73172 2694
rect 73196 2692 73252 2694
rect 80242 2624 80298 2680
rect 77298 2352 77354 2408
rect 88890 3440 88946 3496
rect 88246 2352 88302 2408
rect 88706 1400 88762 1456
rect 90956 4378 91012 4380
rect 91036 4378 91092 4380
rect 91116 4378 91172 4380
rect 91196 4378 91252 4380
rect 90956 4326 90982 4378
rect 90982 4326 91012 4378
rect 91036 4326 91046 4378
rect 91046 4326 91092 4378
rect 91116 4326 91162 4378
rect 91162 4326 91172 4378
rect 91196 4326 91226 4378
rect 91226 4326 91252 4378
rect 90956 4324 91012 4326
rect 91036 4324 91092 4326
rect 91116 4324 91172 4326
rect 91196 4324 91252 4326
rect 104162 12688 104218 12744
rect 107474 10376 107530 10432
rect 107290 8064 107346 8120
rect 107474 6160 107530 6216
rect 107290 5072 107346 5128
rect 104162 4800 104218 4856
rect 100758 3440 100814 3496
rect 90956 3290 91012 3292
rect 91036 3290 91092 3292
rect 91116 3290 91172 3292
rect 91196 3290 91252 3292
rect 90956 3238 90982 3290
rect 90982 3238 91012 3290
rect 91036 3238 91046 3290
rect 91046 3238 91092 3290
rect 91116 3238 91162 3290
rect 91162 3238 91172 3290
rect 91196 3238 91226 3290
rect 91226 3238 91252 3290
rect 90956 3236 91012 3238
rect 91036 3236 91092 3238
rect 91116 3236 91172 3238
rect 91196 3236 91252 3238
rect 90730 2624 90786 2680
rect 89810 40 89866 96
rect 104622 2352 104678 2408
rect 90956 2202 91012 2204
rect 91036 2202 91092 2204
rect 91116 2202 91172 2204
rect 91196 2202 91252 2204
rect 90956 2150 90982 2202
rect 90982 2150 91012 2202
rect 91036 2150 91046 2202
rect 91046 2150 91092 2202
rect 91116 2150 91162 2202
rect 91162 2150 91172 2202
rect 91196 2150 91226 2202
rect 91226 2150 91252 2202
rect 90956 2148 91012 2150
rect 91036 2148 91092 2150
rect 91116 2148 91172 2150
rect 91196 2148 91252 2150
rect 97538 1400 97594 1456
rect 105542 1128 105598 1184
rect 105542 40 105598 96
<< metal3 >>
rect 104157 12746 104223 12749
rect 107520 12746 108000 12776
rect 104157 12744 108000 12746
rect 104157 12688 104162 12744
rect 104218 12688 108000 12744
rect 104157 12686 108000 12688
rect 104157 12683 104223 12686
rect 107520 12656 108000 12686
rect 36944 11456 37264 11457
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 11391 37264 11392
rect 72944 11456 73264 11457
rect 72944 11392 72952 11456
rect 73016 11392 73032 11456
rect 73096 11392 73112 11456
rect 73176 11392 73192 11456
rect 73256 11392 73264 11456
rect 72944 11391 73264 11392
rect 18944 10912 19264 10913
rect 18944 10848 18952 10912
rect 19016 10848 19032 10912
rect 19096 10848 19112 10912
rect 19176 10848 19192 10912
rect 19256 10848 19264 10912
rect 18944 10847 19264 10848
rect 54944 10912 55264 10913
rect 54944 10848 54952 10912
rect 55016 10848 55032 10912
rect 55096 10848 55112 10912
rect 55176 10848 55192 10912
rect 55256 10848 55264 10912
rect 54944 10847 55264 10848
rect 90944 10912 91264 10913
rect 90944 10848 90952 10912
rect 91016 10848 91032 10912
rect 91096 10848 91112 10912
rect 91176 10848 91192 10912
rect 91256 10848 91264 10912
rect 90944 10847 91264 10848
rect 107520 10437 108000 10464
rect 107469 10434 108000 10437
rect 107388 10432 108000 10434
rect 107388 10376 107474 10432
rect 107530 10376 108000 10432
rect 107388 10374 108000 10376
rect 107469 10371 108000 10374
rect 36944 10368 37264 10369
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 10303 37264 10304
rect 72944 10368 73264 10369
rect 72944 10304 72952 10368
rect 73016 10304 73032 10368
rect 73096 10304 73112 10368
rect 73176 10304 73192 10368
rect 73256 10304 73264 10368
rect 107520 10344 108000 10371
rect 72944 10303 73264 10304
rect 18944 9824 19264 9825
rect 18944 9760 18952 9824
rect 19016 9760 19032 9824
rect 19096 9760 19112 9824
rect 19176 9760 19192 9824
rect 19256 9760 19264 9824
rect 18944 9759 19264 9760
rect 54944 9824 55264 9825
rect 54944 9760 54952 9824
rect 55016 9760 55032 9824
rect 55096 9760 55112 9824
rect 55176 9760 55192 9824
rect 55256 9760 55264 9824
rect 54944 9759 55264 9760
rect 90944 9824 91264 9825
rect 90944 9760 90952 9824
rect 91016 9760 91032 9824
rect 91096 9760 91112 9824
rect 91176 9760 91192 9824
rect 91256 9760 91264 9824
rect 90944 9759 91264 9760
rect 36944 9280 37264 9281
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 9215 37264 9216
rect 72944 9280 73264 9281
rect 72944 9216 72952 9280
rect 73016 9216 73032 9280
rect 73096 9216 73112 9280
rect 73176 9216 73192 9280
rect 73256 9216 73264 9280
rect 72944 9215 73264 9216
rect 18944 8736 19264 8737
rect 18944 8672 18952 8736
rect 19016 8672 19032 8736
rect 19096 8672 19112 8736
rect 19176 8672 19192 8736
rect 19256 8672 19264 8736
rect 18944 8671 19264 8672
rect 54944 8736 55264 8737
rect 54944 8672 54952 8736
rect 55016 8672 55032 8736
rect 55096 8672 55112 8736
rect 55176 8672 55192 8736
rect 55256 8672 55264 8736
rect 54944 8671 55264 8672
rect 90944 8736 91264 8737
rect 90944 8672 90952 8736
rect 91016 8672 91032 8736
rect 91096 8672 91112 8736
rect 91176 8672 91192 8736
rect 91256 8672 91264 8736
rect 90944 8671 91264 8672
rect 36944 8192 37264 8193
rect 36944 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37264 8192
rect 36944 8127 37264 8128
rect 72944 8192 73264 8193
rect 72944 8128 72952 8192
rect 73016 8128 73032 8192
rect 73096 8128 73112 8192
rect 73176 8128 73192 8192
rect 73256 8128 73264 8192
rect 72944 8127 73264 8128
rect 107285 8122 107351 8125
rect 107520 8122 108000 8152
rect 107285 8120 108000 8122
rect 107285 8064 107290 8120
rect 107346 8064 108000 8120
rect 107285 8062 108000 8064
rect 107285 8059 107351 8062
rect 107520 8032 108000 8062
rect 18944 7648 19264 7649
rect 18944 7584 18952 7648
rect 19016 7584 19032 7648
rect 19096 7584 19112 7648
rect 19176 7584 19192 7648
rect 19256 7584 19264 7648
rect 18944 7583 19264 7584
rect 54944 7648 55264 7649
rect 54944 7584 54952 7648
rect 55016 7584 55032 7648
rect 55096 7584 55112 7648
rect 55176 7584 55192 7648
rect 55256 7584 55264 7648
rect 54944 7583 55264 7584
rect 90944 7648 91264 7649
rect 90944 7584 90952 7648
rect 91016 7584 91032 7648
rect 91096 7584 91112 7648
rect 91176 7584 91192 7648
rect 91256 7584 91264 7648
rect 90944 7583 91264 7584
rect 36944 7104 37264 7105
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 7039 37264 7040
rect 72944 7104 73264 7105
rect 72944 7040 72952 7104
rect 73016 7040 73032 7104
rect 73096 7040 73112 7104
rect 73176 7040 73192 7104
rect 73256 7040 73264 7104
rect 72944 7039 73264 7040
rect 18944 6560 19264 6561
rect 18944 6496 18952 6560
rect 19016 6496 19032 6560
rect 19096 6496 19112 6560
rect 19176 6496 19192 6560
rect 19256 6496 19264 6560
rect 18944 6495 19264 6496
rect 54944 6560 55264 6561
rect 54944 6496 54952 6560
rect 55016 6496 55032 6560
rect 55096 6496 55112 6560
rect 55176 6496 55192 6560
rect 55256 6496 55264 6560
rect 54944 6495 55264 6496
rect 90944 6560 91264 6561
rect 90944 6496 90952 6560
rect 91016 6496 91032 6560
rect 91096 6496 91112 6560
rect 91176 6496 91192 6560
rect 91256 6496 91264 6560
rect 90944 6495 91264 6496
rect 38561 6354 38627 6357
rect 77753 6354 77819 6357
rect 38561 6352 62130 6354
rect 38561 6296 38566 6352
rect 38622 6296 62130 6352
rect 38561 6294 62130 6296
rect 38561 6291 38627 6294
rect 62070 6218 62130 6294
rect 77753 6352 81450 6354
rect 77753 6296 77758 6352
rect 77814 6296 81450 6352
rect 77753 6294 81450 6296
rect 77753 6291 77819 6294
rect 77477 6218 77543 6221
rect 62070 6216 77543 6218
rect 62070 6160 77482 6216
rect 77538 6160 77543 6216
rect 62070 6158 77543 6160
rect 81390 6218 81450 6294
rect 107469 6218 107535 6221
rect 81390 6216 107535 6218
rect 81390 6160 107474 6216
rect 107530 6160 107535 6216
rect 81390 6158 107535 6160
rect 77477 6155 77543 6158
rect 107469 6155 107535 6158
rect 36944 6016 37264 6017
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 5951 37264 5952
rect 72944 6016 73264 6017
rect 72944 5952 72952 6016
rect 73016 5952 73032 6016
rect 73096 5952 73112 6016
rect 73176 5952 73192 6016
rect 73256 5952 73264 6016
rect 72944 5951 73264 5952
rect 51809 5946 51875 5949
rect 59813 5946 59879 5949
rect 51809 5944 59879 5946
rect 51809 5888 51814 5944
rect 51870 5888 59818 5944
rect 59874 5888 59879 5944
rect 51809 5886 59879 5888
rect 51809 5883 51875 5886
rect 59813 5883 59879 5886
rect 38101 5810 38167 5813
rect 63217 5810 63283 5813
rect 107520 5810 108000 5840
rect 38101 5808 63283 5810
rect 38101 5752 38106 5808
rect 38162 5752 63222 5808
rect 63278 5752 63283 5808
rect 38101 5750 63283 5752
rect 38101 5747 38167 5750
rect 63217 5747 63283 5750
rect 100710 5750 108000 5810
rect 39113 5674 39179 5677
rect 51809 5674 51875 5677
rect 39113 5672 51875 5674
rect 39113 5616 39118 5672
rect 39174 5616 51814 5672
rect 51870 5616 51875 5672
rect 39113 5614 51875 5616
rect 39113 5611 39179 5614
rect 51809 5611 51875 5614
rect 88057 5674 88123 5677
rect 100710 5674 100770 5750
rect 107520 5720 108000 5750
rect 88057 5672 100770 5674
rect 88057 5616 88062 5672
rect 88118 5616 100770 5672
rect 88057 5614 100770 5616
rect 88057 5611 88123 5614
rect 61009 5538 61075 5541
rect 68737 5538 68803 5541
rect 61009 5536 68803 5538
rect 61009 5480 61014 5536
rect 61070 5480 68742 5536
rect 68798 5480 68803 5536
rect 61009 5478 68803 5480
rect 61009 5475 61075 5478
rect 68737 5475 68803 5478
rect 18944 5472 19264 5473
rect 18944 5408 18952 5472
rect 19016 5408 19032 5472
rect 19096 5408 19112 5472
rect 19176 5408 19192 5472
rect 19256 5408 19264 5472
rect 18944 5407 19264 5408
rect 54944 5472 55264 5473
rect 54944 5408 54952 5472
rect 55016 5408 55032 5472
rect 55096 5408 55112 5472
rect 55176 5408 55192 5472
rect 55256 5408 55264 5472
rect 54944 5407 55264 5408
rect 90944 5472 91264 5473
rect 90944 5408 90952 5472
rect 91016 5408 91032 5472
rect 91096 5408 91112 5472
rect 91176 5408 91192 5472
rect 91256 5408 91264 5472
rect 90944 5407 91264 5408
rect 4521 5266 4587 5269
rect 37641 5266 37707 5269
rect 4521 5264 37707 5266
rect 4521 5208 4526 5264
rect 4582 5208 37646 5264
rect 37702 5208 37707 5264
rect 4521 5206 37707 5208
rect 4521 5203 4587 5206
rect 37641 5203 37707 5206
rect 39757 5266 39823 5269
rect 60181 5266 60247 5269
rect 39757 5264 60247 5266
rect 39757 5208 39762 5264
rect 39818 5208 60186 5264
rect 60242 5208 60247 5264
rect 39757 5206 60247 5208
rect 39757 5203 39823 5206
rect 60181 5203 60247 5206
rect 18045 5130 18111 5133
rect 37825 5130 37891 5133
rect 18045 5128 37891 5130
rect 18045 5072 18050 5128
rect 18106 5072 37830 5128
rect 37886 5072 37891 5128
rect 18045 5070 37891 5072
rect 18045 5067 18111 5070
rect 37825 5067 37891 5070
rect 51165 5130 51231 5133
rect 62757 5130 62823 5133
rect 77385 5130 77451 5133
rect 87965 5130 88031 5133
rect 107285 5130 107351 5133
rect 51165 5128 62130 5130
rect 51165 5072 51170 5128
rect 51226 5072 62130 5128
rect 51165 5070 62130 5072
rect 51165 5067 51231 5070
rect 62070 4994 62130 5070
rect 62757 5128 81450 5130
rect 62757 5072 62762 5128
rect 62818 5072 77390 5128
rect 77446 5072 81450 5128
rect 62757 5070 81450 5072
rect 62757 5067 62823 5070
rect 77385 5067 77451 5070
rect 72785 4994 72851 4997
rect 62070 4992 72851 4994
rect 62070 4936 72790 4992
rect 72846 4936 72851 4992
rect 62070 4934 72851 4936
rect 81390 4994 81450 5070
rect 87965 5128 107351 5130
rect 87965 5072 87970 5128
rect 88026 5072 107290 5128
rect 107346 5072 107351 5128
rect 87965 5070 107351 5072
rect 87965 5067 88031 5070
rect 107285 5067 107351 5070
rect 88149 4994 88215 4997
rect 89805 4994 89871 4997
rect 81390 4992 89871 4994
rect 81390 4936 88154 4992
rect 88210 4936 89810 4992
rect 89866 4936 89871 4992
rect 81390 4934 89871 4936
rect 72785 4931 72851 4934
rect 88149 4931 88215 4934
rect 89805 4931 89871 4934
rect 36944 4928 37264 4929
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 4863 37264 4864
rect 72944 4928 73264 4929
rect 72944 4864 72952 4928
rect 73016 4864 73032 4928
rect 73096 4864 73112 4928
rect 73176 4864 73192 4928
rect 73256 4864 73264 4928
rect 72944 4863 73264 4864
rect 38469 4858 38535 4861
rect 49877 4858 49943 4861
rect 38469 4856 49943 4858
rect 38469 4800 38474 4856
rect 38530 4800 49882 4856
rect 49938 4800 49943 4856
rect 38469 4798 49943 4800
rect 38469 4795 38535 4798
rect 49877 4795 49943 4798
rect 88701 4858 88767 4861
rect 104157 4858 104223 4861
rect 88701 4856 104223 4858
rect 88701 4800 88706 4856
rect 88762 4800 104162 4856
rect 104218 4800 104223 4856
rect 88701 4798 104223 4800
rect 88701 4795 88767 4798
rect 104157 4795 104223 4798
rect 39205 4722 39271 4725
rect 51165 4722 51231 4725
rect 39205 4720 51231 4722
rect 39205 4664 39210 4720
rect 39266 4664 51170 4720
rect 51226 4664 51231 4720
rect 39205 4662 51231 4664
rect 39205 4659 39271 4662
rect 51165 4659 51231 4662
rect 68829 4722 68895 4725
rect 77845 4722 77911 4725
rect 68829 4720 77911 4722
rect 68829 4664 68834 4720
rect 68890 4664 77850 4720
rect 77906 4664 77911 4720
rect 68829 4662 77911 4664
rect 68829 4659 68895 4662
rect 77845 4659 77911 4662
rect 18944 4384 19264 4385
rect 18944 4320 18952 4384
rect 19016 4320 19032 4384
rect 19096 4320 19112 4384
rect 19176 4320 19192 4384
rect 19256 4320 19264 4384
rect 18944 4319 19264 4320
rect 54944 4384 55264 4385
rect 54944 4320 54952 4384
rect 55016 4320 55032 4384
rect 55096 4320 55112 4384
rect 55176 4320 55192 4384
rect 55256 4320 55264 4384
rect 54944 4319 55264 4320
rect 90944 4384 91264 4385
rect 90944 4320 90952 4384
rect 91016 4320 91032 4384
rect 91096 4320 91112 4384
rect 91176 4320 91192 4384
rect 91256 4320 91264 4384
rect 90944 4319 91264 4320
rect 12433 4042 12499 4045
rect 19333 4042 19399 4045
rect 12433 4040 19399 4042
rect 12433 3984 12438 4040
rect 12494 3984 19338 4040
rect 19394 3984 19399 4040
rect 12433 3982 19399 3984
rect 12433 3979 12499 3982
rect 19333 3979 19399 3982
rect 80697 4042 80763 4045
rect 86953 4042 87019 4045
rect 80697 4040 87019 4042
rect 80697 3984 80702 4040
rect 80758 3984 86958 4040
rect 87014 3984 87019 4040
rect 80697 3982 87019 3984
rect 80697 3979 80763 3982
rect 86953 3979 87019 3982
rect 4889 3906 4955 3909
rect 17769 3906 17835 3909
rect 35249 3906 35315 3909
rect 4889 3904 35315 3906
rect 4889 3848 4894 3904
rect 4950 3848 17774 3904
rect 17830 3848 35254 3904
rect 35310 3848 35315 3904
rect 4889 3846 35315 3848
rect 4889 3843 4955 3846
rect 17769 3843 17835 3846
rect 35249 3843 35315 3846
rect 56869 3906 56935 3909
rect 65793 3906 65859 3909
rect 56869 3904 65859 3906
rect 56869 3848 56874 3904
rect 56930 3848 65798 3904
rect 65854 3848 65859 3904
rect 56869 3846 65859 3848
rect 56869 3843 56935 3846
rect 65793 3843 65859 3846
rect 78949 3906 79015 3909
rect 88701 3906 88767 3909
rect 78949 3904 88767 3906
rect 78949 3848 78954 3904
rect 79010 3848 88706 3904
rect 88762 3848 88767 3904
rect 78949 3846 88767 3848
rect 78949 3843 79015 3846
rect 88701 3843 88767 3846
rect 36944 3840 37264 3841
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 3775 37264 3776
rect 72944 3840 73264 3841
rect 72944 3776 72952 3840
rect 73016 3776 73032 3840
rect 73096 3776 73112 3840
rect 73176 3776 73192 3840
rect 73256 3776 73264 3840
rect 72944 3775 73264 3776
rect 49969 3770 50035 3773
rect 60365 3770 60431 3773
rect 49969 3768 60431 3770
rect 49969 3712 49974 3768
rect 50030 3712 60370 3768
rect 60426 3712 60431 3768
rect 49969 3710 60431 3712
rect 49969 3707 50035 3710
rect 60365 3707 60431 3710
rect 2313 3634 2379 3637
rect 37825 3634 37891 3637
rect 2313 3632 37891 3634
rect 2313 3576 2318 3632
rect 2374 3576 37830 3632
rect 37886 3576 37891 3632
rect 2313 3574 37891 3576
rect 2313 3571 2379 3574
rect 37825 3571 37891 3574
rect 65793 3634 65859 3637
rect 78949 3634 79015 3637
rect 65793 3632 79015 3634
rect 65793 3576 65798 3632
rect 65854 3576 78954 3632
rect 79010 3576 79015 3632
rect 65793 3574 79015 3576
rect 65793 3571 65859 3574
rect 78949 3571 79015 3574
rect 88885 3498 88951 3501
rect 100753 3498 100819 3501
rect 88885 3496 100819 3498
rect 88885 3440 88890 3496
rect 88946 3440 100758 3496
rect 100814 3440 100819 3496
rect 88885 3438 100819 3440
rect 88885 3435 88951 3438
rect 100753 3435 100819 3438
rect 107520 3408 108000 3528
rect 18944 3296 19264 3297
rect 18944 3232 18952 3296
rect 19016 3232 19032 3296
rect 19096 3232 19112 3296
rect 19176 3232 19192 3296
rect 19256 3232 19264 3296
rect 18944 3231 19264 3232
rect 54944 3296 55264 3297
rect 54944 3232 54952 3296
rect 55016 3232 55032 3296
rect 55096 3232 55112 3296
rect 55176 3232 55192 3296
rect 55256 3232 55264 3296
rect 54944 3231 55264 3232
rect 90944 3296 91264 3297
rect 90944 3232 90952 3296
rect 91016 3232 91032 3296
rect 91096 3232 91112 3296
rect 91176 3232 91192 3296
rect 91256 3232 91264 3296
rect 90944 3231 91264 3232
rect 35249 3090 35315 3093
rect 56869 3090 56935 3093
rect 35249 3088 56935 3090
rect 35249 3032 35254 3088
rect 35310 3032 56874 3088
rect 56930 3032 56935 3088
rect 35249 3030 56935 3032
rect 35249 3027 35315 3030
rect 56869 3027 56935 3030
rect 26141 2954 26207 2957
rect 33133 2954 33199 2957
rect 26141 2952 33199 2954
rect 26141 2896 26146 2952
rect 26202 2896 33138 2952
rect 33194 2896 33199 2952
rect 26141 2894 33199 2896
rect 26141 2891 26207 2894
rect 33133 2891 33199 2894
rect 67449 2954 67515 2957
rect 73337 2954 73403 2957
rect 67449 2952 73403 2954
rect 67449 2896 67454 2952
rect 67510 2896 73342 2952
rect 73398 2896 73403 2952
rect 67449 2894 73403 2896
rect 67449 2891 67515 2894
rect 73337 2891 73403 2894
rect 36944 2752 37264 2753
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2687 37264 2688
rect 72944 2752 73264 2753
rect 72944 2688 72952 2752
rect 73016 2688 73032 2752
rect 73096 2688 73112 2752
rect 73176 2688 73192 2752
rect 73256 2688 73264 2752
rect 72944 2687 73264 2688
rect 25681 2682 25747 2685
rect 36629 2682 36695 2685
rect 25681 2680 36695 2682
rect 25681 2624 25686 2680
rect 25742 2624 36634 2680
rect 36690 2624 36695 2680
rect 25681 2622 36695 2624
rect 25681 2619 25747 2622
rect 36629 2619 36695 2622
rect 80237 2682 80303 2685
rect 90725 2682 90791 2685
rect 80237 2680 90791 2682
rect 80237 2624 80242 2680
rect 80298 2624 90730 2680
rect 90786 2624 90791 2680
rect 80237 2622 90791 2624
rect 80237 2619 80303 2622
rect 90725 2619 90791 2622
rect 6821 2546 6887 2549
rect 16849 2546 16915 2549
rect 6821 2544 16915 2546
rect 6821 2488 6826 2544
rect 6882 2488 16854 2544
rect 16910 2488 16915 2544
rect 6821 2486 16915 2488
rect 6821 2483 6887 2486
rect 16849 2483 16915 2486
rect 36169 2546 36235 2549
rect 43897 2546 43963 2549
rect 36169 2544 43963 2546
rect 36169 2488 36174 2544
rect 36230 2488 43902 2544
rect 43958 2488 43963 2544
rect 36169 2486 43963 2488
rect 36169 2483 36235 2486
rect 43897 2483 43963 2486
rect 12617 2410 12683 2413
rect 23657 2410 23723 2413
rect 12617 2408 23723 2410
rect 12617 2352 12622 2408
rect 12678 2352 23662 2408
rect 23718 2352 23723 2408
rect 12617 2350 23723 2352
rect 12617 2347 12683 2350
rect 23657 2347 23723 2350
rect 67357 2410 67423 2413
rect 77293 2410 77359 2413
rect 67357 2408 77359 2410
rect 67357 2352 67362 2408
rect 67418 2352 77298 2408
rect 77354 2352 77359 2408
rect 67357 2350 77359 2352
rect 67357 2347 67423 2350
rect 77293 2347 77359 2350
rect 88241 2410 88307 2413
rect 104617 2410 104683 2413
rect 88241 2408 104683 2410
rect 88241 2352 88246 2408
rect 88302 2352 104622 2408
rect 104678 2352 104683 2408
rect 88241 2350 104683 2352
rect 88241 2347 88307 2350
rect 104617 2347 104683 2350
rect 18944 2208 19264 2209
rect 18944 2144 18952 2208
rect 19016 2144 19032 2208
rect 19096 2144 19112 2208
rect 19176 2144 19192 2208
rect 19256 2144 19264 2208
rect 18944 2143 19264 2144
rect 54944 2208 55264 2209
rect 54944 2144 54952 2208
rect 55016 2144 55032 2208
rect 55096 2144 55112 2208
rect 55176 2144 55192 2208
rect 55256 2144 55264 2208
rect 54944 2143 55264 2144
rect 90944 2208 91264 2209
rect 90944 2144 90952 2208
rect 91016 2144 91032 2208
rect 91096 2144 91112 2208
rect 91176 2144 91192 2208
rect 91256 2144 91264 2208
rect 90944 2143 91264 2144
rect 1577 1458 1643 1461
rect 9765 1458 9831 1461
rect 1577 1456 9831 1458
rect 1577 1400 1582 1456
rect 1638 1400 9770 1456
rect 9826 1400 9831 1456
rect 1577 1398 9831 1400
rect 1577 1395 1643 1398
rect 9765 1395 9831 1398
rect 20621 1458 20687 1461
rect 30005 1458 30071 1461
rect 20621 1456 30071 1458
rect 20621 1400 20626 1456
rect 20682 1400 30010 1456
rect 30066 1400 30071 1456
rect 20621 1398 30071 1400
rect 20621 1395 20687 1398
rect 30005 1395 30071 1398
rect 88701 1458 88767 1461
rect 97533 1458 97599 1461
rect 88701 1456 97599 1458
rect 88701 1400 88706 1456
rect 88762 1400 97538 1456
rect 97594 1400 97599 1456
rect 88701 1398 97599 1400
rect 88701 1395 88767 1398
rect 97533 1395 97599 1398
rect 39481 1322 39547 1325
rect 50245 1322 50311 1325
rect 39481 1320 50311 1322
rect 39481 1264 39486 1320
rect 39542 1264 50250 1320
rect 50306 1264 50311 1320
rect 39481 1262 50311 1264
rect 39481 1259 39547 1262
rect 50245 1259 50311 1262
rect 53465 1322 53531 1325
rect 64137 1322 64203 1325
rect 53465 1320 64203 1322
rect 53465 1264 53470 1320
rect 53526 1264 64142 1320
rect 64198 1264 64203 1320
rect 53465 1262 64203 1264
rect 53465 1259 53531 1262
rect 64137 1259 64203 1262
rect 105537 1186 105603 1189
rect 107520 1186 108000 1216
rect 105537 1184 108000 1186
rect 105537 1128 105542 1184
rect 105598 1128 108000 1184
rect 105537 1126 108000 1128
rect 105537 1123 105603 1126
rect 107520 1096 108000 1126
rect 89805 98 89871 101
rect 105537 98 105603 101
rect 89805 96 105603 98
rect 89805 40 89810 96
rect 89866 40 105542 96
rect 105598 40 105603 96
rect 89805 38 105603 40
rect 89805 35 89871 38
rect 105537 35 105603 38
<< via3 >>
rect 36952 11452 37016 11456
rect 36952 11396 36956 11452
rect 36956 11396 37012 11452
rect 37012 11396 37016 11452
rect 36952 11392 37016 11396
rect 37032 11452 37096 11456
rect 37032 11396 37036 11452
rect 37036 11396 37092 11452
rect 37092 11396 37096 11452
rect 37032 11392 37096 11396
rect 37112 11452 37176 11456
rect 37112 11396 37116 11452
rect 37116 11396 37172 11452
rect 37172 11396 37176 11452
rect 37112 11392 37176 11396
rect 37192 11452 37256 11456
rect 37192 11396 37196 11452
rect 37196 11396 37252 11452
rect 37252 11396 37256 11452
rect 37192 11392 37256 11396
rect 72952 11452 73016 11456
rect 72952 11396 72956 11452
rect 72956 11396 73012 11452
rect 73012 11396 73016 11452
rect 72952 11392 73016 11396
rect 73032 11452 73096 11456
rect 73032 11396 73036 11452
rect 73036 11396 73092 11452
rect 73092 11396 73096 11452
rect 73032 11392 73096 11396
rect 73112 11452 73176 11456
rect 73112 11396 73116 11452
rect 73116 11396 73172 11452
rect 73172 11396 73176 11452
rect 73112 11392 73176 11396
rect 73192 11452 73256 11456
rect 73192 11396 73196 11452
rect 73196 11396 73252 11452
rect 73252 11396 73256 11452
rect 73192 11392 73256 11396
rect 18952 10908 19016 10912
rect 18952 10852 18956 10908
rect 18956 10852 19012 10908
rect 19012 10852 19016 10908
rect 18952 10848 19016 10852
rect 19032 10908 19096 10912
rect 19032 10852 19036 10908
rect 19036 10852 19092 10908
rect 19092 10852 19096 10908
rect 19032 10848 19096 10852
rect 19112 10908 19176 10912
rect 19112 10852 19116 10908
rect 19116 10852 19172 10908
rect 19172 10852 19176 10908
rect 19112 10848 19176 10852
rect 19192 10908 19256 10912
rect 19192 10852 19196 10908
rect 19196 10852 19252 10908
rect 19252 10852 19256 10908
rect 19192 10848 19256 10852
rect 54952 10908 55016 10912
rect 54952 10852 54956 10908
rect 54956 10852 55012 10908
rect 55012 10852 55016 10908
rect 54952 10848 55016 10852
rect 55032 10908 55096 10912
rect 55032 10852 55036 10908
rect 55036 10852 55092 10908
rect 55092 10852 55096 10908
rect 55032 10848 55096 10852
rect 55112 10908 55176 10912
rect 55112 10852 55116 10908
rect 55116 10852 55172 10908
rect 55172 10852 55176 10908
rect 55112 10848 55176 10852
rect 55192 10908 55256 10912
rect 55192 10852 55196 10908
rect 55196 10852 55252 10908
rect 55252 10852 55256 10908
rect 55192 10848 55256 10852
rect 90952 10908 91016 10912
rect 90952 10852 90956 10908
rect 90956 10852 91012 10908
rect 91012 10852 91016 10908
rect 90952 10848 91016 10852
rect 91032 10908 91096 10912
rect 91032 10852 91036 10908
rect 91036 10852 91092 10908
rect 91092 10852 91096 10908
rect 91032 10848 91096 10852
rect 91112 10908 91176 10912
rect 91112 10852 91116 10908
rect 91116 10852 91172 10908
rect 91172 10852 91176 10908
rect 91112 10848 91176 10852
rect 91192 10908 91256 10912
rect 91192 10852 91196 10908
rect 91196 10852 91252 10908
rect 91252 10852 91256 10908
rect 91192 10848 91256 10852
rect 36952 10364 37016 10368
rect 36952 10308 36956 10364
rect 36956 10308 37012 10364
rect 37012 10308 37016 10364
rect 36952 10304 37016 10308
rect 37032 10364 37096 10368
rect 37032 10308 37036 10364
rect 37036 10308 37092 10364
rect 37092 10308 37096 10364
rect 37032 10304 37096 10308
rect 37112 10364 37176 10368
rect 37112 10308 37116 10364
rect 37116 10308 37172 10364
rect 37172 10308 37176 10364
rect 37112 10304 37176 10308
rect 37192 10364 37256 10368
rect 37192 10308 37196 10364
rect 37196 10308 37252 10364
rect 37252 10308 37256 10364
rect 37192 10304 37256 10308
rect 72952 10364 73016 10368
rect 72952 10308 72956 10364
rect 72956 10308 73012 10364
rect 73012 10308 73016 10364
rect 72952 10304 73016 10308
rect 73032 10364 73096 10368
rect 73032 10308 73036 10364
rect 73036 10308 73092 10364
rect 73092 10308 73096 10364
rect 73032 10304 73096 10308
rect 73112 10364 73176 10368
rect 73112 10308 73116 10364
rect 73116 10308 73172 10364
rect 73172 10308 73176 10364
rect 73112 10304 73176 10308
rect 73192 10364 73256 10368
rect 73192 10308 73196 10364
rect 73196 10308 73252 10364
rect 73252 10308 73256 10364
rect 73192 10304 73256 10308
rect 18952 9820 19016 9824
rect 18952 9764 18956 9820
rect 18956 9764 19012 9820
rect 19012 9764 19016 9820
rect 18952 9760 19016 9764
rect 19032 9820 19096 9824
rect 19032 9764 19036 9820
rect 19036 9764 19092 9820
rect 19092 9764 19096 9820
rect 19032 9760 19096 9764
rect 19112 9820 19176 9824
rect 19112 9764 19116 9820
rect 19116 9764 19172 9820
rect 19172 9764 19176 9820
rect 19112 9760 19176 9764
rect 19192 9820 19256 9824
rect 19192 9764 19196 9820
rect 19196 9764 19252 9820
rect 19252 9764 19256 9820
rect 19192 9760 19256 9764
rect 54952 9820 55016 9824
rect 54952 9764 54956 9820
rect 54956 9764 55012 9820
rect 55012 9764 55016 9820
rect 54952 9760 55016 9764
rect 55032 9820 55096 9824
rect 55032 9764 55036 9820
rect 55036 9764 55092 9820
rect 55092 9764 55096 9820
rect 55032 9760 55096 9764
rect 55112 9820 55176 9824
rect 55112 9764 55116 9820
rect 55116 9764 55172 9820
rect 55172 9764 55176 9820
rect 55112 9760 55176 9764
rect 55192 9820 55256 9824
rect 55192 9764 55196 9820
rect 55196 9764 55252 9820
rect 55252 9764 55256 9820
rect 55192 9760 55256 9764
rect 90952 9820 91016 9824
rect 90952 9764 90956 9820
rect 90956 9764 91012 9820
rect 91012 9764 91016 9820
rect 90952 9760 91016 9764
rect 91032 9820 91096 9824
rect 91032 9764 91036 9820
rect 91036 9764 91092 9820
rect 91092 9764 91096 9820
rect 91032 9760 91096 9764
rect 91112 9820 91176 9824
rect 91112 9764 91116 9820
rect 91116 9764 91172 9820
rect 91172 9764 91176 9820
rect 91112 9760 91176 9764
rect 91192 9820 91256 9824
rect 91192 9764 91196 9820
rect 91196 9764 91252 9820
rect 91252 9764 91256 9820
rect 91192 9760 91256 9764
rect 36952 9276 37016 9280
rect 36952 9220 36956 9276
rect 36956 9220 37012 9276
rect 37012 9220 37016 9276
rect 36952 9216 37016 9220
rect 37032 9276 37096 9280
rect 37032 9220 37036 9276
rect 37036 9220 37092 9276
rect 37092 9220 37096 9276
rect 37032 9216 37096 9220
rect 37112 9276 37176 9280
rect 37112 9220 37116 9276
rect 37116 9220 37172 9276
rect 37172 9220 37176 9276
rect 37112 9216 37176 9220
rect 37192 9276 37256 9280
rect 37192 9220 37196 9276
rect 37196 9220 37252 9276
rect 37252 9220 37256 9276
rect 37192 9216 37256 9220
rect 72952 9276 73016 9280
rect 72952 9220 72956 9276
rect 72956 9220 73012 9276
rect 73012 9220 73016 9276
rect 72952 9216 73016 9220
rect 73032 9276 73096 9280
rect 73032 9220 73036 9276
rect 73036 9220 73092 9276
rect 73092 9220 73096 9276
rect 73032 9216 73096 9220
rect 73112 9276 73176 9280
rect 73112 9220 73116 9276
rect 73116 9220 73172 9276
rect 73172 9220 73176 9276
rect 73112 9216 73176 9220
rect 73192 9276 73256 9280
rect 73192 9220 73196 9276
rect 73196 9220 73252 9276
rect 73252 9220 73256 9276
rect 73192 9216 73256 9220
rect 18952 8732 19016 8736
rect 18952 8676 18956 8732
rect 18956 8676 19012 8732
rect 19012 8676 19016 8732
rect 18952 8672 19016 8676
rect 19032 8732 19096 8736
rect 19032 8676 19036 8732
rect 19036 8676 19092 8732
rect 19092 8676 19096 8732
rect 19032 8672 19096 8676
rect 19112 8732 19176 8736
rect 19112 8676 19116 8732
rect 19116 8676 19172 8732
rect 19172 8676 19176 8732
rect 19112 8672 19176 8676
rect 19192 8732 19256 8736
rect 19192 8676 19196 8732
rect 19196 8676 19252 8732
rect 19252 8676 19256 8732
rect 19192 8672 19256 8676
rect 54952 8732 55016 8736
rect 54952 8676 54956 8732
rect 54956 8676 55012 8732
rect 55012 8676 55016 8732
rect 54952 8672 55016 8676
rect 55032 8732 55096 8736
rect 55032 8676 55036 8732
rect 55036 8676 55092 8732
rect 55092 8676 55096 8732
rect 55032 8672 55096 8676
rect 55112 8732 55176 8736
rect 55112 8676 55116 8732
rect 55116 8676 55172 8732
rect 55172 8676 55176 8732
rect 55112 8672 55176 8676
rect 55192 8732 55256 8736
rect 55192 8676 55196 8732
rect 55196 8676 55252 8732
rect 55252 8676 55256 8732
rect 55192 8672 55256 8676
rect 90952 8732 91016 8736
rect 90952 8676 90956 8732
rect 90956 8676 91012 8732
rect 91012 8676 91016 8732
rect 90952 8672 91016 8676
rect 91032 8732 91096 8736
rect 91032 8676 91036 8732
rect 91036 8676 91092 8732
rect 91092 8676 91096 8732
rect 91032 8672 91096 8676
rect 91112 8732 91176 8736
rect 91112 8676 91116 8732
rect 91116 8676 91172 8732
rect 91172 8676 91176 8732
rect 91112 8672 91176 8676
rect 91192 8732 91256 8736
rect 91192 8676 91196 8732
rect 91196 8676 91252 8732
rect 91252 8676 91256 8732
rect 91192 8672 91256 8676
rect 36952 8188 37016 8192
rect 36952 8132 36956 8188
rect 36956 8132 37012 8188
rect 37012 8132 37016 8188
rect 36952 8128 37016 8132
rect 37032 8188 37096 8192
rect 37032 8132 37036 8188
rect 37036 8132 37092 8188
rect 37092 8132 37096 8188
rect 37032 8128 37096 8132
rect 37112 8188 37176 8192
rect 37112 8132 37116 8188
rect 37116 8132 37172 8188
rect 37172 8132 37176 8188
rect 37112 8128 37176 8132
rect 37192 8188 37256 8192
rect 37192 8132 37196 8188
rect 37196 8132 37252 8188
rect 37252 8132 37256 8188
rect 37192 8128 37256 8132
rect 72952 8188 73016 8192
rect 72952 8132 72956 8188
rect 72956 8132 73012 8188
rect 73012 8132 73016 8188
rect 72952 8128 73016 8132
rect 73032 8188 73096 8192
rect 73032 8132 73036 8188
rect 73036 8132 73092 8188
rect 73092 8132 73096 8188
rect 73032 8128 73096 8132
rect 73112 8188 73176 8192
rect 73112 8132 73116 8188
rect 73116 8132 73172 8188
rect 73172 8132 73176 8188
rect 73112 8128 73176 8132
rect 73192 8188 73256 8192
rect 73192 8132 73196 8188
rect 73196 8132 73252 8188
rect 73252 8132 73256 8188
rect 73192 8128 73256 8132
rect 18952 7644 19016 7648
rect 18952 7588 18956 7644
rect 18956 7588 19012 7644
rect 19012 7588 19016 7644
rect 18952 7584 19016 7588
rect 19032 7644 19096 7648
rect 19032 7588 19036 7644
rect 19036 7588 19092 7644
rect 19092 7588 19096 7644
rect 19032 7584 19096 7588
rect 19112 7644 19176 7648
rect 19112 7588 19116 7644
rect 19116 7588 19172 7644
rect 19172 7588 19176 7644
rect 19112 7584 19176 7588
rect 19192 7644 19256 7648
rect 19192 7588 19196 7644
rect 19196 7588 19252 7644
rect 19252 7588 19256 7644
rect 19192 7584 19256 7588
rect 54952 7644 55016 7648
rect 54952 7588 54956 7644
rect 54956 7588 55012 7644
rect 55012 7588 55016 7644
rect 54952 7584 55016 7588
rect 55032 7644 55096 7648
rect 55032 7588 55036 7644
rect 55036 7588 55092 7644
rect 55092 7588 55096 7644
rect 55032 7584 55096 7588
rect 55112 7644 55176 7648
rect 55112 7588 55116 7644
rect 55116 7588 55172 7644
rect 55172 7588 55176 7644
rect 55112 7584 55176 7588
rect 55192 7644 55256 7648
rect 55192 7588 55196 7644
rect 55196 7588 55252 7644
rect 55252 7588 55256 7644
rect 55192 7584 55256 7588
rect 90952 7644 91016 7648
rect 90952 7588 90956 7644
rect 90956 7588 91012 7644
rect 91012 7588 91016 7644
rect 90952 7584 91016 7588
rect 91032 7644 91096 7648
rect 91032 7588 91036 7644
rect 91036 7588 91092 7644
rect 91092 7588 91096 7644
rect 91032 7584 91096 7588
rect 91112 7644 91176 7648
rect 91112 7588 91116 7644
rect 91116 7588 91172 7644
rect 91172 7588 91176 7644
rect 91112 7584 91176 7588
rect 91192 7644 91256 7648
rect 91192 7588 91196 7644
rect 91196 7588 91252 7644
rect 91252 7588 91256 7644
rect 91192 7584 91256 7588
rect 36952 7100 37016 7104
rect 36952 7044 36956 7100
rect 36956 7044 37012 7100
rect 37012 7044 37016 7100
rect 36952 7040 37016 7044
rect 37032 7100 37096 7104
rect 37032 7044 37036 7100
rect 37036 7044 37092 7100
rect 37092 7044 37096 7100
rect 37032 7040 37096 7044
rect 37112 7100 37176 7104
rect 37112 7044 37116 7100
rect 37116 7044 37172 7100
rect 37172 7044 37176 7100
rect 37112 7040 37176 7044
rect 37192 7100 37256 7104
rect 37192 7044 37196 7100
rect 37196 7044 37252 7100
rect 37252 7044 37256 7100
rect 37192 7040 37256 7044
rect 72952 7100 73016 7104
rect 72952 7044 72956 7100
rect 72956 7044 73012 7100
rect 73012 7044 73016 7100
rect 72952 7040 73016 7044
rect 73032 7100 73096 7104
rect 73032 7044 73036 7100
rect 73036 7044 73092 7100
rect 73092 7044 73096 7100
rect 73032 7040 73096 7044
rect 73112 7100 73176 7104
rect 73112 7044 73116 7100
rect 73116 7044 73172 7100
rect 73172 7044 73176 7100
rect 73112 7040 73176 7044
rect 73192 7100 73256 7104
rect 73192 7044 73196 7100
rect 73196 7044 73252 7100
rect 73252 7044 73256 7100
rect 73192 7040 73256 7044
rect 18952 6556 19016 6560
rect 18952 6500 18956 6556
rect 18956 6500 19012 6556
rect 19012 6500 19016 6556
rect 18952 6496 19016 6500
rect 19032 6556 19096 6560
rect 19032 6500 19036 6556
rect 19036 6500 19092 6556
rect 19092 6500 19096 6556
rect 19032 6496 19096 6500
rect 19112 6556 19176 6560
rect 19112 6500 19116 6556
rect 19116 6500 19172 6556
rect 19172 6500 19176 6556
rect 19112 6496 19176 6500
rect 19192 6556 19256 6560
rect 19192 6500 19196 6556
rect 19196 6500 19252 6556
rect 19252 6500 19256 6556
rect 19192 6496 19256 6500
rect 54952 6556 55016 6560
rect 54952 6500 54956 6556
rect 54956 6500 55012 6556
rect 55012 6500 55016 6556
rect 54952 6496 55016 6500
rect 55032 6556 55096 6560
rect 55032 6500 55036 6556
rect 55036 6500 55092 6556
rect 55092 6500 55096 6556
rect 55032 6496 55096 6500
rect 55112 6556 55176 6560
rect 55112 6500 55116 6556
rect 55116 6500 55172 6556
rect 55172 6500 55176 6556
rect 55112 6496 55176 6500
rect 55192 6556 55256 6560
rect 55192 6500 55196 6556
rect 55196 6500 55252 6556
rect 55252 6500 55256 6556
rect 55192 6496 55256 6500
rect 90952 6556 91016 6560
rect 90952 6500 90956 6556
rect 90956 6500 91012 6556
rect 91012 6500 91016 6556
rect 90952 6496 91016 6500
rect 91032 6556 91096 6560
rect 91032 6500 91036 6556
rect 91036 6500 91092 6556
rect 91092 6500 91096 6556
rect 91032 6496 91096 6500
rect 91112 6556 91176 6560
rect 91112 6500 91116 6556
rect 91116 6500 91172 6556
rect 91172 6500 91176 6556
rect 91112 6496 91176 6500
rect 91192 6556 91256 6560
rect 91192 6500 91196 6556
rect 91196 6500 91252 6556
rect 91252 6500 91256 6556
rect 91192 6496 91256 6500
rect 36952 6012 37016 6016
rect 36952 5956 36956 6012
rect 36956 5956 37012 6012
rect 37012 5956 37016 6012
rect 36952 5952 37016 5956
rect 37032 6012 37096 6016
rect 37032 5956 37036 6012
rect 37036 5956 37092 6012
rect 37092 5956 37096 6012
rect 37032 5952 37096 5956
rect 37112 6012 37176 6016
rect 37112 5956 37116 6012
rect 37116 5956 37172 6012
rect 37172 5956 37176 6012
rect 37112 5952 37176 5956
rect 37192 6012 37256 6016
rect 37192 5956 37196 6012
rect 37196 5956 37252 6012
rect 37252 5956 37256 6012
rect 37192 5952 37256 5956
rect 72952 6012 73016 6016
rect 72952 5956 72956 6012
rect 72956 5956 73012 6012
rect 73012 5956 73016 6012
rect 72952 5952 73016 5956
rect 73032 6012 73096 6016
rect 73032 5956 73036 6012
rect 73036 5956 73092 6012
rect 73092 5956 73096 6012
rect 73032 5952 73096 5956
rect 73112 6012 73176 6016
rect 73112 5956 73116 6012
rect 73116 5956 73172 6012
rect 73172 5956 73176 6012
rect 73112 5952 73176 5956
rect 73192 6012 73256 6016
rect 73192 5956 73196 6012
rect 73196 5956 73252 6012
rect 73252 5956 73256 6012
rect 73192 5952 73256 5956
rect 18952 5468 19016 5472
rect 18952 5412 18956 5468
rect 18956 5412 19012 5468
rect 19012 5412 19016 5468
rect 18952 5408 19016 5412
rect 19032 5468 19096 5472
rect 19032 5412 19036 5468
rect 19036 5412 19092 5468
rect 19092 5412 19096 5468
rect 19032 5408 19096 5412
rect 19112 5468 19176 5472
rect 19112 5412 19116 5468
rect 19116 5412 19172 5468
rect 19172 5412 19176 5468
rect 19112 5408 19176 5412
rect 19192 5468 19256 5472
rect 19192 5412 19196 5468
rect 19196 5412 19252 5468
rect 19252 5412 19256 5468
rect 19192 5408 19256 5412
rect 54952 5468 55016 5472
rect 54952 5412 54956 5468
rect 54956 5412 55012 5468
rect 55012 5412 55016 5468
rect 54952 5408 55016 5412
rect 55032 5468 55096 5472
rect 55032 5412 55036 5468
rect 55036 5412 55092 5468
rect 55092 5412 55096 5468
rect 55032 5408 55096 5412
rect 55112 5468 55176 5472
rect 55112 5412 55116 5468
rect 55116 5412 55172 5468
rect 55172 5412 55176 5468
rect 55112 5408 55176 5412
rect 55192 5468 55256 5472
rect 55192 5412 55196 5468
rect 55196 5412 55252 5468
rect 55252 5412 55256 5468
rect 55192 5408 55256 5412
rect 90952 5468 91016 5472
rect 90952 5412 90956 5468
rect 90956 5412 91012 5468
rect 91012 5412 91016 5468
rect 90952 5408 91016 5412
rect 91032 5468 91096 5472
rect 91032 5412 91036 5468
rect 91036 5412 91092 5468
rect 91092 5412 91096 5468
rect 91032 5408 91096 5412
rect 91112 5468 91176 5472
rect 91112 5412 91116 5468
rect 91116 5412 91172 5468
rect 91172 5412 91176 5468
rect 91112 5408 91176 5412
rect 91192 5468 91256 5472
rect 91192 5412 91196 5468
rect 91196 5412 91252 5468
rect 91252 5412 91256 5468
rect 91192 5408 91256 5412
rect 36952 4924 37016 4928
rect 36952 4868 36956 4924
rect 36956 4868 37012 4924
rect 37012 4868 37016 4924
rect 36952 4864 37016 4868
rect 37032 4924 37096 4928
rect 37032 4868 37036 4924
rect 37036 4868 37092 4924
rect 37092 4868 37096 4924
rect 37032 4864 37096 4868
rect 37112 4924 37176 4928
rect 37112 4868 37116 4924
rect 37116 4868 37172 4924
rect 37172 4868 37176 4924
rect 37112 4864 37176 4868
rect 37192 4924 37256 4928
rect 37192 4868 37196 4924
rect 37196 4868 37252 4924
rect 37252 4868 37256 4924
rect 37192 4864 37256 4868
rect 72952 4924 73016 4928
rect 72952 4868 72956 4924
rect 72956 4868 73012 4924
rect 73012 4868 73016 4924
rect 72952 4864 73016 4868
rect 73032 4924 73096 4928
rect 73032 4868 73036 4924
rect 73036 4868 73092 4924
rect 73092 4868 73096 4924
rect 73032 4864 73096 4868
rect 73112 4924 73176 4928
rect 73112 4868 73116 4924
rect 73116 4868 73172 4924
rect 73172 4868 73176 4924
rect 73112 4864 73176 4868
rect 73192 4924 73256 4928
rect 73192 4868 73196 4924
rect 73196 4868 73252 4924
rect 73252 4868 73256 4924
rect 73192 4864 73256 4868
rect 18952 4380 19016 4384
rect 18952 4324 18956 4380
rect 18956 4324 19012 4380
rect 19012 4324 19016 4380
rect 18952 4320 19016 4324
rect 19032 4380 19096 4384
rect 19032 4324 19036 4380
rect 19036 4324 19092 4380
rect 19092 4324 19096 4380
rect 19032 4320 19096 4324
rect 19112 4380 19176 4384
rect 19112 4324 19116 4380
rect 19116 4324 19172 4380
rect 19172 4324 19176 4380
rect 19112 4320 19176 4324
rect 19192 4380 19256 4384
rect 19192 4324 19196 4380
rect 19196 4324 19252 4380
rect 19252 4324 19256 4380
rect 19192 4320 19256 4324
rect 54952 4380 55016 4384
rect 54952 4324 54956 4380
rect 54956 4324 55012 4380
rect 55012 4324 55016 4380
rect 54952 4320 55016 4324
rect 55032 4380 55096 4384
rect 55032 4324 55036 4380
rect 55036 4324 55092 4380
rect 55092 4324 55096 4380
rect 55032 4320 55096 4324
rect 55112 4380 55176 4384
rect 55112 4324 55116 4380
rect 55116 4324 55172 4380
rect 55172 4324 55176 4380
rect 55112 4320 55176 4324
rect 55192 4380 55256 4384
rect 55192 4324 55196 4380
rect 55196 4324 55252 4380
rect 55252 4324 55256 4380
rect 55192 4320 55256 4324
rect 90952 4380 91016 4384
rect 90952 4324 90956 4380
rect 90956 4324 91012 4380
rect 91012 4324 91016 4380
rect 90952 4320 91016 4324
rect 91032 4380 91096 4384
rect 91032 4324 91036 4380
rect 91036 4324 91092 4380
rect 91092 4324 91096 4380
rect 91032 4320 91096 4324
rect 91112 4380 91176 4384
rect 91112 4324 91116 4380
rect 91116 4324 91172 4380
rect 91172 4324 91176 4380
rect 91112 4320 91176 4324
rect 91192 4380 91256 4384
rect 91192 4324 91196 4380
rect 91196 4324 91252 4380
rect 91252 4324 91256 4380
rect 91192 4320 91256 4324
rect 36952 3836 37016 3840
rect 36952 3780 36956 3836
rect 36956 3780 37012 3836
rect 37012 3780 37016 3836
rect 36952 3776 37016 3780
rect 37032 3836 37096 3840
rect 37032 3780 37036 3836
rect 37036 3780 37092 3836
rect 37092 3780 37096 3836
rect 37032 3776 37096 3780
rect 37112 3836 37176 3840
rect 37112 3780 37116 3836
rect 37116 3780 37172 3836
rect 37172 3780 37176 3836
rect 37112 3776 37176 3780
rect 37192 3836 37256 3840
rect 37192 3780 37196 3836
rect 37196 3780 37252 3836
rect 37252 3780 37256 3836
rect 37192 3776 37256 3780
rect 72952 3836 73016 3840
rect 72952 3780 72956 3836
rect 72956 3780 73012 3836
rect 73012 3780 73016 3836
rect 72952 3776 73016 3780
rect 73032 3836 73096 3840
rect 73032 3780 73036 3836
rect 73036 3780 73092 3836
rect 73092 3780 73096 3836
rect 73032 3776 73096 3780
rect 73112 3836 73176 3840
rect 73112 3780 73116 3836
rect 73116 3780 73172 3836
rect 73172 3780 73176 3836
rect 73112 3776 73176 3780
rect 73192 3836 73256 3840
rect 73192 3780 73196 3836
rect 73196 3780 73252 3836
rect 73252 3780 73256 3836
rect 73192 3776 73256 3780
rect 18952 3292 19016 3296
rect 18952 3236 18956 3292
rect 18956 3236 19012 3292
rect 19012 3236 19016 3292
rect 18952 3232 19016 3236
rect 19032 3292 19096 3296
rect 19032 3236 19036 3292
rect 19036 3236 19092 3292
rect 19092 3236 19096 3292
rect 19032 3232 19096 3236
rect 19112 3292 19176 3296
rect 19112 3236 19116 3292
rect 19116 3236 19172 3292
rect 19172 3236 19176 3292
rect 19112 3232 19176 3236
rect 19192 3292 19256 3296
rect 19192 3236 19196 3292
rect 19196 3236 19252 3292
rect 19252 3236 19256 3292
rect 19192 3232 19256 3236
rect 54952 3292 55016 3296
rect 54952 3236 54956 3292
rect 54956 3236 55012 3292
rect 55012 3236 55016 3292
rect 54952 3232 55016 3236
rect 55032 3292 55096 3296
rect 55032 3236 55036 3292
rect 55036 3236 55092 3292
rect 55092 3236 55096 3292
rect 55032 3232 55096 3236
rect 55112 3292 55176 3296
rect 55112 3236 55116 3292
rect 55116 3236 55172 3292
rect 55172 3236 55176 3292
rect 55112 3232 55176 3236
rect 55192 3292 55256 3296
rect 55192 3236 55196 3292
rect 55196 3236 55252 3292
rect 55252 3236 55256 3292
rect 55192 3232 55256 3236
rect 90952 3292 91016 3296
rect 90952 3236 90956 3292
rect 90956 3236 91012 3292
rect 91012 3236 91016 3292
rect 90952 3232 91016 3236
rect 91032 3292 91096 3296
rect 91032 3236 91036 3292
rect 91036 3236 91092 3292
rect 91092 3236 91096 3292
rect 91032 3232 91096 3236
rect 91112 3292 91176 3296
rect 91112 3236 91116 3292
rect 91116 3236 91172 3292
rect 91172 3236 91176 3292
rect 91112 3232 91176 3236
rect 91192 3292 91256 3296
rect 91192 3236 91196 3292
rect 91196 3236 91252 3292
rect 91252 3236 91256 3292
rect 91192 3232 91256 3236
rect 36952 2748 37016 2752
rect 36952 2692 36956 2748
rect 36956 2692 37012 2748
rect 37012 2692 37016 2748
rect 36952 2688 37016 2692
rect 37032 2748 37096 2752
rect 37032 2692 37036 2748
rect 37036 2692 37092 2748
rect 37092 2692 37096 2748
rect 37032 2688 37096 2692
rect 37112 2748 37176 2752
rect 37112 2692 37116 2748
rect 37116 2692 37172 2748
rect 37172 2692 37176 2748
rect 37112 2688 37176 2692
rect 37192 2748 37256 2752
rect 37192 2692 37196 2748
rect 37196 2692 37252 2748
rect 37252 2692 37256 2748
rect 37192 2688 37256 2692
rect 72952 2748 73016 2752
rect 72952 2692 72956 2748
rect 72956 2692 73012 2748
rect 73012 2692 73016 2748
rect 72952 2688 73016 2692
rect 73032 2748 73096 2752
rect 73032 2692 73036 2748
rect 73036 2692 73092 2748
rect 73092 2692 73096 2748
rect 73032 2688 73096 2692
rect 73112 2748 73176 2752
rect 73112 2692 73116 2748
rect 73116 2692 73172 2748
rect 73172 2692 73176 2748
rect 73112 2688 73176 2692
rect 73192 2748 73256 2752
rect 73192 2692 73196 2748
rect 73196 2692 73252 2748
rect 73252 2692 73256 2748
rect 73192 2688 73256 2692
rect 18952 2204 19016 2208
rect 18952 2148 18956 2204
rect 18956 2148 19012 2204
rect 19012 2148 19016 2204
rect 18952 2144 19016 2148
rect 19032 2204 19096 2208
rect 19032 2148 19036 2204
rect 19036 2148 19092 2204
rect 19092 2148 19096 2204
rect 19032 2144 19096 2148
rect 19112 2204 19176 2208
rect 19112 2148 19116 2204
rect 19116 2148 19172 2204
rect 19172 2148 19176 2204
rect 19112 2144 19176 2148
rect 19192 2204 19256 2208
rect 19192 2148 19196 2204
rect 19196 2148 19252 2204
rect 19252 2148 19256 2204
rect 19192 2144 19256 2148
rect 54952 2204 55016 2208
rect 54952 2148 54956 2204
rect 54956 2148 55012 2204
rect 55012 2148 55016 2204
rect 54952 2144 55016 2148
rect 55032 2204 55096 2208
rect 55032 2148 55036 2204
rect 55036 2148 55092 2204
rect 55092 2148 55096 2204
rect 55032 2144 55096 2148
rect 55112 2204 55176 2208
rect 55112 2148 55116 2204
rect 55116 2148 55172 2204
rect 55172 2148 55176 2204
rect 55112 2144 55176 2148
rect 55192 2204 55256 2208
rect 55192 2148 55196 2204
rect 55196 2148 55252 2204
rect 55252 2148 55256 2204
rect 55192 2144 55256 2148
rect 90952 2204 91016 2208
rect 90952 2148 90956 2204
rect 90956 2148 91012 2204
rect 91012 2148 91016 2204
rect 90952 2144 91016 2148
rect 91032 2204 91096 2208
rect 91032 2148 91036 2204
rect 91036 2148 91092 2204
rect 91092 2148 91096 2204
rect 91032 2144 91096 2148
rect 91112 2204 91176 2208
rect 91112 2148 91116 2204
rect 91116 2148 91172 2204
rect 91172 2148 91176 2204
rect 91112 2144 91176 2148
rect 91192 2204 91256 2208
rect 91192 2148 91196 2204
rect 91196 2148 91252 2204
rect 91252 2148 91256 2204
rect 91192 2144 91256 2148
<< metal4 >>
rect 18944 10912 19264 11472
rect 18944 10848 18952 10912
rect 19016 10848 19032 10912
rect 19096 10848 19112 10912
rect 19176 10848 19192 10912
rect 19256 10848 19264 10912
rect 18944 9824 19264 10848
rect 18944 9760 18952 9824
rect 19016 9760 19032 9824
rect 19096 9760 19112 9824
rect 19176 9760 19192 9824
rect 19256 9760 19264 9824
rect 18944 8736 19264 9760
rect 18944 8672 18952 8736
rect 19016 8672 19032 8736
rect 19096 8672 19112 8736
rect 19176 8672 19192 8736
rect 19256 8672 19264 8736
rect 18944 7648 19264 8672
rect 18944 7584 18952 7648
rect 19016 7584 19032 7648
rect 19096 7584 19112 7648
rect 19176 7584 19192 7648
rect 19256 7584 19264 7648
rect 18944 6560 19264 7584
rect 18944 6496 18952 6560
rect 19016 6496 19032 6560
rect 19096 6496 19112 6560
rect 19176 6496 19192 6560
rect 19256 6496 19264 6560
rect 18944 5472 19264 6496
rect 18944 5408 18952 5472
rect 19016 5408 19032 5472
rect 19096 5408 19112 5472
rect 19176 5408 19192 5472
rect 19256 5408 19264 5472
rect 18944 4384 19264 5408
rect 18944 4320 18952 4384
rect 19016 4320 19032 4384
rect 19096 4320 19112 4384
rect 19176 4320 19192 4384
rect 19256 4320 19264 4384
rect 18944 3296 19264 4320
rect 18944 3232 18952 3296
rect 19016 3232 19032 3296
rect 19096 3232 19112 3296
rect 19176 3232 19192 3296
rect 19256 3232 19264 3296
rect 18944 2208 19264 3232
rect 18944 2144 18952 2208
rect 19016 2144 19032 2208
rect 19096 2144 19112 2208
rect 19176 2144 19192 2208
rect 19256 2144 19264 2208
rect 18944 2128 19264 2144
rect 36944 11456 37264 11472
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 10368 37264 11392
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 9280 37264 10304
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 8192 37264 9216
rect 36944 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37264 8192
rect 36944 7104 37264 8128
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 6016 37264 7040
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 4928 37264 5952
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 3840 37264 4864
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 2752 37264 3776
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2128 37264 2688
rect 54944 10912 55264 11472
rect 54944 10848 54952 10912
rect 55016 10848 55032 10912
rect 55096 10848 55112 10912
rect 55176 10848 55192 10912
rect 55256 10848 55264 10912
rect 54944 9824 55264 10848
rect 54944 9760 54952 9824
rect 55016 9760 55032 9824
rect 55096 9760 55112 9824
rect 55176 9760 55192 9824
rect 55256 9760 55264 9824
rect 54944 8736 55264 9760
rect 54944 8672 54952 8736
rect 55016 8672 55032 8736
rect 55096 8672 55112 8736
rect 55176 8672 55192 8736
rect 55256 8672 55264 8736
rect 54944 7648 55264 8672
rect 54944 7584 54952 7648
rect 55016 7584 55032 7648
rect 55096 7584 55112 7648
rect 55176 7584 55192 7648
rect 55256 7584 55264 7648
rect 54944 6560 55264 7584
rect 54944 6496 54952 6560
rect 55016 6496 55032 6560
rect 55096 6496 55112 6560
rect 55176 6496 55192 6560
rect 55256 6496 55264 6560
rect 54944 5472 55264 6496
rect 54944 5408 54952 5472
rect 55016 5408 55032 5472
rect 55096 5408 55112 5472
rect 55176 5408 55192 5472
rect 55256 5408 55264 5472
rect 54944 4384 55264 5408
rect 54944 4320 54952 4384
rect 55016 4320 55032 4384
rect 55096 4320 55112 4384
rect 55176 4320 55192 4384
rect 55256 4320 55264 4384
rect 54944 3296 55264 4320
rect 54944 3232 54952 3296
rect 55016 3232 55032 3296
rect 55096 3232 55112 3296
rect 55176 3232 55192 3296
rect 55256 3232 55264 3296
rect 54944 2208 55264 3232
rect 54944 2144 54952 2208
rect 55016 2144 55032 2208
rect 55096 2144 55112 2208
rect 55176 2144 55192 2208
rect 55256 2144 55264 2208
rect 54944 2128 55264 2144
rect 72944 11456 73264 11472
rect 72944 11392 72952 11456
rect 73016 11392 73032 11456
rect 73096 11392 73112 11456
rect 73176 11392 73192 11456
rect 73256 11392 73264 11456
rect 72944 10368 73264 11392
rect 72944 10304 72952 10368
rect 73016 10304 73032 10368
rect 73096 10304 73112 10368
rect 73176 10304 73192 10368
rect 73256 10304 73264 10368
rect 72944 9280 73264 10304
rect 72944 9216 72952 9280
rect 73016 9216 73032 9280
rect 73096 9216 73112 9280
rect 73176 9216 73192 9280
rect 73256 9216 73264 9280
rect 72944 8192 73264 9216
rect 72944 8128 72952 8192
rect 73016 8128 73032 8192
rect 73096 8128 73112 8192
rect 73176 8128 73192 8192
rect 73256 8128 73264 8192
rect 72944 7104 73264 8128
rect 72944 7040 72952 7104
rect 73016 7040 73032 7104
rect 73096 7040 73112 7104
rect 73176 7040 73192 7104
rect 73256 7040 73264 7104
rect 72944 6016 73264 7040
rect 72944 5952 72952 6016
rect 73016 5952 73032 6016
rect 73096 5952 73112 6016
rect 73176 5952 73192 6016
rect 73256 5952 73264 6016
rect 72944 4928 73264 5952
rect 72944 4864 72952 4928
rect 73016 4864 73032 4928
rect 73096 4864 73112 4928
rect 73176 4864 73192 4928
rect 73256 4864 73264 4928
rect 72944 3840 73264 4864
rect 72944 3776 72952 3840
rect 73016 3776 73032 3840
rect 73096 3776 73112 3840
rect 73176 3776 73192 3840
rect 73256 3776 73264 3840
rect 72944 2752 73264 3776
rect 72944 2688 72952 2752
rect 73016 2688 73032 2752
rect 73096 2688 73112 2752
rect 73176 2688 73192 2752
rect 73256 2688 73264 2752
rect 72944 2128 73264 2688
rect 90944 10912 91264 11472
rect 90944 10848 90952 10912
rect 91016 10848 91032 10912
rect 91096 10848 91112 10912
rect 91176 10848 91192 10912
rect 91256 10848 91264 10912
rect 90944 9824 91264 10848
rect 90944 9760 90952 9824
rect 91016 9760 91032 9824
rect 91096 9760 91112 9824
rect 91176 9760 91192 9824
rect 91256 9760 91264 9824
rect 90944 8736 91264 9760
rect 90944 8672 90952 8736
rect 91016 8672 91032 8736
rect 91096 8672 91112 8736
rect 91176 8672 91192 8736
rect 91256 8672 91264 8736
rect 90944 7648 91264 8672
rect 90944 7584 90952 7648
rect 91016 7584 91032 7648
rect 91096 7584 91112 7648
rect 91176 7584 91192 7648
rect 91256 7584 91264 7648
rect 90944 6560 91264 7584
rect 90944 6496 90952 6560
rect 91016 6496 91032 6560
rect 91096 6496 91112 6560
rect 91176 6496 91192 6560
rect 91256 6496 91264 6560
rect 90944 5472 91264 6496
rect 90944 5408 90952 5472
rect 91016 5408 91032 5472
rect 91096 5408 91112 5472
rect 91176 5408 91192 5472
rect 91256 5408 91264 5472
rect 90944 4384 91264 5408
rect 90944 4320 90952 4384
rect 91016 4320 91032 4384
rect 91096 4320 91112 4384
rect 91176 4320 91192 4384
rect 91256 4320 91264 4384
rect 90944 3296 91264 4320
rect 90944 3232 90952 3296
rect 91016 3232 91032 3296
rect 91096 3232 91112 3296
rect 91176 3232 91192 3296
rect 91256 3232 91264 3296
rect 90944 2208 91264 3232
rect 90944 2144 90952 2208
rect 91016 2144 91032 2208
rect 91096 2144 91112 2208
rect 91176 2144 91192 2208
rect 91256 2144 91264 2208
rect 90944 2128 91264 2144
use scs8hd_buf_2  _19_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__19__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_11
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_34 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_35
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_36
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_37
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_38
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_155
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_39
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_40
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_41
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_257 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_42
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_273
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_285
timestamp 1586364061
transform 1 0 27324 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 36064 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 36432 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_379 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_382
timestamp 1586364061
transform 1 0 36248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_386
timestamp 1586364061
transform 1 0 36616 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_398
timestamp 1586364061
transform 1 0 37720 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_410
timestamp 1586364061
transform 1 0 38824 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 39284 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 39836 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_412
timestamp 1586364061
transform 1 0 39008 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_419
timestamp 1586364061
transform 1 0 39652 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_423
timestamp 1586364061
transform 1 0 40020 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_422
timestamp 1586364061
transform 1 0 39928 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_426
timestamp 1586364061
transform 1 0 40296 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_428
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_431
timestamp 1586364061
transform 1 0 40756 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_435
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_440
timestamp 1586364061
transform 1 0 41584 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_447
timestamp 1586364061
transform 1 0 42228 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_459
timestamp 1586364061
transform 1 0 43332 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_452
timestamp 1586364061
transform 1 0 42688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_466
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_478
timestamp 1586364061
transform 1 0 45080 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_464
timestamp 1586364061
transform 1 0 43792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_476
timestamp 1586364061
transform 1 0 44896 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_490
timestamp 1586364061
transform 1 0 46184 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 49588 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_521
timestamp 1586364061
transform 1 0 49036 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_528
timestamp 1586364061
transform 1 0 49680 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_525
timestamp 1586364061
transform 1 0 49404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_540
timestamp 1586364061
transform 1 0 50784 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_552
timestamp 1586364061
transform 1 0 51888 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_537
timestamp 1586364061
transform 1 0 50508 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_550
timestamp 1586364061
transform 1 0 51704 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 53268 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 52440 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 52348 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 52716 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_559
timestamp 1586364061
transform 1 0 52532 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_556
timestamp 1586364061
transform 1 0 52256 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_559
timestamp 1586364061
transform 1 0 52532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_563
timestamp 1586364061
transform 1 0 52900 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 53820 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_571
timestamp 1586364061
transform 1 0 53636 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_575
timestamp 1586364061
transform 1 0 54004 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_587
timestamp 1586364061
transform 1 0 55108 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_575
timestamp 1586364061
transform 1 0 54004 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_587
timestamp 1586364061
transform 1 0 55108 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 55292 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_590
timestamp 1586364061
transform 1 0 55384 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_602
timestamp 1586364061
transform 1 0 56488 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_599
timestamp 1586364061
transform 1 0 56212 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 58144 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 57224 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_614
timestamp 1586364061
transform 1 0 57592 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_621
timestamp 1586364061
transform 1 0 58236 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_607
timestamp 1586364061
transform 1 0 56948 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_611
timestamp 1586364061
transform 1 0 57316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_623
timestamp 1586364061
transform 1 0 58420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_633
timestamp 1586364061
transform 1 0 59340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_635
timestamp 1586364061
transform 1 0 59524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 60996 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_645
timestamp 1586364061
transform 1 0 60444 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_652
timestamp 1586364061
transform 1 0 61088 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_647
timestamp 1586364061
transform 1 0 60628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_659
timestamp 1586364061
transform 1 0 61732 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 62836 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_664
timestamp 1586364061
transform 1 0 62192 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_676
timestamp 1586364061
transform 1 0 63296 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_672
timestamp 1586364061
transform 1 0 62928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 63848 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 64216 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 64584 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_683
timestamp 1586364061
transform 1 0 63940 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_695
timestamp 1586364061
transform 1 0 65044 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_684
timestamp 1586364061
transform 1 0 64032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_688
timestamp 1586364061
transform 1 0 64400 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_692
timestamp 1586364061
transform 1 0 64768 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 66700 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_707
timestamp 1586364061
transform 1 0 66148 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_704
timestamp 1586364061
transform 1 0 65872 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 66792 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 67344 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_718
timestamp 1586364061
transform 1 0 67160 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_722
timestamp 1586364061
transform 1 0 67528 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_716
timestamp 1586364061
transform 1 0 66976 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_728
timestamp 1586364061
transform 1 0 68080 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 69552 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 68448 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_734
timestamp 1586364061
transform 1 0 68632 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_742
timestamp 1586364061
transform 1 0 69368 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_745
timestamp 1586364061
transform 1 0 69644 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_733
timestamp 1586364061
transform 1 0 68540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_745
timestamp 1586364061
transform 1 0 69644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_757
timestamp 1586364061
transform 1 0 70748 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_757
timestamp 1586364061
transform 1 0 70748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 72404 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_769
timestamp 1586364061
transform 1 0 71852 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_776
timestamp 1586364061
transform 1 0 72496 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_769
timestamp 1586364061
transform 1 0 71852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_781
timestamp 1586364061
transform 1 0 72956 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 74060 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_788
timestamp 1586364061
transform 1 0 73600 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_800
timestamp 1586364061
transform 1 0 74704 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_794
timestamp 1586364061
transform 1 0 74152 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 75256 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_807
timestamp 1586364061
transform 1 0 75348 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_819
timestamp 1586364061
transform 1 0 76452 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_806
timestamp 1586364061
transform 1 0 75256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_818
timestamp 1586364061
transform 1 0 76360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 78108 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 78016 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_831
timestamp 1586364061
transform 1 0 77556 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_838
timestamp 1586364061
transform 1 0 78200 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_830
timestamp 1586364061
transform 1 0 77464 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_838
timestamp 1586364061
transform 1 0 78200 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 79672 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 78384 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_850
timestamp 1586364061
transform 1 0 79304 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_842
timestamp 1586364061
transform 1 0 78568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_855
timestamp 1586364061
transform 1 0 79764 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 80040 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 80960 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 80592 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_862
timestamp 1586364061
transform 1 0 80408 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_869
timestamp 1586364061
transform 1 0 81052 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_862
timestamp 1586364061
transform 1 0 80408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_866
timestamp 1586364061
transform 1 0 80776 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_881
timestamp 1586364061
transform 1 0 82156 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_878
timestamp 1586364061
transform 1 0 81880 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_890
timestamp 1586364061
transform 1 0 82984 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 83812 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_893
timestamp 1586364061
transform 1 0 83260 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_900
timestamp 1586364061
transform 1 0 83904 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_902
timestamp 1586364061
transform 1 0 84088 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 85284 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_912
timestamp 1586364061
transform 1 0 85008 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_924
timestamp 1586364061
transform 1 0 86112 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_914
timestamp 1586364061
transform 1 0 85192 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_916
timestamp 1586364061
transform 1 0 85376 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 88044 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 86664 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 87860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_931
timestamp 1586364061
transform 1 0 86756 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_943
timestamp 1586364061
transform 1 0 87860 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_928
timestamp 1586364061
transform 1 0 86480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_940
timestamp 1586364061
transform 1 0 87584 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 89516 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 88596 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 88964 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_955
timestamp 1586364061
transform 1 0 88964 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_962
timestamp 1586364061
transform 1 0 89608 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_949
timestamp 1586364061
transform 1 0 88412 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_953
timestamp 1586364061
transform 1 0 88780 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_957
timestamp 1586364061
transform 1 0 89148 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 90896 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_974
timestamp 1586364061
transform 1 0 90712 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_969
timestamp 1586364061
transform 1 0 90252 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_975
timestamp 1586364061
transform 1 0 90804 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_977
timestamp 1586364061
transform 1 0 90988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 92368 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_986
timestamp 1586364061
transform 1 0 91816 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_993
timestamp 1586364061
transform 1 0 92460 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_989
timestamp 1586364061
transform 1 0 92092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1005
timestamp 1586364061
transform 1 0 93564 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1001
timestamp 1586364061
transform 1 0 93196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1013
timestamp 1586364061
transform 1 0 94300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 95220 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1017
timestamp 1586364061
transform 1 0 94668 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1024
timestamp 1586364061
transform 1 0 95312 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1025
timestamp 1586364061
transform 1 0 95404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 96508 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1036
timestamp 1586364061
transform 1 0 96416 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1048
timestamp 1586364061
transform 1 0 97520 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1038
timestamp 1586364061
transform 1 0 96600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1050
timestamp 1586364061
transform 1 0 97704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 98072 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1055
timestamp 1586364061
transform 1 0 98164 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1067
timestamp 1586364061
transform 1 0 99268 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1062
timestamp 1586364061
transform 1 0 98808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 100924 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1079
timestamp 1586364061
transform 1 0 100372 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1086
timestamp 1586364061
transform 1 0 101016 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1074
timestamp 1586364061
transform 1 0 99912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1086
timestamp 1586364061
transform 1 0 101016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 102120 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1098
timestamp 1586364061
transform 1 0 102120 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1099
timestamp 1586364061
transform 1 0 102212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 103776 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1110
timestamp 1586364061
transform 1 0 103224 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1117
timestamp 1586364061
transform 1 0 103868 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1111
timestamp 1586364061
transform 1 0 103316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1123
timestamp 1586364061
transform 1 0 104420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1129
timestamp 1586364061
transform 1 0 104972 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_1141
timestamp 1586364061
transform 1 0 106076 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_1135
timestamp 1586364061
transform 1 0 105524 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 106812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 106812 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_1145
timestamp 1586364061
transform 1 0 106444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_1143
timestamp 1586364061
transform 1 0 106260 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 36064 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_379
timestamp 1586364061
transform 1 0 35972 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_388
timestamp 1586364061
transform 1 0 36800 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_396
timestamp 1586364061
transform 1 0 37536 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_410
timestamp 1586364061
transform 1 0 38824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_422
timestamp 1586364061
transform 1 0 39928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_434
timestamp 1586364061
transform 1 0 41032 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_446
timestamp 1586364061
transform 1 0 42136 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_459
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_471
timestamp 1586364061
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_483
timestamp 1586364061
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_495
timestamp 1586364061
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_507
timestamp 1586364061
transform 1 0 47748 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_520
timestamp 1586364061
transform 1 0 48944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_532
timestamp 1586364061
transform 1 0 50048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_544
timestamp 1586364061
transform 1 0 51152 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 52348 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_556
timestamp 1586364061
transform 1 0 52256 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_565
timestamp 1586364061
transform 1 0 53084 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_577
timestamp 1586364061
transform 1 0 54188 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_581
timestamp 1586364061
transform 1 0 54556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_593
timestamp 1586364061
transform 1 0 55660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_605
timestamp 1586364061
transform 1 0 56764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_617
timestamp 1586364061
transform 1 0 57868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 60076 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_629
timestamp 1586364061
transform 1 0 58972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_642
timestamp 1586364061
transform 1 0 60168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_654
timestamp 1586364061
transform 1 0 61272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_666
timestamp 1586364061
transform 1 0 62376 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 64216 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_678
timestamp 1586364061
transform 1 0 63480 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_694
timestamp 1586364061
transform 1 0 64952 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 65688 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_703
timestamp 1586364061
transform 1 0 65780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_715
timestamp 1586364061
transform 1 0 66884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_727
timestamp 1586364061
transform 1 0 67988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_739
timestamp 1586364061
transform 1 0 69092 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 71300 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_751
timestamp 1586364061
transform 1 0 70196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_764
timestamp 1586364061
transform 1 0 71392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_776
timestamp 1586364061
transform 1 0 72496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_788
timestamp 1586364061
transform 1 0 73600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_800
timestamp 1586364061
transform 1 0 74704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_812
timestamp 1586364061
transform 1 0 75808 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 78016 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 76912 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_825
timestamp 1586364061
transform 1 0 77004 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_833
timestamp 1586364061
transform 1 0 77740 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_844
timestamp 1586364061
transform 1 0 78752 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_856
timestamp 1586364061
transform 1 0 79856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_868
timestamp 1586364061
transform 1 0 80960 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 82524 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_880
timestamp 1586364061
transform 1 0 82064 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_884
timestamp 1586364061
transform 1 0 82432 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_886
timestamp 1586364061
transform 1 0 82616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_898
timestamp 1586364061
transform 1 0 83720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_910
timestamp 1586364061
transform 1 0 84824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_922
timestamp 1586364061
transform 1 0 85928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_934
timestamp 1586364061
transform 1 0 87032 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 88228 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 88136 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_955
timestamp 1586364061
transform 1 0 88964 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_967
timestamp 1586364061
transform 1 0 90068 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_979
timestamp 1586364061
transform 1 0 91172 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_991
timestamp 1586364061
transform 1 0 92276 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 93748 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_1003
timestamp 1586364061
transform 1 0 93380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_1008
timestamp 1586364061
transform 1 0 93840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1020
timestamp 1586364061
transform 1 0 94944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1032
timestamp 1586364061
transform 1 0 96048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1044
timestamp 1586364061
transform 1 0 97152 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 99360 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1056
timestamp 1586364061
transform 1 0 98256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1069
timestamp 1586364061
transform 1 0 99452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1081
timestamp 1586364061
transform 1 0 100556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1093
timestamp 1586364061
transform 1 0 101660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1105
timestamp 1586364061
transform 1 0 102764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1117
timestamp 1586364061
transform 1 0 103868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 104972 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1130
timestamp 1586364061
transform 1 0 105064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 106812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_1142
timestamp 1586364061
transform 1 0 106168 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_11
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_70
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_82
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 774 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_209
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_221
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35236 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_373
timestamp 1586364061
transform 1 0 35420 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35604 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_377
timestamp 1586364061
transform 1 0 35788 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_389
timestamp 1586364061
transform 1 0 36892 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 37720 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__D
timestamp 1586364061
transform 1 0 38088 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__C
timestamp 1586364061
transform 1 0 38456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__B
timestamp 1586364061
transform 1 0 37352 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_393
timestamp 1586364061
transform 1 0 37260 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_396
timestamp 1586364061
transform 1 0 37536 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_400
timestamp 1586364061
transform 1 0 37904 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_404
timestamp 1586364061
transform 1 0 38272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_408
timestamp 1586364061
transform 1 0 38640 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_420
timestamp 1586364061
transform 1 0 39744 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_426
timestamp 1586364061
transform 1 0 40296 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_428
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_440
timestamp 1586364061
transform 1 0 41584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_452
timestamp 1586364061
transform 1 0 42688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_464
timestamp 1586364061
transform 1 0 43792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_476
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 49864 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_525
timestamp 1586364061
transform 1 0 49404 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_529
timestamp 1586364061
transform 1 0 49772 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_532
timestamp 1586364061
transform 1 0 50048 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_544
timestamp 1586364061
transform 1 0 51152 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_548
timestamp 1586364061
transform 1 0 51520 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_550
timestamp 1586364061
transform 1 0 51704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_562
timestamp 1586364061
transform 1 0 52808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_574
timestamp 1586364061
transform 1 0 53912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_586
timestamp 1586364061
transform 1 0 55016 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 56856 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_598
timestamp 1586364061
transform 1 0 56120 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 57224 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 57500 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_608
timestamp 1586364061
transform 1 0 57040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_611
timestamp 1586364061
transform 1 0 57316 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_615
timestamp 1586364061
transform 1 0 57684 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_627
timestamp 1586364061
transform 1 0 58788 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_639
timestamp 1586364061
transform 1 0 59892 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_651
timestamp 1586364061
transform 1 0 60996 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 62836 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_663
timestamp 1586364061
transform 1 0 62100 0 1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_3_672
timestamp 1586364061
transform 1 0 62928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_684
timestamp 1586364061
transform 1 0 64032 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 65780 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 66148 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_696
timestamp 1586364061
transform 1 0 65136 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_702
timestamp 1586364061
transform 1 0 65688 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_705
timestamp 1586364061
transform 1 0 65964 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_709
timestamp 1586364061
transform 1 0 66332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_721
timestamp 1586364061
transform 1 0 67436 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_729
timestamp 1586364061
transform 1 0 68172 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 68448 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_733
timestamp 1586364061
transform 1 0 68540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_745
timestamp 1586364061
transform 1 0 69644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_757
timestamp 1586364061
transform 1 0 70748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_769
timestamp 1586364061
transform 1 0 71852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_781
timestamp 1586364061
transform 1 0 72956 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 74060 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_794
timestamp 1586364061
transform 1 0 74152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_806
timestamp 1586364061
transform 1 0 75256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_818
timestamp 1586364061
transform 1 0 76360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_830
timestamp 1586364061
transform 1 0 77464 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 79672 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 78844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 79212 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_842
timestamp 1586364061
transform 1 0 78568 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_847
timestamp 1586364061
transform 1 0 79028 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_851
timestamp 1586364061
transform 1 0 79396 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_855
timestamp 1586364061
transform 1 0 79764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_867
timestamp 1586364061
transform 1 0 80868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_879
timestamp 1586364061
transform 1 0 81972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_891
timestamp 1586364061
transform 1 0 83076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_903
timestamp 1586364061
transform 1 0 84180 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 85284 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_916
timestamp 1586364061
transform 1 0 85376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_928
timestamp 1586364061
transform 1 0 86480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_940
timestamp 1586364061
transform 1 0 87584 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 88228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 88596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_946
timestamp 1586364061
transform 1 0 88136 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_949
timestamp 1586364061
transform 1 0 88412 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_953
timestamp 1586364061
transform 1 0 88780 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 90896 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_965
timestamp 1586364061
transform 1 0 89884 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_973
timestamp 1586364061
transform 1 0 90620 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_977
timestamp 1586364061
transform 1 0 90988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_989
timestamp 1586364061
transform 1 0 92092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1001
timestamp 1586364061
transform 1 0 93196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1013
timestamp 1586364061
transform 1 0 94300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1025
timestamp 1586364061
transform 1 0 95404 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 96508 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1038
timestamp 1586364061
transform 1 0 96600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1050
timestamp 1586364061
transform 1 0 97704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1062
timestamp 1586364061
transform 1 0 98808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1074
timestamp 1586364061
transform 1 0 99912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1086
timestamp 1586364061
transform 1 0 101016 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 102120 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1099
timestamp 1586364061
transform 1 0 102212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1111
timestamp 1586364061
transform 1 0 103316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1123
timestamp 1586364061
transform 1 0 104420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_1135
timestamp 1586364061
transform 1 0 105524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 106812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_1143
timestamp 1586364061
transform 1 0 106260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_11
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_14
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_39
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_63
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 35236 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_369
timestamp 1586364061
transform 1 0 35052 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 37076 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_382
timestamp 1586364061
transform 1 0 36248 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_390
timestamp 1586364061
transform 1 0 36984 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _15_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 37444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_393
timestamp 1586364061
transform 1 0 37260 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_415
timestamp 1586364061
transform 1 0 39284 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_427
timestamp 1586364061
transform 1 0 40388 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_439
timestamp 1586364061
transform 1 0 41492 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_451
timestamp 1586364061
transform 1 0 42596 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_457
timestamp 1586364061
transform 1 0 43148 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_483
timestamp 1586364061
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_495
timestamp 1586364061
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_507
timestamp 1586364061
transform 1 0 47748 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _11_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 49864 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_520
timestamp 1586364061
transform 1 0 48944 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_528
timestamp 1586364061
transform 1 0 49680 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_539
timestamp 1586364061
transform 1 0 50692 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_551
timestamp 1586364061
transform 1 0 51796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_563
timestamp 1586364061
transform 1 0 52900 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_575
timestamp 1586364061
transform 1 0 54004 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_579
timestamp 1586364061
transform 1 0 54372 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_581
timestamp 1586364061
transform 1 0 54556 0 -1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 56856 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_4_593
timestamp 1586364061
transform 1 0 55660 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_605
timestamp 1586364061
transform 1 0 56764 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_617
timestamp 1586364061
transform 1 0 57868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 60076 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_629
timestamp 1586364061
transform 1 0 58972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_642
timestamp 1586364061
transform 1 0 60168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_654
timestamp 1586364061
transform 1 0 61272 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 62836 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_666
timestamp 1586364061
transform 1 0 62376 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_670
timestamp 1586364061
transform 1 0 62744 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_673
timestamp 1586364061
transform 1 0 63020 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_685
timestamp 1586364061
transform 1 0 64124 0 -1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 65780 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 65688 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_697
timestamp 1586364061
transform 1 0 65228 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_701
timestamp 1586364061
transform 1 0 65596 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_714
timestamp 1586364061
transform 1 0 66792 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_726
timestamp 1586364061
transform 1 0 67896 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_738
timestamp 1586364061
transform 1 0 69000 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 71300 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_750
timestamp 1586364061
transform 1 0 70104 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_762
timestamp 1586364061
transform 1 0 71208 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_764
timestamp 1586364061
transform 1 0 71392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_776
timestamp 1586364061
transform 1 0 72496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_788
timestamp 1586364061
transform 1 0 73600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_800
timestamp 1586364061
transform 1 0 74704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_812
timestamp 1586364061
transform 1 0 75808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 76912 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 77372 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_825
timestamp 1586364061
transform 1 0 77004 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_831
timestamp 1586364061
transform 1 0 77556 0 -1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 78844 0 -1 4896
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_4_843
timestamp 1586364061
transform 1 0 78660 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_856
timestamp 1586364061
transform 1 0 79856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_868
timestamp 1586364061
transform 1 0 80960 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 82524 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_880
timestamp 1586364061
transform 1 0 82064 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_884
timestamp 1586364061
transform 1 0 82432 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_886
timestamp 1586364061
transform 1 0 82616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_898
timestamp 1586364061
transform 1 0 83720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_910
timestamp 1586364061
transform 1 0 84824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_922
timestamp 1586364061
transform 1 0 85928 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__05__B
timestamp 1586364061
transform 1 0 87768 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_934
timestamp 1586364061
transform 1 0 87032 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_944
timestamp 1586364061
transform 1 0 87952 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 88228 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 88136 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_958
timestamp 1586364061
transform 1 0 89240 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_970
timestamp 1586364061
transform 1 0 90344 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_982
timestamp 1586364061
transform 1 0 91448 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_994
timestamp 1586364061
transform 1 0 92552 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 93748 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_1006
timestamp 1586364061
transform 1 0 93656 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1008
timestamp 1586364061
transform 1 0 93840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1020
timestamp 1586364061
transform 1 0 94944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1032
timestamp 1586364061
transform 1 0 96048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1044
timestamp 1586364061
transform 1 0 97152 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 99360 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1056
timestamp 1586364061
transform 1 0 98256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1069
timestamp 1586364061
transform 1 0 99452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1081
timestamp 1586364061
transform 1 0 100556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1093
timestamp 1586364061
transform 1 0 101660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1105
timestamp 1586364061
transform 1 0 102764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1117
timestamp 1586364061
transform 1 0 103868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 104972 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1130
timestamp 1586364061
transform 1 0 105064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 106812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_1142
timestamp 1586364061
transform 1 0 106168 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_9
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_5_48
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_207
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_219
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 36984 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 36616 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_385
timestamp 1586364061
transform 1 0 36524 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_388
timestamp 1586364061
transform 1 0 36800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_392
timestamp 1586364061
transform 1 0 37168 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 37904 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 37720 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 37352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_396
timestamp 1586364061
transform 1 0 37536 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 39652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_417
timestamp 1586364061
transform 1 0 39468 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_421
timestamp 1586364061
transform 1 0 39836 0 1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_5_428
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_440
timestamp 1586364061
transform 1 0 41584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_452
timestamp 1586364061
transform 1 0 42688 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_464
timestamp 1586364061
transform 1 0 43792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_476
timestamp 1586364061
transform 1 0 44896 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_525
timestamp 1586364061
transform 1 0 49404 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 51060 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_537
timestamp 1586364061
transform 1 0 50508 0 1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_5_545
timestamp 1586364061
transform 1 0 51244 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_550
timestamp 1586364061
transform 1 0 51704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_562
timestamp 1586364061
transform 1 0 52808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_574
timestamp 1586364061
transform 1 0 53912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_586
timestamp 1586364061
transform 1 0 55016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_598
timestamp 1586364061
transform 1 0 56120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 57224 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_611
timestamp 1586364061
transform 1 0 57316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_623
timestamp 1586364061
transform 1 0 58420 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 60168 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 59800 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_635
timestamp 1586364061
transform 1 0 59524 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_640
timestamp 1586364061
transform 1 0 59984 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 60536 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 60904 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_644
timestamp 1586364061
transform 1 0 60352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_648
timestamp 1586364061
transform 1 0 60720 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_652
timestamp 1586364061
transform 1 0 61088 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 62836 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 63112 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 62652 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_664
timestamp 1586364061
transform 1 0 62192 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_668
timestamp 1586364061
transform 1 0 62560 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_672
timestamp 1586364061
transform 1 0 62928 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_676
timestamp 1586364061
transform 1 0 63296 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 63480 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_680
timestamp 1586364061
transform 1 0 63664 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_692
timestamp 1586364061
transform 1 0 64768 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_704
timestamp 1586364061
transform 1 0 65872 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_716
timestamp 1586364061
transform 1 0 66976 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_728
timestamp 1586364061
transform 1 0 68080 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 68448 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 68724 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_733
timestamp 1586364061
transform 1 0 68540 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_737
timestamp 1586364061
transform 1 0 68908 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_749
timestamp 1586364061
transform 1 0 70012 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_761
timestamp 1586364061
transform 1 0 71116 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_773
timestamp 1586364061
transform 1 0 72220 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 74060 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_785
timestamp 1586364061
transform 1 0 73324 0 1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_5_794
timestamp 1586364061
transform 1 0 74152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_806
timestamp 1586364061
transform 1 0 75256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_818
timestamp 1586364061
transform 1 0 76360 0 1 4896
box -38 -48 406 592
use scs8hd_and4_4  _07_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 77372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 77188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 76820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_822
timestamp 1586364061
transform 1 0 76728 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_825
timestamp 1586364061
transform 1 0 77004 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_838
timestamp 1586364061
transform 1 0 78200 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 79672 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_850
timestamp 1586364061
transform 1 0 79304 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_855
timestamp 1586364061
transform 1 0 79764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_867
timestamp 1586364061
transform 1 0 80868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_879
timestamp 1586364061
transform 1 0 81972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_891
timestamp 1586364061
transform 1 0 83076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_903
timestamp 1586364061
transform 1 0 84180 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 85284 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_916
timestamp 1586364061
transform 1 0 85376 0 1 4896
box -38 -48 1142 592
use scs8hd_and4_4  _05_
timestamp 1586364061
transform 1 0 87768 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__05__C
timestamp 1586364061
transform 1 0 87584 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 87216 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_928
timestamp 1586364061
transform 1 0 86480 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_938
timestamp 1586364061
transform 1 0 87400 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_951
timestamp 1586364061
transform 1 0 88596 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_963
timestamp 1586364061
transform 1 0 89700 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 90896 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_975
timestamp 1586364061
transform 1 0 90804 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_977
timestamp 1586364061
transform 1 0 90988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_989
timestamp 1586364061
transform 1 0 92092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1001
timestamp 1586364061
transform 1 0 93196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1013
timestamp 1586364061
transform 1 0 94300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1025
timestamp 1586364061
transform 1 0 95404 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 96508 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1038
timestamp 1586364061
transform 1 0 96600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1050
timestamp 1586364061
transform 1 0 97704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1062
timestamp 1586364061
transform 1 0 98808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1074
timestamp 1586364061
transform 1 0 99912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1086
timestamp 1586364061
transform 1 0 101016 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 102120 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1099
timestamp 1586364061
transform 1 0 102212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1111
timestamp 1586364061
transform 1 0 103316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1123
timestamp 1586364061
transform 1 0 104420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_1135
timestamp 1586364061
transform 1 0 105524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 106812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_1143
timestamp 1586364061
transform 1 0 106260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_300
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__14__C
timestamp 1586364061
transform 1 0 36984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__B
timestamp 1586364061
transform 1 0 36616 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_6  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_385
timestamp 1586364061
transform 1 0 36524 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_388
timestamp 1586364061
transform 1 0 36800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_392
timestamp 1586364061
transform 1 0 37168 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _13_
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _14_
timestamp 1586364061
transform 1 0 37536 0 1 5984
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__14__D
timestamp 1586364061
transform 1 0 37352 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 37444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_393
timestamp 1586364061
transform 1 0 37260 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_415
timestamp 1586364061
transform 1 0 39284 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_427
timestamp 1586364061
transform 1 0 40388 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_413
timestamp 1586364061
transform 1 0 39100 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_425
timestamp 1586364061
transform 1 0 40204 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_439
timestamp 1586364061
transform 1 0 41492 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_440
timestamp 1586364061
transform 1 0 41584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_451
timestamp 1586364061
transform 1 0 42596 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_457
timestamp 1586364061
transform 1 0 43148 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_459
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_452
timestamp 1586364061
transform 1 0 42688 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_471
timestamp 1586364061
transform 1 0 44436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_464
timestamp 1586364061
transform 1 0 43792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_476
timestamp 1586364061
transform 1 0 44896 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_483
timestamp 1586364061
transform 1 0 45540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_495
timestamp 1586364061
transform 1 0 46644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_489
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_507
timestamp 1586364061
transform 1 0 47748 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_501
timestamp 1586364061
transform 1 0 47196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_513
timestamp 1586364061
transform 1 0 48300 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_520
timestamp 1586364061
transform 1 0 48944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_532
timestamp 1586364061
transform 1 0 50048 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_525
timestamp 1586364061
transform 1 0 49404 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _08_
timestamp 1586364061
transform 1 0 51060 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_540
timestamp 1586364061
transform 1 0 50784 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_552
timestamp 1586364061
transform 1 0 51888 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_537
timestamp 1586364061
transform 1 0 50508 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_550
timestamp 1586364061
transform 1 0 51704 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_564
timestamp 1586364061
transform 1 0 52992 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_562
timestamp 1586364061
transform 1 0 52808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_576
timestamp 1586364061
transform 1 0 54096 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_581
timestamp 1586364061
transform 1 0 54556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_574
timestamp 1586364061
transform 1 0 53912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_586
timestamp 1586364061
transform 1 0 55016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_593
timestamp 1586364061
transform 1 0 55660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_605
timestamp 1586364061
transform 1 0 56764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_598
timestamp 1586364061
transform 1 0 56120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 57224 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_617
timestamp 1586364061
transform 1 0 57868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_611
timestamp 1586364061
transform 1 0 57316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_623
timestamp 1586364061
transform 1 0 58420 0 1 5984
box -38 -48 1142 592
use scs8hd_and4_4  _10_
timestamp 1586364061
transform 1 0 60168 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 60076 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_629
timestamp 1586364061
transform 1 0 58972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_635
timestamp 1586364061
transform 1 0 59524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_651
timestamp 1586364061
transform 1 0 60996 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_647
timestamp 1586364061
transform 1 0 60628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_659
timestamp 1586364061
transform 1 0 61732 0 1 5984
box -38 -48 1142 592
use scs8hd_and4_4  _09_
timestamp 1586364061
transform 1 0 62836 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 62836 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_663
timestamp 1586364061
transform 1 0 62100 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_672
timestamp 1586364061
transform 1 0 62928 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_680
timestamp 1586364061
transform 1 0 63664 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_692
timestamp 1586364061
transform 1 0 64768 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_684
timestamp 1586364061
transform 1 0 64032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 65688 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_700
timestamp 1586364061
transform 1 0 65504 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_703
timestamp 1586364061
transform 1 0 65780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_696
timestamp 1586364061
transform 1 0 65136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_708
timestamp 1586364061
transform 1 0 66240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_715
timestamp 1586364061
transform 1 0 66884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_727
timestamp 1586364061
transform 1 0 67988 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_720
timestamp 1586364061
transform 1 0 67344 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _06_
timestamp 1586364061
transform 1 0 68724 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 68448 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_744
timestamp 1586364061
transform 1 0 69552 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_733
timestamp 1586364061
transform 1 0 68540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_745
timestamp 1586364061
transform 1 0 69644 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 71300 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_756
timestamp 1586364061
transform 1 0 70656 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_762
timestamp 1586364061
transform 1 0 71208 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_764
timestamp 1586364061
transform 1 0 71392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_757
timestamp 1586364061
transform 1 0 70748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_776
timestamp 1586364061
transform 1 0 72496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_769
timestamp 1586364061
transform 1 0 71852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_781
timestamp 1586364061
transform 1 0 72956 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 74060 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_788
timestamp 1586364061
transform 1 0 73600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_800
timestamp 1586364061
transform 1 0 74704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_794
timestamp 1586364061
transform 1 0 74152 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_812
timestamp 1586364061
transform 1 0 75808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_806
timestamp 1586364061
transform 1 0 75256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_818
timestamp 1586364061
transform 1 0 76360 0 1 5984
box -38 -48 774 592
use scs8hd_buf_1  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 77280 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 77740 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 77372 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_825
timestamp 1586364061
transform 1 0 77004 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_831
timestamp 1586364061
transform 1 0 77556 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_826
timestamp 1586364061
transform 1 0 77096 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_831
timestamp 1586364061
transform 1 0 77556 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_835
timestamp 1586364061
transform 1 0 77924 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 79672 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_843
timestamp 1586364061
transform 1 0 78660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_855
timestamp 1586364061
transform 1 0 79764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_847
timestamp 1586364061
transform 1 0 79028 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_853
timestamp 1586364061
transform 1 0 79580 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_855
timestamp 1586364061
transform 1 0 79764 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_867
timestamp 1586364061
transform 1 0 80868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_867
timestamp 1586364061
transform 1 0 80868 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 82524 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_879
timestamp 1586364061
transform 1 0 81972 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_6_886
timestamp 1586364061
transform 1 0 82616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_879
timestamp 1586364061
transform 1 0 81972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_891
timestamp 1586364061
transform 1 0 83076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_898
timestamp 1586364061
transform 1 0 83720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_903
timestamp 1586364061
transform 1 0 84180 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 85284 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_910
timestamp 1586364061
transform 1 0 84824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_922
timestamp 1586364061
transform 1 0 85928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_916
timestamp 1586364061
transform 1 0 85376 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__05__D
timestamp 1586364061
transform 1 0 87768 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_934
timestamp 1586364061
transform 1 0 87032 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_944
timestamp 1586364061
transform 1 0 87952 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_928
timestamp 1586364061
transform 1 0 86480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_940
timestamp 1586364061
transform 1 0 87584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 88136 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_947
timestamp 1586364061
transform 1 0 88228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_959
timestamp 1586364061
transform 1 0 89332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_952
timestamp 1586364061
transform 1 0 88688 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 90896 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_971
timestamp 1586364061
transform 1 0 90436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_964
timestamp 1586364061
transform 1 0 89792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_977
timestamp 1586364061
transform 1 0 90988 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_983
timestamp 1586364061
transform 1 0 91540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_995
timestamp 1586364061
transform 1 0 92644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_989
timestamp 1586364061
transform 1 0 92092 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 93748 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1008
timestamp 1586364061
transform 1 0 93840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1001
timestamp 1586364061
transform 1 0 93196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1013
timestamp 1586364061
transform 1 0 94300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1020
timestamp 1586364061
transform 1 0 94944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1032
timestamp 1586364061
transform 1 0 96048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1025
timestamp 1586364061
transform 1 0 95404 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 96508 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1044
timestamp 1586364061
transform 1 0 97152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1038
timestamp 1586364061
transform 1 0 96600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1050
timestamp 1586364061
transform 1 0 97704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 99360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1056
timestamp 1586364061
transform 1 0 98256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1069
timestamp 1586364061
transform 1 0 99452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1062
timestamp 1586364061
transform 1 0 98808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1081
timestamp 1586364061
transform 1 0 100556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1074
timestamp 1586364061
transform 1 0 99912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1086
timestamp 1586364061
transform 1 0 101016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 102120 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1093
timestamp 1586364061
transform 1 0 101660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1105
timestamp 1586364061
transform 1 0 102764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1099
timestamp 1586364061
transform 1 0 102212 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1117
timestamp 1586364061
transform 1 0 103868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1111
timestamp 1586364061
transform 1 0 103316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1123
timestamp 1586364061
transform 1 0 104420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 104972 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1130
timestamp 1586364061
transform 1 0 105064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_1135
timestamp 1586364061
transform 1 0 105524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 106812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 106812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_1142
timestamp 1586364061
transform 1 0 106168 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_1143
timestamp 1586364061
transform 1 0 106260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 37904 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_402
timestamp 1586364061
transform 1 0 38088 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_414
timestamp 1586364061
transform 1 0 39192 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_426
timestamp 1586364061
transform 1 0 40296 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_438
timestamp 1586364061
transform 1 0 41400 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_450
timestamp 1586364061
transform 1 0 42504 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_459
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_471
timestamp 1586364061
transform 1 0 44436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_483
timestamp 1586364061
transform 1 0 45540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_495
timestamp 1586364061
transform 1 0 46644 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_507
timestamp 1586364061
transform 1 0 47748 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_520
timestamp 1586364061
transform 1 0 48944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_532
timestamp 1586364061
transform 1 0 50048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_544
timestamp 1586364061
transform 1 0 51152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_556
timestamp 1586364061
transform 1 0 52256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_568
timestamp 1586364061
transform 1 0 53360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_581
timestamp 1586364061
transform 1 0 54556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_593
timestamp 1586364061
transform 1 0 55660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_605
timestamp 1586364061
transform 1 0 56764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_617
timestamp 1586364061
transform 1 0 57868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 60076 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_629
timestamp 1586364061
transform 1 0 58972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_642
timestamp 1586364061
transform 1 0 60168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_654
timestamp 1586364061
transform 1 0 61272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_666
timestamp 1586364061
transform 1 0 62376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_678
timestamp 1586364061
transform 1 0 63480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_690
timestamp 1586364061
transform 1 0 64584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 65688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_703
timestamp 1586364061
transform 1 0 65780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_715
timestamp 1586364061
transform 1 0 66884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_727
timestamp 1586364061
transform 1 0 67988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_739
timestamp 1586364061
transform 1 0 69092 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 71300 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_751
timestamp 1586364061
transform 1 0 70196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_764
timestamp 1586364061
transform 1 0 71392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_776
timestamp 1586364061
transform 1 0 72496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_788
timestamp 1586364061
transform 1 0 73600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_800
timestamp 1586364061
transform 1 0 74704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_812
timestamp 1586364061
transform 1 0 75808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_825
timestamp 1586364061
transform 1 0 77004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_837
timestamp 1586364061
transform 1 0 78108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_849
timestamp 1586364061
transform 1 0 79212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_861
timestamp 1586364061
transform 1 0 80316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_873
timestamp 1586364061
transform 1 0 81420 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 82524 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_886
timestamp 1586364061
transform 1 0 82616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_898
timestamp 1586364061
transform 1 0 83720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_910
timestamp 1586364061
transform 1 0 84824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_922
timestamp 1586364061
transform 1 0 85928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_934
timestamp 1586364061
transform 1 0 87032 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 88136 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_947
timestamp 1586364061
transform 1 0 88228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_959
timestamp 1586364061
transform 1 0 89332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_971
timestamp 1586364061
transform 1 0 90436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_983
timestamp 1586364061
transform 1 0 91540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_995
timestamp 1586364061
transform 1 0 92644 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 93748 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1008
timestamp 1586364061
transform 1 0 93840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1020
timestamp 1586364061
transform 1 0 94944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1032
timestamp 1586364061
transform 1 0 96048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1044
timestamp 1586364061
transform 1 0 97152 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 99360 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1056
timestamp 1586364061
transform 1 0 98256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1069
timestamp 1586364061
transform 1 0 99452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1081
timestamp 1586364061
transform 1 0 100556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1093
timestamp 1586364061
transform 1 0 101660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1105
timestamp 1586364061
transform 1 0 102764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1117
timestamp 1586364061
transform 1 0 103868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 104972 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1130
timestamp 1586364061
transform 1 0 105064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 106812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_1142
timestamp 1586364061
transform 1 0 106168 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_415
timestamp 1586364061
transform 1 0 39284 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_428
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_440
timestamp 1586364061
transform 1 0 41584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_452
timestamp 1586364061
transform 1 0 42688 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_464
timestamp 1586364061
transform 1 0 43792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_476
timestamp 1586364061
transform 1 0 44896 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_489
timestamp 1586364061
transform 1 0 46092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_501
timestamp 1586364061
transform 1 0 47196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_513
timestamp 1586364061
transform 1 0 48300 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_525
timestamp 1586364061
transform 1 0 49404 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 51612 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_537
timestamp 1586364061
transform 1 0 50508 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_550
timestamp 1586364061
transform 1 0 51704 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_562
timestamp 1586364061
transform 1 0 52808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_574
timestamp 1586364061
transform 1 0 53912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_586
timestamp 1586364061
transform 1 0 55016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_598
timestamp 1586364061
transform 1 0 56120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 57224 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_611
timestamp 1586364061
transform 1 0 57316 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_623
timestamp 1586364061
transform 1 0 58420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_635
timestamp 1586364061
transform 1 0 59524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_647
timestamp 1586364061
transform 1 0 60628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_659
timestamp 1586364061
transform 1 0 61732 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 62836 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_672
timestamp 1586364061
transform 1 0 62928 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_684
timestamp 1586364061
transform 1 0 64032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_696
timestamp 1586364061
transform 1 0 65136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_708
timestamp 1586364061
transform 1 0 66240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_720
timestamp 1586364061
transform 1 0 67344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 68448 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_733
timestamp 1586364061
transform 1 0 68540 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_745
timestamp 1586364061
transform 1 0 69644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_757
timestamp 1586364061
transform 1 0 70748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_769
timestamp 1586364061
transform 1 0 71852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_781
timestamp 1586364061
transform 1 0 72956 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 74060 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_794
timestamp 1586364061
transform 1 0 74152 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_806
timestamp 1586364061
transform 1 0 75256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_818
timestamp 1586364061
transform 1 0 76360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_830
timestamp 1586364061
transform 1 0 77464 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 79672 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_842
timestamp 1586364061
transform 1 0 78568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_855
timestamp 1586364061
transform 1 0 79764 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_867
timestamp 1586364061
transform 1 0 80868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_879
timestamp 1586364061
transform 1 0 81972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_891
timestamp 1586364061
transform 1 0 83076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_903
timestamp 1586364061
transform 1 0 84180 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 85284 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_916
timestamp 1586364061
transform 1 0 85376 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_928
timestamp 1586364061
transform 1 0 86480 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_940
timestamp 1586364061
transform 1 0 87584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_952
timestamp 1586364061
transform 1 0 88688 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 90896 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_964
timestamp 1586364061
transform 1 0 89792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_977
timestamp 1586364061
transform 1 0 90988 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_989
timestamp 1586364061
transform 1 0 92092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1001
timestamp 1586364061
transform 1 0 93196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1013
timestamp 1586364061
transform 1 0 94300 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1025
timestamp 1586364061
transform 1 0 95404 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 96508 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1038
timestamp 1586364061
transform 1 0 96600 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1050
timestamp 1586364061
transform 1 0 97704 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1062
timestamp 1586364061
transform 1 0 98808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1074
timestamp 1586364061
transform 1 0 99912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1086
timestamp 1586364061
transform 1 0 101016 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 102120 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1099
timestamp 1586364061
transform 1 0 102212 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1111
timestamp 1586364061
transform 1 0 103316 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1123
timestamp 1586364061
transform 1 0 104420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_1135
timestamp 1586364061
transform 1 0 105524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 106812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_1143
timestamp 1586364061
transform 1 0 106260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_373
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_385
timestamp 1586364061
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_410
timestamp 1586364061
transform 1 0 38824 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_422
timestamp 1586364061
transform 1 0 39928 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_434
timestamp 1586364061
transform 1 0 41032 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_446
timestamp 1586364061
transform 1 0 42136 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_459
timestamp 1586364061
transform 1 0 43332 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_471
timestamp 1586364061
transform 1 0 44436 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_483
timestamp 1586364061
transform 1 0 45540 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_495
timestamp 1586364061
transform 1 0 46644 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_507
timestamp 1586364061
transform 1 0 47748 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 48852 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_520
timestamp 1586364061
transform 1 0 48944 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_532
timestamp 1586364061
transform 1 0 50048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_544
timestamp 1586364061
transform 1 0 51152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_556
timestamp 1586364061
transform 1 0 52256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_568
timestamp 1586364061
transform 1 0 53360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 54464 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_581
timestamp 1586364061
transform 1 0 54556 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_593
timestamp 1586364061
transform 1 0 55660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_605
timestamp 1586364061
transform 1 0 56764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_617
timestamp 1586364061
transform 1 0 57868 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 60076 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_629
timestamp 1586364061
transform 1 0 58972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_642
timestamp 1586364061
transform 1 0 60168 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_654
timestamp 1586364061
transform 1 0 61272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_666
timestamp 1586364061
transform 1 0 62376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_678
timestamp 1586364061
transform 1 0 63480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_690
timestamp 1586364061
transform 1 0 64584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 65688 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_703
timestamp 1586364061
transform 1 0 65780 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_715
timestamp 1586364061
transform 1 0 66884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_727
timestamp 1586364061
transform 1 0 67988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_739
timestamp 1586364061
transform 1 0 69092 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 71300 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_751
timestamp 1586364061
transform 1 0 70196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_764
timestamp 1586364061
transform 1 0 71392 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_776
timestamp 1586364061
transform 1 0 72496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_788
timestamp 1586364061
transform 1 0 73600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_800
timestamp 1586364061
transform 1 0 74704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_812
timestamp 1586364061
transform 1 0 75808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 76912 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_825
timestamp 1586364061
transform 1 0 77004 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_837
timestamp 1586364061
transform 1 0 78108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_849
timestamp 1586364061
transform 1 0 79212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_861
timestamp 1586364061
transform 1 0 80316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_873
timestamp 1586364061
transform 1 0 81420 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 82524 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_886
timestamp 1586364061
transform 1 0 82616 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_898
timestamp 1586364061
transform 1 0 83720 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_910
timestamp 1586364061
transform 1 0 84824 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_922
timestamp 1586364061
transform 1 0 85928 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_934
timestamp 1586364061
transform 1 0 87032 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 88136 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_947
timestamp 1586364061
transform 1 0 88228 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_959
timestamp 1586364061
transform 1 0 89332 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_971
timestamp 1586364061
transform 1 0 90436 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_983
timestamp 1586364061
transform 1 0 91540 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_995
timestamp 1586364061
transform 1 0 92644 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 93748 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_1008
timestamp 1586364061
transform 1 0 93840 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1020
timestamp 1586364061
transform 1 0 94944 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1032
timestamp 1586364061
transform 1 0 96048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1044
timestamp 1586364061
transform 1 0 97152 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 99360 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_1056
timestamp 1586364061
transform 1 0 98256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1069
timestamp 1586364061
transform 1 0 99452 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1081
timestamp 1586364061
transform 1 0 100556 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1093
timestamp 1586364061
transform 1 0 101660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1105
timestamp 1586364061
transform 1 0 102764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1117
timestamp 1586364061
transform 1 0 103868 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 104972 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_1130
timestamp 1586364061
transform 1 0 105064 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 106812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_1142
timestamp 1586364061
transform 1 0 106168 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_354
timestamp 1586364061
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_379
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_391
timestamp 1586364061
transform 1 0 37076 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_415
timestamp 1586364061
transform 1 0 39284 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_428
timestamp 1586364061
transform 1 0 40480 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_440
timestamp 1586364061
transform 1 0 41584 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_452
timestamp 1586364061
transform 1 0 42688 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_464
timestamp 1586364061
transform 1 0 43792 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_476
timestamp 1586364061
transform 1 0 44896 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_489
timestamp 1586364061
transform 1 0 46092 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_501
timestamp 1586364061
transform 1 0 47196 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_513
timestamp 1586364061
transform 1 0 48300 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_525
timestamp 1586364061
transform 1 0 49404 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 51612 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_537
timestamp 1586364061
transform 1 0 50508 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_550
timestamp 1586364061
transform 1 0 51704 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_562
timestamp 1586364061
transform 1 0 52808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_574
timestamp 1586364061
transform 1 0 53912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_586
timestamp 1586364061
transform 1 0 55016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_598
timestamp 1586364061
transform 1 0 56120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 57224 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_611
timestamp 1586364061
transform 1 0 57316 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_623
timestamp 1586364061
transform 1 0 58420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_635
timestamp 1586364061
transform 1 0 59524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_647
timestamp 1586364061
transform 1 0 60628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_659
timestamp 1586364061
transform 1 0 61732 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 62836 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_672
timestamp 1586364061
transform 1 0 62928 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_684
timestamp 1586364061
transform 1 0 64032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_696
timestamp 1586364061
transform 1 0 65136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_708
timestamp 1586364061
transform 1 0 66240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_720
timestamp 1586364061
transform 1 0 67344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 68448 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_733
timestamp 1586364061
transform 1 0 68540 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_745
timestamp 1586364061
transform 1 0 69644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_757
timestamp 1586364061
transform 1 0 70748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_769
timestamp 1586364061
transform 1 0 71852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_781
timestamp 1586364061
transform 1 0 72956 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 74060 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_794
timestamp 1586364061
transform 1 0 74152 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_806
timestamp 1586364061
transform 1 0 75256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_818
timestamp 1586364061
transform 1 0 76360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_830
timestamp 1586364061
transform 1 0 77464 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 79672 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_842
timestamp 1586364061
transform 1 0 78568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_855
timestamp 1586364061
transform 1 0 79764 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_867
timestamp 1586364061
transform 1 0 80868 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_879
timestamp 1586364061
transform 1 0 81972 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_891
timestamp 1586364061
transform 1 0 83076 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_903
timestamp 1586364061
transform 1 0 84180 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 85284 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_916
timestamp 1586364061
transform 1 0 85376 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_928
timestamp 1586364061
transform 1 0 86480 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_940
timestamp 1586364061
transform 1 0 87584 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_952
timestamp 1586364061
transform 1 0 88688 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 90896 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_964
timestamp 1586364061
transform 1 0 89792 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_977
timestamp 1586364061
transform 1 0 90988 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_989
timestamp 1586364061
transform 1 0 92092 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1001
timestamp 1586364061
transform 1 0 93196 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1013
timestamp 1586364061
transform 1 0 94300 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1025
timestamp 1586364061
transform 1 0 95404 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 96508 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_1038
timestamp 1586364061
transform 1 0 96600 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1050
timestamp 1586364061
transform 1 0 97704 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1062
timestamp 1586364061
transform 1 0 98808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1074
timestamp 1586364061
transform 1 0 99912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1086
timestamp 1586364061
transform 1 0 101016 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 102120 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_1099
timestamp 1586364061
transform 1 0 102212 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1111
timestamp 1586364061
transform 1 0 103316 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1123
timestamp 1586364061
transform 1 0 104420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_1135
timestamp 1586364061
transform 1 0 105524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 106812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_1143
timestamp 1586364061
transform 1 0 106260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_373
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_385
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_410
timestamp 1586364061
transform 1 0 38824 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_422
timestamp 1586364061
transform 1 0 39928 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_434
timestamp 1586364061
transform 1 0 41032 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_446
timestamp 1586364061
transform 1 0 42136 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_459
timestamp 1586364061
transform 1 0 43332 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_471
timestamp 1586364061
transform 1 0 44436 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_483
timestamp 1586364061
transform 1 0 45540 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_495
timestamp 1586364061
transform 1 0 46644 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_507
timestamp 1586364061
transform 1 0 47748 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 48852 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_520
timestamp 1586364061
transform 1 0 48944 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_532
timestamp 1586364061
transform 1 0 50048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_544
timestamp 1586364061
transform 1 0 51152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_556
timestamp 1586364061
transform 1 0 52256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_568
timestamp 1586364061
transform 1 0 53360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 54464 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_581
timestamp 1586364061
transform 1 0 54556 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_593
timestamp 1586364061
transform 1 0 55660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_605
timestamp 1586364061
transform 1 0 56764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_617
timestamp 1586364061
transform 1 0 57868 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 60076 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_629
timestamp 1586364061
transform 1 0 58972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_642
timestamp 1586364061
transform 1 0 60168 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_654
timestamp 1586364061
transform 1 0 61272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_666
timestamp 1586364061
transform 1 0 62376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_678
timestamp 1586364061
transform 1 0 63480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_690
timestamp 1586364061
transform 1 0 64584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 65688 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_703
timestamp 1586364061
transform 1 0 65780 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_715
timestamp 1586364061
transform 1 0 66884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_727
timestamp 1586364061
transform 1 0 67988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_739
timestamp 1586364061
transform 1 0 69092 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 71300 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_751
timestamp 1586364061
transform 1 0 70196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_764
timestamp 1586364061
transform 1 0 71392 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_776
timestamp 1586364061
transform 1 0 72496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_788
timestamp 1586364061
transform 1 0 73600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_800
timestamp 1586364061
transform 1 0 74704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_812
timestamp 1586364061
transform 1 0 75808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 76912 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_825
timestamp 1586364061
transform 1 0 77004 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_837
timestamp 1586364061
transform 1 0 78108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_849
timestamp 1586364061
transform 1 0 79212 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_861
timestamp 1586364061
transform 1 0 80316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_873
timestamp 1586364061
transform 1 0 81420 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 82524 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_886
timestamp 1586364061
transform 1 0 82616 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_898
timestamp 1586364061
transform 1 0 83720 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_910
timestamp 1586364061
transform 1 0 84824 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_922
timestamp 1586364061
transform 1 0 85928 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_934
timestamp 1586364061
transform 1 0 87032 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 88136 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_947
timestamp 1586364061
transform 1 0 88228 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_959
timestamp 1586364061
transform 1 0 89332 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_971
timestamp 1586364061
transform 1 0 90436 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_983
timestamp 1586364061
transform 1 0 91540 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_995
timestamp 1586364061
transform 1 0 92644 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 93748 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_1008
timestamp 1586364061
transform 1 0 93840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1020
timestamp 1586364061
transform 1 0 94944 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1032
timestamp 1586364061
transform 1 0 96048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1044
timestamp 1586364061
transform 1 0 97152 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 99360 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_1056
timestamp 1586364061
transform 1 0 98256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1069
timestamp 1586364061
transform 1 0 99452 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1081
timestamp 1586364061
transform 1 0 100556 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1093
timestamp 1586364061
transform 1 0 101660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1105
timestamp 1586364061
transform 1 0 102764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1117
timestamp 1586364061
transform 1 0 103868 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 104972 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_1130
timestamp 1586364061
transform 1 0 105064 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 106812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_1142
timestamp 1586364061
transform 1 0 106168 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_373
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_379
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_391
timestamp 1586364061
transform 1 0 37076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_385
timestamp 1586364061
transform 1 0 36524 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_403
timestamp 1586364061
transform 1 0 38180 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_410
timestamp 1586364061
transform 1 0 38824 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_415
timestamp 1586364061
transform 1 0 39284 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_428
timestamp 1586364061
transform 1 0 40480 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_422
timestamp 1586364061
transform 1 0 39928 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_440
timestamp 1586364061
transform 1 0 41584 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_434
timestamp 1586364061
transform 1 0 41032 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_452
timestamp 1586364061
transform 1 0 42688 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_446
timestamp 1586364061
transform 1 0 42136 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_459
timestamp 1586364061
transform 1 0 43332 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_464
timestamp 1586364061
transform 1 0 43792 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_476
timestamp 1586364061
transform 1 0 44896 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_471
timestamp 1586364061
transform 1 0 44436 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_489
timestamp 1586364061
transform 1 0 46092 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_483
timestamp 1586364061
transform 1 0 45540 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_495
timestamp 1586364061
transform 1 0 46644 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_501
timestamp 1586364061
transform 1 0 47196 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_513
timestamp 1586364061
transform 1 0 48300 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_507
timestamp 1586364061
transform 1 0 47748 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 48852 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_525
timestamp 1586364061
transform 1 0 49404 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_520
timestamp 1586364061
transform 1 0 48944 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_532
timestamp 1586364061
transform 1 0 50048 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 51612 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_537
timestamp 1586364061
transform 1 0 50508 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_550
timestamp 1586364061
transform 1 0 51704 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_544
timestamp 1586364061
transform 1 0 51152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_562
timestamp 1586364061
transform 1 0 52808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_556
timestamp 1586364061
transform 1 0 52256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_568
timestamp 1586364061
transform 1 0 53360 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 54464 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_574
timestamp 1586364061
transform 1 0 53912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_586
timestamp 1586364061
transform 1 0 55016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_581
timestamp 1586364061
transform 1 0 54556 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_598
timestamp 1586364061
transform 1 0 56120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_593
timestamp 1586364061
transform 1 0 55660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_605
timestamp 1586364061
transform 1 0 56764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 57224 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_611
timestamp 1586364061
transform 1 0 57316 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_623
timestamp 1586364061
transform 1 0 58420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_617
timestamp 1586364061
transform 1 0 57868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 60076 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_635
timestamp 1586364061
transform 1 0 59524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_629
timestamp 1586364061
transform 1 0 58972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_642
timestamp 1586364061
transform 1 0 60168 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_647
timestamp 1586364061
transform 1 0 60628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_659
timestamp 1586364061
transform 1 0 61732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_654
timestamp 1586364061
transform 1 0 61272 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 62836 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_672
timestamp 1586364061
transform 1 0 62928 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_666
timestamp 1586364061
transform 1 0 62376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_684
timestamp 1586364061
transform 1 0 64032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_678
timestamp 1586364061
transform 1 0 63480 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_690
timestamp 1586364061
transform 1 0 64584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 65688 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_696
timestamp 1586364061
transform 1 0 65136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_708
timestamp 1586364061
transform 1 0 66240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_703
timestamp 1586364061
transform 1 0 65780 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_720
timestamp 1586364061
transform 1 0 67344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_715
timestamp 1586364061
transform 1 0 66884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_727
timestamp 1586364061
transform 1 0 67988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 68448 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_733
timestamp 1586364061
transform 1 0 68540 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_745
timestamp 1586364061
transform 1 0 69644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_739
timestamp 1586364061
transform 1 0 69092 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 71300 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_757
timestamp 1586364061
transform 1 0 70748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_751
timestamp 1586364061
transform 1 0 70196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_764
timestamp 1586364061
transform 1 0 71392 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_769
timestamp 1586364061
transform 1 0 71852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_781
timestamp 1586364061
transform 1 0 72956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_776
timestamp 1586364061
transform 1 0 72496 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 74060 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_794
timestamp 1586364061
transform 1 0 74152 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_788
timestamp 1586364061
transform 1 0 73600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_800
timestamp 1586364061
transform 1 0 74704 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_806
timestamp 1586364061
transform 1 0 75256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_818
timestamp 1586364061
transform 1 0 76360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_812
timestamp 1586364061
transform 1 0 75808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 76912 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_830
timestamp 1586364061
transform 1 0 77464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_825
timestamp 1586364061
transform 1 0 77004 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_837
timestamp 1586364061
transform 1 0 78108 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 79672 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_842
timestamp 1586364061
transform 1 0 78568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_855
timestamp 1586364061
transform 1 0 79764 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_849
timestamp 1586364061
transform 1 0 79212 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_867
timestamp 1586364061
transform 1 0 80868 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_861
timestamp 1586364061
transform 1 0 80316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_873
timestamp 1586364061
transform 1 0 81420 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 82524 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_879
timestamp 1586364061
transform 1 0 81972 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_891
timestamp 1586364061
transform 1 0 83076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_886
timestamp 1586364061
transform 1 0 82616 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_903
timestamp 1586364061
transform 1 0 84180 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_898
timestamp 1586364061
transform 1 0 83720 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 85284 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_916
timestamp 1586364061
transform 1 0 85376 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_910
timestamp 1586364061
transform 1 0 84824 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_922
timestamp 1586364061
transform 1 0 85928 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_928
timestamp 1586364061
transform 1 0 86480 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_940
timestamp 1586364061
transform 1 0 87584 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_934
timestamp 1586364061
transform 1 0 87032 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 88136 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_952
timestamp 1586364061
transform 1 0 88688 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_947
timestamp 1586364061
transform 1 0 88228 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_959
timestamp 1586364061
transform 1 0 89332 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 90896 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_964
timestamp 1586364061
transform 1 0 89792 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_977
timestamp 1586364061
transform 1 0 90988 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_971
timestamp 1586364061
transform 1 0 90436 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_989
timestamp 1586364061
transform 1 0 92092 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_983
timestamp 1586364061
transform 1 0 91540 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_995
timestamp 1586364061
transform 1 0 92644 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 93748 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1001
timestamp 1586364061
transform 1 0 93196 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1013
timestamp 1586364061
transform 1 0 94300 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1008
timestamp 1586364061
transform 1 0 93840 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1025
timestamp 1586364061
transform 1 0 95404 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1020
timestamp 1586364061
transform 1 0 94944 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1032
timestamp 1586364061
transform 1 0 96048 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 96508 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1038
timestamp 1586364061
transform 1 0 96600 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1050
timestamp 1586364061
transform 1 0 97704 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1044
timestamp 1586364061
transform 1 0 97152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 99360 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1062
timestamp 1586364061
transform 1 0 98808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1056
timestamp 1586364061
transform 1 0 98256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1069
timestamp 1586364061
transform 1 0 99452 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1074
timestamp 1586364061
transform 1 0 99912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1086
timestamp 1586364061
transform 1 0 101016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1081
timestamp 1586364061
transform 1 0 100556 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 102120 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1099
timestamp 1586364061
transform 1 0 102212 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1093
timestamp 1586364061
transform 1 0 101660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1105
timestamp 1586364061
transform 1 0 102764 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1111
timestamp 1586364061
transform 1 0 103316 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1123
timestamp 1586364061
transform 1 0 104420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1117
timestamp 1586364061
transform 1 0 103868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 104972 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_1135
timestamp 1586364061
transform 1 0 105524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_1130
timestamp 1586364061
transform 1 0 105064 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 106812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 106812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_1143
timestamp 1586364061
transform 1 0 106260 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_1142
timestamp 1586364061
transform 1 0 106168 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_379
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_415
timestamp 1586364061
transform 1 0 39284 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_428
timestamp 1586364061
transform 1 0 40480 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_440
timestamp 1586364061
transform 1 0 41584 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_452
timestamp 1586364061
transform 1 0 42688 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_464
timestamp 1586364061
transform 1 0 43792 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_476
timestamp 1586364061
transform 1 0 44896 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_489
timestamp 1586364061
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_501
timestamp 1586364061
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_513
timestamp 1586364061
transform 1 0 48300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_525
timestamp 1586364061
transform 1 0 49404 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 51612 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_537
timestamp 1586364061
transform 1 0 50508 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_550
timestamp 1586364061
transform 1 0 51704 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_562
timestamp 1586364061
transform 1 0 52808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_574
timestamp 1586364061
transform 1 0 53912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_586
timestamp 1586364061
transform 1 0 55016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_598
timestamp 1586364061
transform 1 0 56120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 57224 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_611
timestamp 1586364061
transform 1 0 57316 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_623
timestamp 1586364061
transform 1 0 58420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_635
timestamp 1586364061
transform 1 0 59524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_647
timestamp 1586364061
transform 1 0 60628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_659
timestamp 1586364061
transform 1 0 61732 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 62836 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_672
timestamp 1586364061
transform 1 0 62928 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_684
timestamp 1586364061
transform 1 0 64032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_696
timestamp 1586364061
transform 1 0 65136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_708
timestamp 1586364061
transform 1 0 66240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_720
timestamp 1586364061
transform 1 0 67344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 68448 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_733
timestamp 1586364061
transform 1 0 68540 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_745
timestamp 1586364061
transform 1 0 69644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_757
timestamp 1586364061
transform 1 0 70748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_769
timestamp 1586364061
transform 1 0 71852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_781
timestamp 1586364061
transform 1 0 72956 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 74060 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_794
timestamp 1586364061
transform 1 0 74152 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_806
timestamp 1586364061
transform 1 0 75256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_818
timestamp 1586364061
transform 1 0 76360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_830
timestamp 1586364061
transform 1 0 77464 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 79672 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_842
timestamp 1586364061
transform 1 0 78568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_855
timestamp 1586364061
transform 1 0 79764 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_867
timestamp 1586364061
transform 1 0 80868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_879
timestamp 1586364061
transform 1 0 81972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_891
timestamp 1586364061
transform 1 0 83076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_903
timestamp 1586364061
transform 1 0 84180 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 85284 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_916
timestamp 1586364061
transform 1 0 85376 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_928
timestamp 1586364061
transform 1 0 86480 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_940
timestamp 1586364061
transform 1 0 87584 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_952
timestamp 1586364061
transform 1 0 88688 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 90896 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_964
timestamp 1586364061
transform 1 0 89792 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_977
timestamp 1586364061
transform 1 0 90988 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_989
timestamp 1586364061
transform 1 0 92092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1001
timestamp 1586364061
transform 1 0 93196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1013
timestamp 1586364061
transform 1 0 94300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1025
timestamp 1586364061
transform 1 0 95404 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 96508 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_1038
timestamp 1586364061
transform 1 0 96600 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1050
timestamp 1586364061
transform 1 0 97704 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1062
timestamp 1586364061
transform 1 0 98808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1074
timestamp 1586364061
transform 1 0 99912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1086
timestamp 1586364061
transform 1 0 101016 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 102120 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_1099
timestamp 1586364061
transform 1 0 102212 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1111
timestamp 1586364061
transform 1 0 103316 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1123
timestamp 1586364061
transform 1 0 104420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_1135
timestamp 1586364061
transform 1 0 105524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 106812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_1143
timestamp 1586364061
transform 1 0 106260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_75
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_94
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_118
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 15364 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_156
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_242
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_249
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_261
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 26772 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_273
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_280
timestamp 1586364061
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_292
timestamp 1586364061
transform 1 0 27968 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 29624 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_304
timestamp 1586364061
transform 1 0 29072 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_311
timestamp 1586364061
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_323
timestamp 1586364061
transform 1 0 30820 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_335
timestamp 1586364061
transform 1 0 31924 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 32476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_342
timestamp 1586364061
transform 1 0 32568 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_354
timestamp 1586364061
transform 1 0 33672 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 35328 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_366
timestamp 1586364061
transform 1 0 34776 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_385
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 38180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_397
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_404
timestamp 1586364061
transform 1 0 38272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_416
timestamp 1586364061
transform 1 0 39376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_428
timestamp 1586364061
transform 1 0 40480 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 41032 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_435
timestamp 1586364061
transform 1 0 41124 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_447
timestamp 1586364061
transform 1 0 42228 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_459
timestamp 1586364061
transform 1 0 43332 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 43884 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_466
timestamp 1586364061
transform 1 0 43976 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_478
timestamp 1586364061
transform 1 0 45080 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 46736 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_490
timestamp 1586364061
transform 1 0 46184 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_497
timestamp 1586364061
transform 1 0 46828 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_509
timestamp 1586364061
transform 1 0 47932 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 49588 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_521
timestamp 1586364061
transform 1 0 49036 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_528
timestamp 1586364061
transform 1 0 49680 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_540
timestamp 1586364061
transform 1 0 50784 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_552
timestamp 1586364061
transform 1 0 51888 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 52440 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_559
timestamp 1586364061
transform 1 0 52532 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_571
timestamp 1586364061
transform 1 0 53636 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_583
timestamp 1586364061
transform 1 0 54740 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 55292 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_590
timestamp 1586364061
transform 1 0 55384 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_602
timestamp 1586364061
transform 1 0 56488 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 58144 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_614
timestamp 1586364061
transform 1 0 57592 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_621
timestamp 1586364061
transform 1 0 58236 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_633
timestamp 1586364061
transform 1 0 59340 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 60996 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_645
timestamp 1586364061
transform 1 0 60444 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_652
timestamp 1586364061
transform 1 0 61088 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_664
timestamp 1586364061
transform 1 0 62192 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_676
timestamp 1586364061
transform 1 0 63296 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 63848 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_683
timestamp 1586364061
transform 1 0 63940 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_695
timestamp 1586364061
transform 1 0 65044 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 66700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_707
timestamp 1586364061
transform 1 0 66148 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_714
timestamp 1586364061
transform 1 0 66792 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_726
timestamp 1586364061
transform 1 0 67896 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 69552 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_738
timestamp 1586364061
transform 1 0 69000 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_745
timestamp 1586364061
transform 1 0 69644 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_757
timestamp 1586364061
transform 1 0 70748 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 72404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_769
timestamp 1586364061
transform 1 0 71852 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_776
timestamp 1586364061
transform 1 0 72496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_788
timestamp 1586364061
transform 1 0 73600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_800
timestamp 1586364061
transform 1 0 74704 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 75256 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_807
timestamp 1586364061
transform 1 0 75348 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_819
timestamp 1586364061
transform 1 0 76452 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 78108 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_831
timestamp 1586364061
transform 1 0 77556 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_838
timestamp 1586364061
transform 1 0 78200 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_850
timestamp 1586364061
transform 1 0 79304 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 80960 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_862
timestamp 1586364061
transform 1 0 80408 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_869
timestamp 1586364061
transform 1 0 81052 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_881
timestamp 1586364061
transform 1 0 82156 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 83812 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_893
timestamp 1586364061
transform 1 0 83260 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_900
timestamp 1586364061
transform 1 0 83904 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_912
timestamp 1586364061
transform 1 0 85008 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_924
timestamp 1586364061
transform 1 0 86112 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 86664 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_931
timestamp 1586364061
transform 1 0 86756 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_943
timestamp 1586364061
transform 1 0 87860 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 89516 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_955
timestamp 1586364061
transform 1 0 88964 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_962
timestamp 1586364061
transform 1 0 89608 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_974
timestamp 1586364061
transform 1 0 90712 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 92368 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_986
timestamp 1586364061
transform 1 0 91816 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_993
timestamp 1586364061
transform 1 0 92460 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1005
timestamp 1586364061
transform 1 0 93564 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 95220 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_1017
timestamp 1586364061
transform 1 0 94668 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_1024
timestamp 1586364061
transform 1 0 95312 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1036
timestamp 1586364061
transform 1 0 96416 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_1048
timestamp 1586364061
transform 1 0 97520 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 98072 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_1055
timestamp 1586364061
transform 1 0 98164 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1067
timestamp 1586364061
transform 1 0 99268 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 100924 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_1079
timestamp 1586364061
transform 1 0 100372 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_1086
timestamp 1586364061
transform 1 0 101016 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1098
timestamp 1586364061
transform 1 0 102120 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 103776 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_1110
timestamp 1586364061
transform 1 0 103224 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_1117
timestamp 1586364061
transform 1 0 103868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1129
timestamp 1586364061
transform 1 0 104972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_1141
timestamp 1586364061
transform 1 0 106076 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 106812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_1145
timestamp 1586364061
transform 1 0 106444 0 -1 11424
box -38 -48 130 592
<< labels >>
rlabel metal3 s 107520 3408 108000 3528 6 address[0]
port 0 nsew default input
rlabel metal3 s 107520 5720 108000 5840 6 address[1]
port 1 nsew default input
rlabel metal3 s 107520 8032 108000 8152 6 address[2]
port 2 nsew default input
rlabel metal3 s 107520 10344 108000 10464 6 address[3]
port 3 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_width_0_height_0__pin_0_
port 4 nsew default input
rlabel metal2 s 70766 0 70822 480 6 bottom_width_0_height_0__pin_10_
port 5 nsew default input
rlabel metal2 s 77574 0 77630 480 6 bottom_width_0_height_0__pin_11_
port 6 nsew default tristate
rlabel metal2 s 84290 0 84346 480 6 bottom_width_0_height_0__pin_12_
port 7 nsew default input
rlabel metal2 s 91006 0 91062 480 6 bottom_width_0_height_0__pin_13_
port 8 nsew default tristate
rlabel metal2 s 97814 0 97870 480 6 bottom_width_0_height_0__pin_14_
port 9 nsew default input
rlabel metal2 s 104530 0 104586 480 6 bottom_width_0_height_0__pin_15_
port 10 nsew default tristate
rlabel metal2 s 10046 0 10102 480 6 bottom_width_0_height_0__pin_1_
port 11 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 bottom_width_0_height_0__pin_2_
port 12 nsew default input
rlabel metal2 s 23570 0 23626 480 6 bottom_width_0_height_0__pin_3_
port 13 nsew default tristate
rlabel metal2 s 30286 0 30342 480 6 bottom_width_0_height_0__pin_4_
port 14 nsew default input
rlabel metal2 s 37002 0 37058 480 6 bottom_width_0_height_0__pin_5_
port 15 nsew default tristate
rlabel metal2 s 43810 0 43866 480 6 bottom_width_0_height_0__pin_6_
port 16 nsew default input
rlabel metal2 s 50526 0 50582 480 6 bottom_width_0_height_0__pin_7_
port 17 nsew default tristate
rlabel metal2 s 57334 0 57390 480 6 bottom_width_0_height_0__pin_8_
port 18 nsew default input
rlabel metal2 s 64050 0 64106 480 6 bottom_width_0_height_0__pin_9_
port 19 nsew default tristate
rlabel metal3 s 107520 12656 108000 12776 6 data_in
port 20 nsew default input
rlabel metal3 s 107520 1096 108000 1216 6 enable
port 21 nsew default input
rlabel metal2 s 6734 13520 6790 14000 6 gfpga_pad_GPIO_PAD[0]
port 22 nsew default bidirectional
rlabel metal2 s 20166 13520 20222 14000 6 gfpga_pad_GPIO_PAD[1]
port 23 nsew default bidirectional
rlabel metal2 s 33690 13520 33746 14000 6 gfpga_pad_GPIO_PAD[2]
port 24 nsew default bidirectional
rlabel metal2 s 47214 13520 47270 14000 6 gfpga_pad_GPIO_PAD[3]
port 25 nsew default bidirectional
rlabel metal2 s 60738 13520 60794 14000 6 gfpga_pad_GPIO_PAD[4]
port 26 nsew default bidirectional
rlabel metal2 s 74170 13520 74226 14000 6 gfpga_pad_GPIO_PAD[5]
port 27 nsew default bidirectional
rlabel metal2 s 87694 13520 87750 14000 6 gfpga_pad_GPIO_PAD[6]
port 28 nsew default bidirectional
rlabel metal2 s 101218 13520 101274 14000 6 gfpga_pad_GPIO_PAD[7]
port 29 nsew default bidirectional
rlabel metal4 s 18944 2128 19264 11472 6 vpwr
port 30 nsew default input
rlabel metal4 s 36944 2128 37264 11472 6 vgnd
port 31 nsew default input
<< end >>
