* NGSPICE file created from sb_0__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt sb_0__1_ bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk_0_E_in right_bottom_grid_pin_34_ right_bottom_grid_pin_35_
+ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_
+ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ top_left_grid_pin_1_ VPWR VGND
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_20.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_3.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[4] mux_bottom_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _067_/A sky130_fd_sc_hd__buf_4
X_062_ VGND VGND VPWR VPWR _062_/HI _062_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_114_ chany_bottom_in[10] VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _104_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_1_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ VGND VGND VPWR VPWR _061_/HI _061_/LO sky130_fd_sc_hd__conb_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_26.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_113_ _113_/A VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_mem_bottom_track_1.prog_clk clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_10.mux_l3_in_0_ mux_right_track_10.mux_l2_in_1_/X mux_right_track_10.mux_l2_in_0_/X
+ mux_right_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ VGND VGND VPWR VPWR _060_/HI _060_/LO sky130_fd_sc_hd__conb_1
X_112_ chany_bottom_in[12] VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_10.mux_l2_in_1_ _062_/HI chany_bottom_in[9] mux_right_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xprog_clk_0_FTB00 prog_clk_0_E_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_111_ chany_bottom_in[13] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xmux_right_track_10.mux_l2_in_0_ right_bottom_grid_pin_35_ mux_right_track_10.mux_l1_in_0_/X
+ mux_right_track_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ _046_/HI chany_bottom_in[8] mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l2_in_1_ _047_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_0.mux_l1_in_2_ chany_bottom_in[12] chany_bottom_in[2] mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _117_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_110_ chany_bottom_in[14] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _125_/A sky130_fd_sc_hd__buf_4
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_10.mux_l1_in_0_ chany_top_in[11] chany_top_in[9] mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ right_bottom_grid_pin_34_ mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_22.mux_l2_in_0_ mux_right_track_22.mux_l1_in_1_/X mux_right_track_22.mux_l1_in_0_/X
+ mux_right_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_1_ chanx_right_in[15] chanx_right_in[8] mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_22.mux_l1_in_1_ _036_/HI chany_bottom_in[17] mux_right_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__buf_4
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _089_/A sky130_fd_sc_hd__buf_4
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_18.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_22.mux_l1_in_0_ right_bottom_grid_pin_41_ chany_top_in[17] mux_right_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_0_ chanx_right_in[1] top_left_grid_pin_1_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_34.mux_l2_in_0_ _042_/HI mux_right_track_34.mux_l1_in_0_/X mux_right_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__buf_4
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_1_ _056_/HI chanx_right_in[14] mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_099_ chany_top_in[5] VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_9.mux_l2_in_1_ _060_/HI mux_bottom_track_9.mux_l1_in_2_/X mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__buf_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[16] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__buf_4
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_30.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_34.mux_l1_in_0_ chany_bottom_in[1] right_bottom_grid_pin_39_ mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_098_ chany_top_in[6] VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l1_in_1_ chanx_right_in[7] chanx_right_in[0] mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.mux_l1_in_1_ chanx_right_in[9] chanx_right_in[2] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_28.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l2_in_1_ _048_/HI chany_bottom_in[17] mux_top_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_097_ _097_/A VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_36.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _101_/A sky130_fd_sc_hd__buf_4
XFILLER_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_096_ chany_top_in[8] VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_079_ _079_/A VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_4.mux_l1_in_3_ _044_/HI chany_bottom_in[5] mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_ chany_bottom_in[8] chanx_right_in[19] mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_34.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_095_ chany_top_in[9] VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_078_ _078_/A VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[5] mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_094_ chany_top_in[10] VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_077_ _077_/A VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_1_ _065_/HI chany_bottom_in[13] mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_22.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_093_ _093_/A VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_076_ _076_/A VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_38_ chany_top_in[13] mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[5] chany_top_in[1] mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__buf_4
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_28.mux_l2_in_0_ _039_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_30.mux_l2_in_0_ _040_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_059_ VGND VGND VPWR VPWR _059_/HI _059_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _097_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_1_ _059_/HI mux_bottom_track_5.mux_l1_in_2_/X mux_bottom_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__buf_4
X_092_ chany_top_in[12] VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[17] mux_bottom_track_5.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_075_ _075_/A VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_28.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__buf_4
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ VGND VGND VPWR VPWR _058_/HI _058_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_28.mux_l1_in_0_ chany_bottom_in[11] right_bottom_grid_pin_36_ mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_30.mux_l1_in_0_ chany_bottom_in[7] right_bottom_grid_pin_37_ mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_091_ chany_top_in[13] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_074_ _074_/A VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_1_ chanx_right_in[10] chanx_right_in[3] mux_bottom_track_5.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_26.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
X_057_ VGND VGND VPWR VPWR _057_/HI _057_/LO sky130_fd_sc_hd__conb_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_109_ _109_/A VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ ccff_tail VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_090_ chany_top_in[14] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _103_/A sky130_fd_sc_hd__buf_4
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_33.mux_l1_in_1_ _058_/HI chanx_right_in[13] mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_073_ _073_/A VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_125_ _125_/A VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_056_ VGND VGND VPWR VPWR _056_/HI _056_/LO sky130_fd_sc_hd__conb_1
Xclkbuf_3_1_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_108_ chany_bottom_in[16] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.mux_l2_in_1_ _050_/HI chany_bottom_in[18] mux_top_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_0_ chanx_right_in[6] chany_top_in[10] mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_072_ _072_/A VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_124_ _124_/A VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_12.mux_l3_in_0_ mux_right_track_12.mux_l2_in_1_/X mux_right_track_12.mux_l2_in_0_/X
+ mux_right_track_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_107_ chany_bottom_in[17] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_12.mux_l2_in_1_ _063_/HI chany_bottom_in[10] mux_right_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_1_ _061_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[2] right_bottom_grid_pin_40_ mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l2_in_0_ chany_bottom_in[9] mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_071_ _071_/A VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ _123_/A VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_106_ chany_bottom_in[18] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_12.mux_l2_in_0_ right_bottom_grid_pin_36_ mux_right_track_12.mux_l1_in_0_/X
+ mux_right_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_38_ right_bottom_grid_pin_36_
+ mux_right_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.mux_l2_in_1_ _037_/HI chany_bottom_in[19] mux_right_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ _049_/HI chany_bottom_in[13] mux_top_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_070_ _070_/A VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _113_/A sky130_fd_sc_hd__buf_4
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_122_ chany_bottom_in[2] VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[6] mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_105_ _105_/A VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__buf_4
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_12.mux_l1_in_0_ chany_top_in[15] chany_top_in[10] mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_34_ chany_top_in[2] mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_24.mux_l2_in_0_ chany_bottom_in[18] mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _124_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_1_ chany_bottom_in[4] chanx_right_in[16] mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_121_ _121_/A VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_1_ _054_/HI mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_104_ _104_/A VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__buf_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[19] mux_bottom_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_34_ chany_top_in[18] mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_0_ chanx_right_in[9] chanx_right_in[2] mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_120_ chany_bottom_in[4] VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_36.mux_l2_in_0_ _043_/HI mux_right_track_36.mux_l1_in_0_/X mux_right_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_30.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_103_ _103_/A VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l1_in_1_ chanx_right_in[12] chanx_right_in[5] mux_bottom_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _068_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _071_/A sky130_fd_sc_hd__buf_4
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _105_/A sky130_fd_sc_hd__buf_4
X_102_ chany_top_in[2] VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xmux_right_track_36.mux_l1_in_0_ chany_bottom_in[0] right_bottom_grid_pin_40_ mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_101_ _101_/A VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_100_ chany_top_in[4] VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_mem_bottom_track_1.prog_clk clkbuf_1_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l1_in_3_ _045_/HI chany_bottom_in[6] mux_right_track_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_32.mux_l2_in_1_ _051_/HI chany_bottom_in[10] mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_1_ mux_right_track_6.mux_l1_in_3_/X mux_right_track_6.mux_l1_in_2_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l1_in_2_ right_bottom_grid_pin_41_ right_bottom_grid_pin_39_
+ mux_right_track_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_32.mux_l2_in_0_ chanx_right_in[14] mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_18.mux_l2_in_0_ mux_right_track_18.mux_l1_in_1_/X mux_right_track_18.mux_l1_in_0_/X
+ mux_right_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_089_ _089_/A VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_20.mux_l2_in_0_ mux_right_track_20.mux_l1_in_1_/X mux_right_track_20.mux_l1_in_0_/X
+ mux_right_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.mux_l1_in_1_ _033_/HI chany_bottom_in[14] mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l1_in_1_ right_bottom_grid_pin_37_ right_bottom_grid_pin_35_
+ mux_right_track_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_20.mux_l1_in_1_ _035_/HI chany_bottom_in[16] mux_right_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l2_in_1_ _053_/HI mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_ chany_bottom_in[16] chany_bottom_in[6] mux_top_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_32.mux_l1_in_0_ chanx_right_in[7] chanx_right_in[0] mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_088_ chany_top_in[16] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_18.mux_l1_in_0_ right_bottom_grid_pin_39_ chany_top_in[14] mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_6.mux_l1_in_0_ chany_top_in[6] chany_top_in[3] mux_right_track_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l1_in_0_ right_bottom_grid_pin_40_ chany_top_in[16] mux_right_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _093_/A sky130_fd_sc_hd__buf_4
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_36.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__buf_4
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_32.mux_l2_in_0_ _041_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _121_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_8.mux_l1_in_1_ chanx_right_in[18] chanx_right_in[11] mux_top_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _070_/A sky130_fd_sc_hd__buf_4
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_087_ chany_top_in[17] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__buf_4
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[4] top_left_grid_pin_1_ mux_top_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_0_0_mem_bottom_track_1.prog_clk clkbuf_1_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.mux_l1_in_0_ chany_bottom_in[3] right_bottom_grid_pin_38_ mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_086_ chany_top_in[18] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ _069_/A VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ _085_/A VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_068_ _068_/A VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l1_in_3_ _034_/HI chany_bottom_in[4] mux_right_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_084_ _084_/A VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ _067_/A VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_119_ chany_bottom_in[5] VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_14.mux_l3_in_0_ mux_right_track_14.mux_l2_in_1_/X mux_right_track_14.mux_l2_in_0_/X
+ mux_right_track_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_0 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_14.mux_l2_in_1_ _064_/HI chany_bottom_in[12] mux_right_track_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l1_in_2_ right_bottom_grid_pin_41_ right_bottom_grid_pin_39_
+ mux_right_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
X_083_ _083_/A VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_066_ right_bottom_grid_pin_41_ VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_34.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_118_ chany_bottom_in[6] VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l1_in_1_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_14.mux_l2_in_0_ right_bottom_grid_pin_37_ mux_right_track_14.mux_l1_in_0_/X
+ mux_right_track_14.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_082_ _082_/A VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_37_ right_bottom_grid_pin_35_
+ mux_right_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _109_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_4.mux_l2_in_1_ _052_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ VGND VGND VPWR VPWR _065_/HI _065_/LO sky130_fd_sc_hd__conb_1
Xclkbuf_3_5_0_mem_bottom_track_1.prog_clk clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_117_ _117_/A VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xmux_top_track_4.mux_l1_in_2_ chany_bottom_in[14] chany_bottom_in[5] mux_top_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_14.mux_l1_in_0_ chany_top_in[19] chany_top_in[12] mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_081_ _081_/A VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__buf_4
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[4] chany_top_in[0] mux_right_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_26.mux_l2_in_0_ _038_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_064_ VGND VGND VPWR VPWR _064_/HI _064_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _123_/A sky130_fd_sc_hd__buf_4
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_17.mux_l2_in_1_ _055_/HI chanx_right_in[15] mux_bottom_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_1_ chanx_right_in[17] chanx_right_in[10] mux_top_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_116_ chany_bottom_in[8] VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l2_in_1_ _057_/HI chanx_right_in[18] mux_bottom_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__buf_4
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__buf_4
X_080_ _080_/A VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XFILLER_10_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_063_ VGND VGND VPWR VPWR _063_/HI _063_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_0_ chanx_right_in[3] top_left_grid_pin_1_ mux_top_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ chany_bottom_in[9] VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_26.mux_l1_in_0_ chany_bottom_in[15] right_bottom_grid_pin_35_ mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ chanx_right_in[8] chanx_right_in[1] mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

