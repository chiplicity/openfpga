* NGSPICE file created from cbx_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

.subckt cbx_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_14_ top_grid_pin_2_ top_grid_pin_6_ vpwr vgnd
XFILLER_22_144 vpwr vgnd scs8hd_fill_2
XFILLER_22_166 vgnd vpwr scs8hd_decap_8
XFILLER_7_7 vgnd vpwr scs8hd_decap_8
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_188 vgnd vpwr scs8hd_decap_3
XFILLER_3_23 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _111_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_103 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__108__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _117_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_3_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _041_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_20 vpwr vgnd scs8hd_fill_2
XFILLER_15_217 vgnd vpwr scs8hd_decap_12
X_131_ _131_/HI _131_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_31 vpwr vgnd scs8hd_fill_2
X_062_ address[4] _122_/B _069_/C _062_/X vgnd vpwr scs8hd_or3_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_9 vgnd vpwr scs8hd_fill_1
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_66 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_045_ address[6] _083_/A vgnd vpwr scs8hd_inv_8
XANTENNA__105__C address[5] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_5.LATCH_0_.latch data_in mem_top_ipin_5.LATCH_0_.latch/Q _090_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_114_ _075_/A _111_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _136_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_205 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_43 vpwr vgnd scs8hd_fill_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_7.LATCH_3_.latch data_in mem_top_ipin_7.LATCH_3_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__116__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_45 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_109 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _129_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_4
XFILLER_19_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB _053_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_186 vgnd vpwr scs8hd_fill_1
XANTENNA__042__A address[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_25_164 vpwr vgnd scs8hd_fill_2
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_186 vgnd vpwr scs8hd_decap_4
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_123 vgnd vpwr scs8hd_decap_8
XFILLER_9_127 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_108 vgnd vpwr scs8hd_decap_4
XFILLER_10_137 vpwr vgnd scs8hd_fill_2
XFILLER_12_22 vgnd vpwr scs8hd_decap_8
XFILLER_12_44 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XANTENNA__108__C _122_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_141 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _122_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__140__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA__050__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _130_/HI _130_/LO vgnd vpwr scs8hd_conb_1
XFILLER_15_229 vgnd vpwr scs8hd_decap_4
XFILLER_23_98 vpwr vgnd scs8hd_fill_2
XFILLER_23_87 vpwr vgnd scs8hd_fill_2
XFILLER_23_76 vpwr vgnd scs8hd_fill_2
X_061_ _051_/B _075_/A _061_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_199 vgnd vpwr scs8hd_decap_4
XFILLER_2_166 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_47 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vgnd vpwr scs8hd_decap_4
XFILLER_20_232 vgnd vpwr scs8hd_fill_1
XANTENNA__045__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_3
XFILLER_11_232 vgnd vpwr scs8hd_fill_1
X_113_ _120_/A _111_/B _113_/Y vgnd vpwr scs8hd_nor2_4
X_044_ enable _098_/C vgnd vpwr scs8hd_inv_8
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_55 vgnd vpwr scs8hd_decap_3
XFILLER_28_184 vgnd vpwr scs8hd_fill_1
XFILLER_6_68 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_143 vgnd vpwr scs8hd_decap_4
XFILLER_25_132 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_ipin_3.LATCH_3_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_31_43 vpwr vgnd scs8hd_fill_2
XFILLER_16_110 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _122_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_143 vgnd vpwr scs8hd_decap_8
XFILLER_16_154 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__143__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__053__A _051_/B vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _124_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_117 vgnd vpwr scs8hd_decap_3
XFILLER_13_102 vpwr vgnd scs8hd_fill_2
XFILLER_13_113 vgnd vpwr scs8hd_decap_4
XFILLER_13_157 vgnd vpwr scs8hd_decap_3
XFILLER_13_179 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__048__A address[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_205 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_7.LATCH_4_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_5_197 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__050__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_44 vpwr vgnd scs8hd_fill_2
XFILLER_23_11 vgnd vpwr scs8hd_decap_3
XFILLER_3_3 vgnd vpwr scs8hd_decap_4
X_060_ address[1] address[2] address[0] _075_/A vgnd vpwr scs8hd_or3_4
XFILLER_2_145 vgnd vpwr scs8hd_decap_6
XFILLER_2_178 vpwr vgnd scs8hd_fill_2
XFILLER_9_13 vpwr vgnd scs8hd_fill_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vgnd vpwr scs8hd_decap_4
XANTENNA__151__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__061__A _051_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vgnd vpwr scs8hd_decap_3
XFILLER_18_44 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
XFILLER_34_76 vgnd vpwr scs8hd_fill_1
X_043_ address[2] _043_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_200 vpwr vgnd scs8hd_fill_2
X_112_ _119_/A _111_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _137_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__056__A _056_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB _077_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_8
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_0_.latch data_in mem_top_ipin_1.LATCH_0_.latch/Q _061_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_232 vgnd vpwr scs8hd_fill_1
XFILLER_16_122 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_ipin_3.LATCH_3_.latch data_in mem_top_ipin_3.LATCH_3_.latch/Q _072_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__053__B _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_66 vgnd vpwr scs8hd_decap_3
XFILLER_26_88 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_184 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__048__B _043_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__064__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_57 vpwr vgnd scs8hd_fill_2
XFILLER_33_209 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_0_.latch data_in _041_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_154 vpwr vgnd scs8hd_fill_2
XANTENNA__149__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__050__C _069_/C vgnd vpwr scs8hd_diode_2
XANTENNA__059__A _051_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_124 vgnd vpwr scs8hd_fill_1
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_9_25 vgnd vpwr scs8hd_fill_1
XFILLER_14_231 vpwr vgnd scs8hd_fill_2
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_3_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__061__B _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_8
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_042_ address[1] _056_/A vgnd vpwr scs8hd_inv_8
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_111_ _118_/A _111_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_92 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_208 vgnd vpwr scs8hd_decap_3
XANTENNA__056__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_13 vgnd vpwr scs8hd_fill_1
XFILLER_29_33 vpwr vgnd scs8hd_fill_2
XFILLER_29_99 vpwr vgnd scs8hd_fill_2
XFILLER_29_77 vgnd vpwr scs8hd_decap_4
XFILLER_29_55 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_3
XFILLER_20_7 vgnd vpwr scs8hd_decap_6
XFILLER_34_178 vgnd vpwr scs8hd_decap_8
XANTENNA__157__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_153 vgnd vpwr scs8hd_decap_6
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A _120_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_6.LATCH_2_.latch data_in mem_top_ipin_6.LATCH_2_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_67 vpwr vgnd scs8hd_fill_2
XFILLER_31_23 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_4_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_0_222 vpwr vgnd scs8hd_fill_2
XFILLER_0_200 vpwr vgnd scs8hd_fill_2
XFILLER_31_115 vgnd vpwr scs8hd_decap_6
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_159 vgnd vpwr scs8hd_decap_4
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _040_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
XFILLER_22_148 vgnd vpwr scs8hd_decap_4
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XFILLER_26_45 vgnd vpwr scs8hd_decap_12
XFILLER_3_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_130 vpwr vgnd scs8hd_fill_2
XFILLER_12_170 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB _075_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__048__C _058_/C vgnd vpwr scs8hd_diode_2
XANTENNA__064__B _062_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_107 vgnd vpwr scs8hd_fill_1
XANTENNA__080__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_221 vgnd vpwr scs8hd_decap_12
XANTENNA__059__B _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_48 vgnd vpwr scs8hd_decap_3
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _117_/A _111_/B _110_/Y vgnd vpwr scs8hd_nor2_4
X_041_ _041_/A _041_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _129_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _138_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__056__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__072__B _072_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _059_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_47 vgnd vpwr scs8hd_decap_8
XFILLER_20_69 vpwr vgnd scs8hd_fill_2
XFILLER_28_176 vgnd vpwr scs8hd_decap_8
XFILLER_28_165 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_231 vpwr vgnd scs8hd_fill_2
XFILLER_13_7 vgnd vpwr scs8hd_fill_1
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XFILLER_25_168 vgnd vpwr scs8hd_decap_4
XANTENNA__067__B _062_/X vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XFILLER_0_212 vgnd vpwr scs8hd_decap_4
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_135 vpwr vgnd scs8hd_fill_2
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_57 vgnd vpwr scs8hd_fill_1
XANTENNA__078__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_138 vpwr vgnd scs8hd_fill_2
XFILLER_13_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_ipin_1.LATCH_3_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_182 vgnd vpwr scs8hd_fill_1
XFILLER_35_230 vgnd vpwr scs8hd_decap_3
XFILLER_27_219 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_119 vgnd vpwr scs8hd_decap_3
XANTENNA__080__B _080_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_219 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_5_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_60 vgnd vpwr scs8hd_fill_1
XANTENNA__075__B _072_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__091__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_14_200 vpwr vgnd scs8hd_fill_2
XFILLER_13_91 vpwr vgnd scs8hd_fill_2
XFILLER_1_170 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_4_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_18_69 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_8
XFILLER_7_207 vgnd vpwr scs8hd_fill_1
XANTENNA__086__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_040_ _040_/A _040_/Y vgnd vpwr scs8hd_inv_8
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_133 vgnd vpwr scs8hd_decap_3
XFILLER_6_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_31_47 vpwr vgnd scs8hd_fill_2
XANTENNA__083__B address[5] vgnd vpwr scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_15_180 vgnd vpwr scs8hd_fill_1
XFILLER_7_60 vgnd vpwr scs8hd_fill_1
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__078__B _080_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_106 vpwr vgnd scs8hd_fill_2
XFILLER_13_117 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_2_.latch data_in mem_top_ipin_2.LATCH_2_.latch/Q _066_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_194 vpwr vgnd scs8hd_fill_2
XFILLER_8_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_176 vgnd vpwr scs8hd_decap_8
XFILLER_8_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_38 vgnd vpwr scs8hd_decap_4
XANTENNA__089__A _120_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_5_.latch data_in mem_top_ipin_4.LATCH_5_.latch/Q _077_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_27_90 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_72 vpwr vgnd scs8hd_fill_2
XFILLER_4_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_48 vgnd vpwr scs8hd_decap_3
XFILLER_3_7 vgnd vpwr scs8hd_fill_1
XFILLER_2_127 vpwr vgnd scs8hd_fill_2
XANTENNA__091__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__086__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_48 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_219 vpwr vgnd scs8hd_fill_2
XFILLER_11_204 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_099_ _116_/A _104_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _139_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_4
XANTENNA__097__A _075_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_10_60 vgnd vpwr scs8hd_decap_4
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XFILLER_19_101 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_192 vpwr vgnd scs8hd_fill_2
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_107 vpwr vgnd scs8hd_fill_2
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_81 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_15_170 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_5.LATCH_1_.latch data_in mem_top_ipin_5.LATCH_1_.latch/Q _089_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA__094__B _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_151 vpwr vgnd scs8hd_fill_2
XFILLER_3_19 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_4_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_4_.latch data_in mem_top_ipin_7.LATCH_4_.latch/Q _100_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB _065_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_210 vgnd vpwr scs8hd_decap_4
XFILLER_5_158 vpwr vgnd scs8hd_fill_2
XFILLER_17_221 vpwr vgnd scs8hd_fill_2
XFILLER_4_84 vgnd vpwr scs8hd_decap_6
XFILLER_4_40 vgnd vpwr scs8hd_fill_1
XFILLER_23_27 vpwr vgnd scs8hd_fill_2
XFILLER_23_16 vpwr vgnd scs8hd_fill_2
XFILLER_2_106 vgnd vpwr scs8hd_decap_3
XANTENNA__091__C _098_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_216 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_24_70 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_098_ _122_/A address[3] _098_/C _084_/D _104_/B vgnd vpwr scs8hd_or4_4
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_29_37 vpwr vgnd scs8hd_fill_2
XFILLER_28_113 vgnd vpwr scs8hd_decap_3
XANTENNA__097__B _091_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_83 vgnd vpwr scs8hd_decap_6
XFILLER_19_113 vpwr vgnd scs8hd_fill_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_182 vgnd vpwr scs8hd_fill_1
XFILLER_15_17 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_226 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
XFILLER_22_108 vgnd vpwr scs8hd_decap_4
XFILLER_30_185 vpwr vgnd scs8hd_fill_2
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_123 vgnd vpwr scs8hd_fill_1
XFILLER_8_134 vpwr vgnd scs8hd_fill_2
XFILLER_8_145 vpwr vgnd scs8hd_fill_2
XFILLER_12_130 vpwr vgnd scs8hd_fill_2
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_137 vpwr vgnd scs8hd_fill_2
XFILLER_4_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__091__D _084_/D vgnd vpwr scs8hd_diode_2
XFILLER_13_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
XFILLER_6_210 vgnd vpwr scs8hd_fill_1
X_097_ _075_/A _091_/X _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_232 vgnd vpwr scs8hd_fill_1
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XFILLER_1_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _131_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_ipin_3.LATCH_4_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
X_149_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_28 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_139 vpwr vgnd scs8hd_fill_2
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_94 vpwr vgnd scs8hd_fill_2
XFILLER_30_120 vgnd vpwr scs8hd_decap_3
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_52 vgnd vpwr scs8hd_decap_6
Xmux_top_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_120 vpwr vgnd scs8hd_fill_2
XFILLER_21_164 vpwr vgnd scs8hd_fill_2
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _139_/HI mem_top_ipin_7.LATCH_5_.latch/Q
+ mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_12_ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_1.LATCH_1_.latch data_in mem_top_ipin_1.LATCH_1_.latch/Q _059_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_116 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_60 vgnd vpwr scs8hd_fill_1
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_204 vgnd vpwr scs8hd_decap_6
Xmem_top_ipin_3.LATCH_4_.latch data_in mem_top_ipin_3.LATCH_4_.latch/Q _071_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_204 vgnd vpwr scs8hd_decap_8
XFILLER_13_51 vgnd vpwr scs8hd_decap_4
XFILLER_13_62 vgnd vpwr scs8hd_fill_1
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
XFILLER_1_174 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _117_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
X_096_ _120_/A _091_/X _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_21 vgnd vpwr scs8hd_fill_1
XFILLER_1_54 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_1_.latch data_in _040_/A _106_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_104 vpwr vgnd scs8hd_fill_2
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XFILLER_19_94 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
X_148_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_079_ _118_/A _080_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_8
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_62 vpwr vgnd scs8hd_fill_2
XFILLER_11_9 vpwr vgnd scs8hd_fill_2
XFILLER_30_165 vgnd vpwr scs8hd_fill_1
XFILLER_30_110 vgnd vpwr scs8hd_fill_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_75 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XFILLER_29_232 vgnd vpwr scs8hd_fill_1
XFILLER_12_143 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vgnd vpwr scs8hd_fill_1
XFILLER_16_73 vpwr vgnd scs8hd_fill_2
XFILLER_16_84 vgnd vpwr scs8hd_decap_8
XFILLER_32_72 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_169 vgnd vpwr scs8hd_decap_4
XFILLER_12_198 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_4.LATCH_0_.latch data_in mem_top_ipin_4.LATCH_0_.latch/Q _082_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__103__A _120_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_6
Xmem_top_ipin_6.LATCH_3_.latch data_in mem_top_ipin_6.LATCH_3_.latch/Q _094_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_76 vgnd vpwr scs8hd_decap_3
XFILLER_4_54 vgnd vpwr scs8hd_decap_6
XFILLER_4_32 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_4_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_1_131 vgnd vpwr scs8hd_decap_3
XANTENNA__100__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_197 vpwr vgnd scs8hd_fill_2
XFILLER_1_153 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_24_62 vpwr vgnd scs8hd_fill_2
X_095_ _119_/A _091_/X _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_33 vgnd vpwr scs8hd_decap_4
XANTENNA__111__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_149 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _138_/HI mem_top_ipin_6.LATCH_5_.latch/Q
+ mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_64 vgnd vpwr scs8hd_fill_1
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XFILLER_19_149 vpwr vgnd scs8hd_fill_2
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
X_147_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__106__A address[4] vgnd vpwr scs8hd_diode_2
X_078_ _117_/A _080_/B _078_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_3 vgnd vpwr scs8hd_decap_8
XFILLER_33_130 vgnd vpwr scs8hd_decap_12
XFILLER_18_182 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_163 vgnd vpwr scs8hd_decap_3
XFILLER_24_130 vgnd vpwr scs8hd_decap_6
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_199 vgnd vpwr scs8hd_decap_12
XFILLER_30_177 vgnd vpwr scs8hd_decap_8
XFILLER_15_174 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _068_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_126 vpwr vgnd scs8hd_fill_2
XFILLER_12_166 vpwr vgnd scs8hd_fill_2
XFILLER_32_84 vgnd vpwr scs8hd_decap_8
XANTENNA__103__B _104_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_170 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_73 vgnd vpwr scs8hd_decap_4
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_225 vgnd vpwr scs8hd_decap_8
XFILLER_4_173 vgnd vpwr scs8hd_decap_8
XANTENNA__114__A _075_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _116_/A vgnd vpwr scs8hd_diode_2
X_094_ _118_/A _091_/X _094_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_202 vgnd vpwr scs8hd_decap_8
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__111__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_19 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_21 vgnd vpwr scs8hd_decap_8
XFILLER_27_150 vgnd vpwr scs8hd_decap_4
XFILLER_19_117 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_146_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__106__B _122_/B vgnd vpwr scs8hd_diode_2
X_077_ _116_/A _080_/B _077_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_142 vgnd vpwr scs8hd_decap_12
XFILLER_25_109 vgnd vpwr scs8hd_decap_3
XFILLER_18_172 vgnd vpwr scs8hd_fill_1
XFILLER_18_194 vgnd vpwr scs8hd_fill_1
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_42 vgnd vpwr scs8hd_decap_3
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_142 vpwr vgnd scs8hd_fill_2
XFILLER_15_153 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_1.LATCH_4_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_30_189 vgnd vpwr scs8hd_fill_1
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_33 vpwr vgnd scs8hd_fill_2
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_129_ _129_/HI _129_/LO vgnd vpwr scs8hd_conb_1
XFILLER_21_112 vpwr vgnd scs8hd_fill_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_29_212 vgnd vpwr scs8hd_decap_12
XFILLER_32_52 vgnd vpwr scs8hd_decap_12
XFILLER_8_149 vgnd vpwr scs8hd_decap_4
XFILLER_16_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_108 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _137_/HI mem_top_ipin_5.LATCH_5_.latch/Q
+ mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _128_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__040__A _040_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_10 vgnd vpwr scs8hd_fill_1
XFILLER_13_76 vpwr vgnd scs8hd_fill_2
XFILLER_1_111 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _118_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_3_.latch data_in mem_top_ipin_2.LATCH_3_.latch/Q _065_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_093_ _117_/A _091_/X _093_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_129 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_99 vpwr vgnd scs8hd_fill_2
XFILLER_19_20 vgnd vpwr scs8hd_decap_3
XFILLER_19_53 vgnd vpwr scs8hd_fill_1
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_145_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__106__C _122_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_076_ _122_/A _122_/B _069_/C _080_/B vgnd vpwr scs8hd_or3_4
XANTENNA__122__B _122_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_33_198 vpwr vgnd scs8hd_fill_2
XFILLER_33_154 vgnd vpwr scs8hd_decap_12
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_198 vgnd vpwr scs8hd_decap_12
XFILLER_24_187 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_98 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_30_157 vgnd vpwr scs8hd_decap_8
XANTENNA__117__B _118_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
X_128_ _075_/A _122_/X _128_/Y vgnd vpwr scs8hd_nor2_4
X_059_ _051_/B _120_/A _059_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_168 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XANTENNA__043__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_224 vgnd vpwr scs8hd_decap_8
XFILLER_12_102 vgnd vpwr scs8hd_decap_12
XFILLER_16_10 vgnd vpwr scs8hd_decap_4
XFILLER_16_21 vgnd vpwr scs8hd_fill_1
XFILLER_16_43 vpwr vgnd scs8hd_fill_2
XFILLER_16_54 vgnd vpwr scs8hd_decap_8
XFILLER_32_64 vgnd vpwr scs8hd_decap_8
XANTENNA__128__A _075_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_227 vgnd vpwr scs8hd_decap_6
XFILLER_27_86 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vgnd vpwr scs8hd_fill_1
XFILLER_27_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_208 vgnd vpwr scs8hd_decap_6
XFILLER_4_142 vgnd vpwr scs8hd_decap_3
XFILLER_4_197 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_230 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_219 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_5.LATCH_2_.latch data_in mem_top_ipin_5.LATCH_2_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_178 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA__141__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__051__A _116_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_5_.latch data_in mem_top_ipin_7.LATCH_5_.latch/Q _099_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_24_87 vgnd vpwr scs8hd_decap_4
XFILLER_24_43 vgnd vpwr scs8hd_decap_8
XFILLER_10_211 vgnd vpwr scs8hd_decap_3
X_092_ _116_/A _091_/X _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_58 vgnd vpwr scs8hd_decap_3
XFILLER_1_69 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_108 vgnd vpwr scs8hd_decap_3
XANTENNA__046__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_45 vpwr vgnd scs8hd_fill_2
XFILLER_10_67 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_89 vgnd vpwr scs8hd_fill_1
XFILLER_19_32 vpwr vgnd scs8hd_fill_2
XFILLER_19_98 vgnd vpwr scs8hd_fill_1
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
X_075_ _075_/A _072_/B _075_/Y vgnd vpwr scs8hd_nor2_4
X_144_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__106__D _058_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__122__C _122_/C vgnd vpwr scs8hd_diode_2
XFILLER_33_111 vpwr vgnd scs8hd_fill_2
XFILLER_33_166 vgnd vpwr scs8hd_decap_12
XFILLER_24_111 vgnd vpwr scs8hd_decap_12
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_11 vgnd vpwr scs8hd_decap_12
XFILLER_21_66 vpwr vgnd scs8hd_fill_2
XFILLER_21_77 vpwr vgnd scs8hd_fill_2
XFILLER_30_125 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _136_/HI mem_top_ipin_4.LATCH_5_.latch/Q
+ mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_166 vpwr vgnd scs8hd_fill_2
X_058_ address[1] address[2] _058_/C _120_/A vgnd vpwr scs8hd_or3_4
X_127_ _120_/A _122_/X _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_147 vpwr vgnd scs8hd_fill_2
XFILLER_12_114 vgnd vpwr scs8hd_fill_1
XFILLER_12_147 vgnd vpwr scs8hd_decap_6
XFILLER_16_77 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB _055_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_98 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__144__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_fill_1
XFILLER_7_184 vpwr vgnd scs8hd_fill_2
XANTENNA__054__A _056_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_43 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_4
XFILLER_4_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__049__A enable vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__051__B _051_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_11 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_66 vpwr vgnd scs8hd_fill_2
X_091_ address[4] _122_/B _098_/C _084_/D _091_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_6
XANTENNA__152__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_3_219 vgnd vpwr scs8hd_decap_12
XANTENNA__062__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_79 vpwr vgnd scs8hd_fill_2
XFILLER_19_11 vgnd vpwr scs8hd_decap_3
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
XFILLER_27_175 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_074_ _120_/A _072_/B _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_101 vgnd vpwr scs8hd_decap_6
XFILLER_18_131 vgnd vpwr scs8hd_decap_3
XFILLER_18_197 vgnd vpwr scs8hd_fill_1
XFILLER_33_178 vgnd vpwr scs8hd_decap_4
XANTENNA__147__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vgnd vpwr scs8hd_decap_4
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__057__A _051_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_4
XFILLER_30_137 vgnd vpwr scs8hd_decap_12
X_126_ _119_/A _122_/X _126_/Y vgnd vpwr scs8hd_nor2_4
X_057_ _051_/B _119_/A _057_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_108 vgnd vpwr scs8hd_decap_8
XFILLER_8_119 vgnd vpwr scs8hd_decap_4
XFILLER_12_126 vpwr vgnd scs8hd_fill_2
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XFILLER_7_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_109_ _116_/A _111_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__054__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_4
XANTENNA__155__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__049__B _083_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__065__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_24 vpwr vgnd scs8hd_fill_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _135_/HI mem_top_ipin_3.LATCH_5_.latch/Q
+ mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_8
X_090_ _075_/A _088_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_2_.latch data_in mem_top_ipin_1.LATCH_2_.latch/Q _057_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__062__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_165 vpwr vgnd scs8hd_fill_2
XFILLER_19_45 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vpwr vgnd scs8hd_fill_2
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
X_142_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_3.LATCH_5_.latch data_in mem_top_ipin_3.LATCH_5_.latch/Q _070_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_073_ _119_/A _072_/B _073_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_165 vgnd vpwr scs8hd_fill_1
XFILLER_24_168 vgnd vpwr scs8hd_decap_8
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__057__B _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA__073__A _119_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_15_113 vpwr vgnd scs8hd_fill_2
XFILLER_30_149 vgnd vpwr scs8hd_decap_4
XFILLER_7_15 vgnd vpwr scs8hd_fill_1
XFILLER_7_48 vpwr vgnd scs8hd_fill_2
X_125_ _118_/A _122_/X _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_7 vgnd vpwr scs8hd_decap_12
X_056_ _056_/A address[2] address[0] _119_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_116 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_24 vgnd vpwr scs8hd_decap_4
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
X_108_ address[4] address[3] _122_/C _111_/B vgnd vpwr scs8hd_or3_4
X_039_ address[0] _058_/C vgnd vpwr scs8hd_inv_8
XANTENNA__070__B _072_/B vgnd vpwr scs8hd_diode_2
XANTENNA__054__C _058_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_56 vpwr vgnd scs8hd_fill_2
XFILLER_16_230 vgnd vpwr scs8hd_decap_3
XFILLER_31_222 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__049__C address[5] vgnd vpwr scs8hd_diode_2
XFILLER_22_200 vgnd vpwr scs8hd_decap_6
XANTENNA__065__B _062_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_47 vpwr vgnd scs8hd_fill_2
XFILLER_1_159 vpwr vgnd scs8hd_fill_2
XFILLER_1_115 vgnd vpwr scs8hd_decap_4
XANTENNA__081__A _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_204 vpwr vgnd scs8hd_fill_2
XFILLER_13_200 vpwr vgnd scs8hd_fill_2
XFILLER_0_170 vgnd vpwr scs8hd_decap_4
XFILLER_5_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB _063_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_1_.latch data_in mem_top_ipin_4.LATCH_1_.latch/Q _081_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_203 vgnd vpwr scs8hd_decap_8
XANTENNA__076__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_6.LATCH_4_.latch data_in mem_top_ipin_6.LATCH_4_.latch/Q _093_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__062__C _069_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XFILLER_27_188 vpwr vgnd scs8hd_fill_2
X_141_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
X_072_ _118_/A _072_/B _072_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_82 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_25 vpwr vgnd scs8hd_fill_2
XFILLER_21_47 vpwr vgnd scs8hd_fill_2
XANTENNA__073__B _072_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_106 vgnd vpwr scs8hd_decap_4
X_124_ _117_/A _122_/X _124_/Y vgnd vpwr scs8hd_nor2_4
X_055_ _051_/B _118_/A _055_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_128 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__068__B _062_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_47 vgnd vpwr scs8hd_decap_4
XFILLER_32_35 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__084__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_194 vgnd vpwr scs8hd_fill_1
X_107_ address[4] _122_/B _122_/C address[0] _107_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_11_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _134_/HI mem_top_ipin_2.LATCH_5_.latch/Q
+ mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_81 vgnd vpwr scs8hd_decap_8
XFILLER_27_24 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_209 vgnd vpwr scs8hd_decap_8
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__081__B _080_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_7.LATCH_0_.latch data_in mem_top_ipin_7.LATCH_0_.latch/Q _104_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_212 vgnd vpwr scs8hd_decap_3
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_0_160 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA__076__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_49 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vgnd vpwr scs8hd_decap_3
XANTENNA__087__A _118_/A vgnd vpwr scs8hd_diode_2
X_071_ _117_/A _072_/B _071_/Y vgnd vpwr scs8hd_nor2_4
X_140_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_18_123 vgnd vpwr scs8hd_decap_6
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_33_126 vpwr vgnd scs8hd_fill_2
XFILLER_33_115 vgnd vpwr scs8hd_decap_6
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
X_054_ _056_/A address[2] _058_/C _118_/A vgnd vpwr scs8hd_or3_4
X_123_ _116_/A _122_/X _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _061_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__084__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_162 vgnd vpwr scs8hd_fill_1
X_106_ address[4] _122_/B _122_/C _058_/C _106_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_133 vgnd vpwr scs8hd_decap_3
XFILLER_7_166 vpwr vgnd scs8hd_fill_2
XFILLER_7_199 vgnd vpwr scs8hd_decap_8
XFILLER_11_184 vpwr vgnd scs8hd_fill_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_47 vgnd vpwr scs8hd_decap_6
XFILLER_25_232 vgnd vpwr scs8hd_fill_1
XANTENNA__079__B _080_/B vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _119_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_147 vgnd vpwr scs8hd_decap_6
XFILLER_4_125 vpwr vgnd scs8hd_fill_2
XFILLER_4_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_217 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_150 vgnd vpwr scs8hd_decap_3
XANTENNA__092__B _091_/X vgnd vpwr scs8hd_diode_2
XANTENNA__076__C _069_/C vgnd vpwr scs8hd_diode_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_220 vpwr vgnd scs8hd_fill_2
XFILLER_14_70 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_135 vpwr vgnd scs8hd_fill_2
XFILLER_27_146 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _088_/B vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ _116_/A _072_/B _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _133_/HI mem_top_ipin_1.LATCH_5_.latch/Q
+ mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_102 vgnd vpwr scs8hd_fill_1
XFILLER_18_113 vgnd vpwr scs8hd_fill_1
XFILLER_18_157 vgnd vpwr scs8hd_decap_8
XFILLER_18_168 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_4_.latch data_in mem_top_ipin_2.LATCH_4_.latch/Q _064_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__098__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
XFILLER_23_160 vgnd vpwr scs8hd_decap_4
XFILLER_15_138 vpwr vgnd scs8hd_fill_2
XFILLER_15_149 vpwr vgnd scs8hd_fill_2
XFILLER_7_29 vpwr vgnd scs8hd_fill_2
X_122_ _122_/A _122_/B _122_/C _122_/X vgnd vpwr scs8hd_or3_4
X_053_ _051_/B _117_/A _053_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_193 vpwr vgnd scs8hd_fill_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__084__C _098_/C vgnd vpwr scs8hd_diode_2
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_20_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_fill_1
X_105_ _098_/C address[6] address[5] _122_/C vgnd vpwr scs8hd_or3_4
XFILLER_7_156 vgnd vpwr scs8hd_fill_1
XFILLER_11_174 vgnd vpwr scs8hd_decap_6
XFILLER_22_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_8_50 vgnd vpwr scs8hd_decap_8
XFILLER_8_61 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__095__B _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vpwr vgnd scs8hd_fill_2
XFILLER_4_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_28 vgnd vpwr scs8hd_decap_8
XFILLER_1_107 vpwr vgnd scs8hd_fill_2
XFILLER_9_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_4
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XFILLER_30_70 vgnd vpwr scs8hd_fill_1
XFILLER_5_232 vgnd vpwr scs8hd_fill_1
Xmem_top_ipin_3.LATCH_0_.latch data_in mem_top_ipin_3.LATCH_0_.latch/Q _075_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_29 vpwr vgnd scs8hd_fill_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_27_103 vpwr vgnd scs8hd_fill_2
XFILLER_19_16 vpwr vgnd scs8hd_fill_2
XFILLER_19_49 vgnd vpwr scs8hd_decap_4
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_27_169 vgnd vpwr scs8hd_decap_4
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vgnd vpwr scs8hd_decap_4
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_ipin_5.LATCH_3_.latch data_in mem_top_ipin_5.LATCH_3_.latch/Q _087_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XFILLER_2_52 vgnd vpwr scs8hd_decap_4
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_191 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__098__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_15_117 vgnd vpwr scs8hd_decap_3
X_121_ _075_/A _118_/B _121_/Y vgnd vpwr scs8hd_nor2_4
X_052_ address[1] _043_/Y address[0] _117_/A vgnd vpwr scs8hd_or3_4
XFILLER_11_50 vpwr vgnd scs8hd_fill_2
XFILLER_14_172 vgnd vpwr scs8hd_decap_8
XFILLER_16_17 vgnd vpwr scs8hd_decap_4
XFILLER_16_28 vgnd vpwr scs8hd_fill_1
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA__084__D _084_/D vgnd vpwr scs8hd_diode_2
XFILLER_20_142 vpwr vgnd scs8hd_fill_2
XFILLER_20_186 vgnd vpwr scs8hd_decap_8
XFILLER_28_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_104_ _075_/A _104_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_19_231 vpwr vgnd scs8hd_fill_2
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XFILLER_27_16 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_201 vgnd vpwr scs8hd_decap_4
XFILLER_4_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
XFILLER_17_93 vpwr vgnd scs8hd_fill_2
XFILLER_3_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_1_119 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _132_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB _066_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_208 vgnd vpwr scs8hd_decap_6
XFILLER_13_204 vgnd vpwr scs8hd_decap_8
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XFILLER_8_230 vgnd vpwr scs8hd_decap_3
XFILLER_5_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_28 vpwr vgnd scs8hd_fill_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XFILLER_25_60 vgnd vpwr scs8hd_fill_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_107 vpwr vgnd scs8hd_fill_2
XFILLER_2_86 vgnd vpwr scs8hd_decap_4
XFILLER_21_29 vpwr vgnd scs8hd_fill_2
XANTENNA__098__C _098_/C vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_051_ _116_/A _051_/B _051_/Y vgnd vpwr scs8hd_nor2_4
X_120_ _120_/A _118_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_184 vgnd vpwr scs8hd_decap_3
XFILLER_23_151 vgnd vpwr scs8hd_decap_3
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_110 vpwr vgnd scs8hd_fill_2
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
X_103_ _120_/A _104_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_14_7 vgnd vpwr scs8hd_fill_1
XFILLER_19_210 vgnd vpwr scs8hd_decap_3
XFILLER_6_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_28 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_202 vpwr vgnd scs8hd_fill_2
XFILLER_17_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _040_/A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_42 vpwr vgnd scs8hd_fill_2
XFILLER_14_40 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_8
XANTENNA__101__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_105 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_65 vpwr vgnd scs8hd_fill_2
XFILLER_32_196 vgnd vpwr scs8hd_decap_12
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__D _084_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_050_ address[4] address[3] _069_/C _051_/B vgnd vpwr scs8hd_or3_4
XFILLER_2_3 vgnd vpwr scs8hd_decap_6
XFILLER_11_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_3_.latch data_in mem_top_ipin_1.LATCH_3_.latch/Q _055_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_200 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_7_148 vpwr vgnd scs8hd_fill_2
XFILLER_11_188 vgnd vpwr scs8hd_decap_3
X_102_ _119_/A _104_/B _102_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_62 vgnd vpwr scs8hd_decap_6
XFILLER_33_72 vpwr vgnd scs8hd_fill_2
XANTENNA__104__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_173 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_217 vgnd vpwr scs8hd_decap_12
XFILLER_0_176 vgnd vpwr scs8hd_decap_4
XFILLER_5_10 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_224 vgnd vpwr scs8hd_decap_8
XFILLER_30_84 vgnd vpwr scs8hd_decap_8
XFILLER_30_73 vpwr vgnd scs8hd_fill_2
XANTENNA__101__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_139 vpwr vgnd scs8hd_fill_2
XFILLER_2_205 vpwr vgnd scs8hd_fill_2
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_194 vpwr vgnd scs8hd_fill_2
XFILLER_26_150 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA__112__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_186 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_15_109 vgnd vpwr scs8hd_fill_1
XFILLER_11_31 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_4.LATCH_2_.latch data_in mem_top_ipin_4.LATCH_2_.latch/Q _080_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_131 vgnd vpwr scs8hd_decap_3
XANTENNA__107__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_8
XFILLER_20_178 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_6.LATCH_5_.latch data_in mem_top_ipin_6.LATCH_5_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_101_ _118_/A _104_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_138 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_223 vgnd vpwr scs8hd_decap_8
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_6
XFILLER_8_65 vgnd vpwr scs8hd_decap_4
XFILLER_4_108 vpwr vgnd scs8hd_fill_2
XFILLER_31_218 vpwr vgnd scs8hd_fill_2
XFILLER_31_207 vgnd vpwr scs8hd_decap_8
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XANTENNA__104__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_152 vpwr vgnd scs8hd_fill_2
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB _051_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_73 vpwr vgnd scs8hd_fill_2
XFILLER_28_51 vgnd vpwr scs8hd_decap_4
XANTENNA__115__A _122_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_88 vgnd vpwr scs8hd_decap_4
XFILLER_10_3 vgnd vpwr scs8hd_decap_4
XFILLER_14_53 vgnd vpwr scs8hd_decap_8
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_2_12 vgnd vpwr scs8hd_decap_12
XANTENNA__112__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_7.LATCH_1_.latch data_in mem_top_ipin_7.LATCH_1_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_162 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_132 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_54 vgnd vpwr scs8hd_decap_4
XFILLER_11_65 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_3
XANTENNA__107__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_20_146 vgnd vpwr scs8hd_decap_6
XFILLER_9_191 vpwr vgnd scs8hd_fill_2
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
X_100_ _117_/A _104_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_157 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_6
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_190 vgnd vpwr scs8hd_fill_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_86 vgnd vpwr scs8hd_decap_4
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_131 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_208 vgnd vpwr scs8hd_decap_4
XFILLER_22_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vpwr vgnd scs8hd_fill_2
XFILLER_0_101 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_34 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__041__A _041_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_218 vgnd vpwr scs8hd_decap_12
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_31 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vgnd vpwr scs8hd_decap_4
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_22 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__107__C _122_/C vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_125 vgnd vpwr scs8hd_decap_4
XFILLER_20_158 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_11_136 vgnd vpwr scs8hd_decap_8
XFILLER_22_54 vgnd vpwr scs8hd_decap_8
XFILLER_22_65 vgnd vpwr scs8hd_decap_3
XFILLER_22_76 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _126_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_195 vgnd vpwr scs8hd_decap_4
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
XANTENNA__044__A enable vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_8
XFILLER_17_54 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_2.LATCH_5_.latch data_in mem_top_ipin_2.LATCH_5_.latch/Q _063_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_198 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_90 vgnd vpwr scs8hd_fill_1
XANTENNA__039__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_231 vpwr vgnd scs8hd_fill_2
XFILLER_0_146 vpwr vgnd scs8hd_fill_2
XFILLER_28_86 vgnd vpwr scs8hd_decap_6
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_46 vpwr vgnd scs8hd_fill_2
XANTENNA__115__C _122_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__052__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_18_109 vpwr vgnd scs8hd_fill_2
XPHY_65 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_21 vgnd vpwr scs8hd_fill_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_98 vpwr vgnd scs8hd_fill_2
XFILLER_2_69 vpwr vgnd scs8hd_fill_2
XFILLER_2_36 vgnd vpwr scs8hd_fill_1
XFILLER_32_178 vgnd vpwr scs8hd_decap_6
XFILLER_32_112 vgnd vpwr scs8hd_decap_12
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_23_156 vpwr vgnd scs8hd_fill_2
XFILLER_23_189 vpwr vgnd scs8hd_fill_2
XANTENNA__047__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_89 vgnd vpwr scs8hd_decap_4
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
XFILLER_14_189 vpwr vgnd scs8hd_fill_2
XANTENNA__107__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_9_171 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_3.LATCH_1_.latch data_in mem_top_ipin_3.LATCH_1_.latch/Q _074_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_90 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _041_/A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_108 vgnd vpwr scs8hd_decap_4
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_174 vgnd vpwr scs8hd_decap_8
X_089_ _120_/A _088_/B _089_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_5.LATCH_4_.latch data_in mem_top_ipin_5.LATCH_4_.latch/Q _086_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__060__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_218 vgnd vpwr scs8hd_decap_12
XFILLER_17_33 vpwr vgnd scs8hd_fill_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_76 vpwr vgnd scs8hd_fill_2
XFILLER_33_43 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_188 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__055__A _051_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_43 vpwr vgnd scs8hd_fill_2
XFILLER_5_14 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_14_78 vgnd vpwr scs8hd_decap_3
XFILLER_30_66 vgnd vpwr scs8hd_decap_4
XFILLER_29_195 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
XFILLER_2_209 vgnd vpwr scs8hd_decap_4
XANTENNA__052__B _043_/Y vgnd vpwr scs8hd_diode_2
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_198 vgnd vpwr scs8hd_decap_12
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_44 vpwr vgnd scs8hd_fill_2
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_48 vpwr vgnd scs8hd_fill_2
XFILLER_2_26 vgnd vpwr scs8hd_decap_4
XFILLER_32_102 vgnd vpwr scs8hd_fill_1
XFILLER_17_187 vpwr vgnd scs8hd_fill_2
XFILLER_32_124 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__153__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_23_113 vgnd vpwr scs8hd_decap_3
XFILLER_23_102 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_46 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_102 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_6.LATCH_0_.latch data_in mem_top_ipin_6.LATCH_0_.latch/Q _097_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_138 vpwr vgnd scs8hd_fill_2
XFILLER_28_205 vgnd vpwr scs8hd_decap_8
XANTENNA__058__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_157_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_142 vpwr vgnd scs8hd_fill_2
XFILLER_8_69 vgnd vpwr scs8hd_fill_1
XFILLER_10_171 vgnd vpwr scs8hd_decap_6
XFILLER_10_193 vgnd vpwr scs8hd_fill_1
X_088_ _119_/A _088_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__060__B address[2] vgnd vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XFILLER_33_66 vgnd vpwr scs8hd_fill_1
XFILLER_33_11 vgnd vpwr scs8hd_decap_12
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
XFILLER_30_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB _057_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__055__B _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _117_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_55 vgnd vpwr scs8hd_fill_1
XFILLER_28_11 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_7 vgnd vpwr scs8hd_fill_1
XANTENNA__156__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__066__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_23 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_174 vgnd vpwr scs8hd_decap_3
XFILLER_29_163 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__052__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
XFILLER_26_144 vgnd vpwr scs8hd_decap_6
XFILLER_26_133 vgnd vpwr scs8hd_decap_8
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_56 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_32_136 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__063__B _062_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_58 vgnd vpwr scs8hd_fill_1
XFILLER_11_69 vgnd vpwr scs8hd_decap_3
XFILLER_2_9 vgnd vpwr scs8hd_fill_1
XFILLER_14_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__058__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_206 vpwr vgnd scs8hd_fill_2
X_156_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_087_ _118_/A _088_/B _087_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_154 vgnd vpwr scs8hd_decap_3
XFILLER_10_150 vgnd vpwr scs8hd_decap_3
XFILLER_12_90 vpwr vgnd scs8hd_fill_2
XANTENNA__060__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _122_/A vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_23 vgnd vpwr scs8hd_decap_12
XFILLER_17_68 vgnd vpwr scs8hd_fill_1
XFILLER_33_89 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _130_/HI _040_/Y mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
X_139_ _139_/HI _139_/LO vgnd vpwr scs8hd_conb_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_82 vpwr vgnd scs8hd_fill_2
XFILLER_21_201 vgnd vpwr scs8hd_decap_3
XFILLER_9_91 vgnd vpwr scs8hd_decap_4
XANTENNA__071__B _072_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_1.LATCH_4_.latch data_in mem_top_ipin_1.LATCH_4_.latch/Q _053_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_38 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _132_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__066__B _062_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_36 vpwr vgnd scs8hd_fill_2
XANTENNA__082__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_230 vgnd vpwr scs8hd_decap_3
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_81 vpwr vgnd scs8hd_fill_2
XFILLER_26_167 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3 vgnd vpwr scs8hd_decap_6
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_32_148 vgnd vpwr scs8hd_decap_4
XFILLER_17_145 vgnd vpwr scs8hd_decap_8
XFILLER_15_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _130_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_159 vpwr vgnd scs8hd_fill_2
XFILLER_9_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__058__C _058_/C vgnd vpwr scs8hd_diode_2
XANTENNA__074__B _072_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_0_7 vgnd vpwr scs8hd_fill_1
XANTENNA__090__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_38 vgnd vpwr scs8hd_fill_1
X_155_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_086_ _117_/A _088_/B _086_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_2.LATCH_0_.latch data_in mem_top_ipin_2.LATCH_0_.latch/Q _068_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__069__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_35 vgnd vpwr scs8hd_decap_8
XFILLER_24_210 vgnd vpwr scs8hd_decap_4
XANTENNA__085__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_58 vgnd vpwr scs8hd_decap_3
XFILLER_15_210 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_138_ _138_/HI _138_/LO vgnd vpwr scs8hd_conb_1
X_069_ _122_/A address[3] _069_/C _072_/B vgnd vpwr scs8hd_or3_4
Xmem_top_ipin_4.LATCH_3_.latch data_in mem_top_ipin_4.LATCH_3_.latch/Q _079_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _080_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_80 vgnd vpwr scs8hd_decap_4
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XFILLER_6_60 vpwr vgnd scs8hd_fill_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_179 vgnd vpwr scs8hd_decap_6
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _080_/B vgnd vpwr scs8hd_diode_2
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_212 vgnd vpwr scs8hd_decap_3
XFILLER_1_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _041_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_138 vpwr vgnd scs8hd_fill_2
XFILLER_16_190 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__088__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_127 vpwr vgnd scs8hd_fill_2
XFILLER_14_149 vgnd vpwr scs8hd_decap_4
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vpwr vgnd scs8hd_fill_2
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
XFILLER_28_219 vgnd vpwr scs8hd_decap_12
XANTENNA__090__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_219 vpwr vgnd scs8hd_fill_2
XFILLER_10_141 vgnd vpwr scs8hd_fill_1
X_154_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_123 vpwr vgnd scs8hd_fill_2
X_085_ _116_/A _088_/B _085_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_2_.latch data_in mem_top_ipin_7.LATCH_2_.latch/Q _102_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__069__C _069_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_37 vpwr vgnd scs8hd_fill_2
XANTENNA__085__B _088_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_91 vpwr vgnd scs8hd_fill_2
XFILLER_23_80 vgnd vpwr scs8hd_decap_4
X_137_ _137_/HI _137_/LO vgnd vpwr scs8hd_conb_1
X_068_ _075_/A _062_/X _068_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_170 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_6
XFILLER_28_47 vpwr vgnd scs8hd_fill_2
XFILLER_28_69 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_218 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _133_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_26 vgnd vpwr scs8hd_decap_4
XFILLER_29_199 vpwr vgnd scs8hd_fill_2
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_48 vgnd vpwr scs8hd_decap_6
XFILLER_25_15 vgnd vpwr scs8hd_decap_6
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _091_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_158 vpwr vgnd scs8hd_fill_2
XFILLER_31_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_183 vgnd vpwr scs8hd_decap_8
XFILLER_26_80 vgnd vpwr scs8hd_fill_1
XFILLER_9_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_73 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_231 vpwr vgnd scs8hd_fill_2
XFILLER_10_186 vgnd vpwr scs8hd_decap_4
X_153_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_146 vgnd vpwr scs8hd_decap_6
X_084_ address[4] address[3] _098_/C _084_/D _088_/B vgnd vpwr scs8hd_or4_4
XFILLER_12_82 vgnd vpwr scs8hd_decap_8
XFILLER_18_231 vpwr vgnd scs8hd_fill_2
XFILLER_17_16 vgnd vpwr scs8hd_decap_4
XFILLER_3_127 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
X_136_ _136_/HI _136_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_7.LATCH_3_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
X_067_ _120_/A _062_/X _067_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_9_72 vpwr vgnd scs8hd_fill_2
XFILLER_21_215 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_119_ _119_/A _118_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _125_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_49 vgnd vpwr scs8hd_decap_8
XFILLER_29_167 vgnd vpwr scs8hd_fill_1
XFILLER_29_134 vgnd vpwr scs8hd_decap_12
XFILLER_29_112 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_115 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_27 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_126 vpwr vgnd scs8hd_fill_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_15_82 vpwr vgnd scs8hd_fill_2
XFILLER_31_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_195 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_22_140 vpwr vgnd scs8hd_fill_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_188 vgnd vpwr scs8hd_fill_1
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_52 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_39 vgnd vpwr scs8hd_decap_6
XANTENNA__099__B _104_/B vgnd vpwr scs8hd_diode_2
X_152_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_083_ _083_/A address[5] _084_/D vgnd vpwr scs8hd_or2_4
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_61 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_202 vgnd vpwr scs8hd_decap_4
XFILLER_33_213 vgnd vpwr scs8hd_decap_12
XFILLER_33_49 vpwr vgnd scs8hd_fill_2
XFILLER_3_117 vgnd vpwr scs8hd_decap_3
XFILLER_30_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_135_ _135_/HI _135_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_71 vgnd vpwr scs8hd_decap_3
X_066_ _119_/A _062_/X _066_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_86 vgnd vpwr scs8hd_decap_4
XFILLER_0_97 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
XFILLER_9_95 vgnd vpwr scs8hd_fill_1
XFILLER_12_205 vgnd vpwr scs8hd_decap_8
XFILLER_12_227 vgnd vpwr scs8hd_decap_6
Xmem_top_ipin_3.LATCH_2_.latch data_in mem_top_ipin_3.LATCH_2_.latch/Q _073_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_231 vpwr vgnd scs8hd_fill_2
X_118_ _118_/A _118_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _134_/HI vgnd vpwr
+ scs8hd_diode_2
X_049_ enable _083_/A address[5] _069_/C vgnd vpwr scs8hd_nand3_4
XFILLER_14_29 vpwr vgnd scs8hd_fill_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_146 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_5.LATCH_5_.latch data_in mem_top_ipin_5.LATCH_5_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_81 vgnd vpwr scs8hd_fill_1
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vpwr vgnd scs8hd_fill_2
XFILLER_6_85 vgnd vpwr scs8hd_decap_6
XFILLER_26_105 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_25_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_163 vgnd vpwr scs8hd_fill_1
XFILLER_16_182 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _041_/Y mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_3_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_3
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_9_145 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_151_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_104 vpwr vgnd scs8hd_fill_2
XFILLER_6_159 vpwr vgnd scs8hd_fill_2
XFILLER_10_111 vgnd vpwr scs8hd_decap_6
XFILLER_10_133 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_082_ _075_/A _080_/B _082_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_225 vgnd vpwr scs8hd_decap_8
XFILLER_15_214 vgnd vpwr scs8hd_fill_1
X_065_ _118_/A _062_/X _065_/Y vgnd vpwr scs8hd_nor2_4
X_134_ _134_/HI _134_/LO vgnd vpwr scs8hd_conb_1
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_6.LATCH_1_.latch data_in mem_top_ipin_6.LATCH_1_.latch/Q _096_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _040_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _131_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_61 vgnd vpwr scs8hd_decap_8
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
X_117_ _117_/A _118_/B _117_/Y vgnd vpwr scs8hd_nor2_4
X_048_ address[1] _043_/Y _058_/C _116_/A vgnd vpwr scs8hd_or3_4
XFILLER_15_3 vgnd vpwr scs8hd_decap_3
XFILLER_14_19 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_20_73 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vgnd vpwr scs8hd_fill_1
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_29_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_20 vgnd vpwr scs8hd_decap_8
XFILLER_6_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _067_/Y vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_191 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_109 vpwr vgnd scs8hd_fill_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_72 vgnd vpwr scs8hd_decap_8
XFILLER_26_61 vgnd vpwr scs8hd_decap_3
XFILLER_9_113 vpwr vgnd scs8hd_fill_2
XFILLER_13_120 vpwr vgnd scs8hd_fill_2
XFILLER_13_153 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vgnd vpwr scs8hd_decap_4
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_43 vpwr vgnd scs8hd_fill_2
XFILLER_22_19 vgnd vpwr scs8hd_decap_12
XFILLER_27_223 vgnd vpwr scs8hd_decap_8
XFILLER_27_201 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_150_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_127 vgnd vpwr scs8hd_decap_4
XFILLER_10_145 vgnd vpwr scs8hd_decap_3
XFILLER_10_167 vpwr vgnd scs8hd_fill_2
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_12_74 vgnd vpwr scs8hd_decap_6
X_081_ _120_/A _080_/B _081_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_201 vpwr vgnd scs8hd_fill_2
XFILLER_5_171 vpwr vgnd scs8hd_fill_2
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_133_ _133_/HI _133_/LO vgnd vpwr scs8hd_conb_1
X_064_ _117_/A _062_/X _064_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__110__A _117_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_18_73 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _116_/A _118_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _098_/C vgnd vpwr scs8hd_diode_2
X_047_ address[3] _122_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _135_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_19 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_3_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_29_159 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_29_50 vgnd vpwr scs8hd_decap_3
XFILLER_26_118 vgnd vpwr scs8hd_decap_4
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_217 vgnd vpwr scs8hd_decap_12
XFILLER_9_9 vgnd vpwr scs8hd_fill_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_25_140 vgnd vpwr scs8hd_fill_1
XFILLER_31_84 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_3
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_1.LATCH_5_.latch data_in mem_top_ipin_1.LATCH_5_.latch/Q _051_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__102__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XFILLER_16_162 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_3
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_9_158 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vgnd vpwr scs8hd_decap_4
XANTENNA__113__A _120_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_99 vgnd vpwr scs8hd_decap_3
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_080_ _119_/A _080_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
X_063_ _116_/A _062_/X _063_/Y vgnd vpwr scs8hd_nor2_4
X_132_ _132_/HI _132_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_186 vpwr vgnd scs8hd_fill_2
XFILLER_2_131 vgnd vpwr scs8hd_decap_3
XFILLER_2_120 vgnd vpwr scs8hd_decap_4
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_21 vgnd vpwr scs8hd_decap_4
XFILLER_9_76 vpwr vgnd scs8hd_fill_2
XFILLER_21_219 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_96 vgnd vpwr scs8hd_decap_6
XANTENNA__105__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_7_223 vgnd vpwr scs8hd_decap_8
X_046_ address[4] _122_/A vgnd vpwr scs8hd_inv_8
X_115_ _122_/A address[3] _122_/C _118_/B vgnd vpwr scs8hd_or3_4
XANTENNA__121__A _075_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_116 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_2.LATCH_1_.latch data_in mem_top_ipin_2.LATCH_1_.latch/Q _067_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_4.LATCH_4_.latch data_in mem_top_ipin_4.LATCH_4_.latch/Q _078_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XFILLER_15_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_111 vpwr vgnd scs8hd_fill_2
XFILLER_16_174 vgnd vpwr scs8hd_decap_8
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

