* NGSPICE file created from cbx_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

.subckt cbx_1__1_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] prog_clk
+ top_grid_pin_16_ top_grid_pin_17_ top_grid_pin_18_ top_grid_pin_19_ top_grid_pin_20_
+ top_grid_pin_21_ top_grid_pin_22_ top_grid_pin_23_ top_grid_pin_24_ top_grid_pin_25_
+ top_grid_pin_26_ top_grid_pin_27_ top_grid_pin_28_ top_grid_pin_29_ top_grid_pin_30_
+ top_grid_pin_31_ VPWR VGND
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_12.mux_l2_in_3_ _23_/HI chanx_right_in[16] mux_bottom_ipin_12.mux_l2_in_2_/S
+ mux_bottom_ipin_12.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_7.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_bottom_ipin_7.mux_l2_in_1_/S
+ mux_bottom_ipin_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_66_ chanx_left_in[5] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S mux_bottom_ipin_4.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_12.mux_l3_in_1_/S
+ mux_bottom_ipin_12.mux_l4_in_0_/S mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_49_ chanx_right_in[2] chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_15.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_2.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_12.mux_l4_in_0_ mux_bottom_ipin_12.mux_l3_in_1_/X mux_bottom_ipin_12.mux_l3_in_0_/X
+ mux_bottom_ipin_12.mux_l4_in_0_/S mux_bottom_ipin_12.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_2.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_2.mux_l1_in_0_/X
+ mux_bottom_ipin_2.mux_l2_in_3_/S mux_bottom_ipin_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S mux_bottom_ipin_13.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S mux_bottom_ipin_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_12.mux_l3_in_1_ mux_bottom_ipin_12.mux_l2_in_3_/X mux_bottom_ipin_12.mux_l2_in_2_/X
+ mux_bottom_ipin_12.mux_l3_in_1_/S mux_bottom_ipin_12.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S mux_bottom_ipin_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1 mux_bottom_ipin_15.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0 _29_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S mux_bottom_ipin_2.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_12.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[12] mux_bottom_ipin_12.mux_l2_in_2_/S
+ mux_bottom_ipin_12.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0 mux_bottom_ipin_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_15.mux_l3_in_1_/S
+ ccff_tail mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_bottom_ipin_7.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_7.mux_l1_in_0_/X
+ mux_bottom_ipin_7.mux_l2_in_1_/S mux_bottom_ipin_7.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S mux_bottom_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_5.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_5.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_65_ chanx_left_in[6] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S mux_bottom_ipin_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S mux_bottom_ipin_1.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_7.mux_l4_in_0_/X top_grid_pin_23_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_12.mux_l2_in_2_/S
+ mux_bottom_ipin_12.mux_l3_in_1_/S mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_2.mux_l3_in_1_/S mux_bottom_ipin_2.mux_l4_in_0_/S
+ mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_48_ chanx_right_in[3] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S mux_bottom_ipin_7.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0 mux_bottom_ipin_10.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_12.mux_l3_in_0_ mux_bottom_ipin_12.mux_l2_in_1_/X mux_bottom_ipin_12.mux_l2_in_0_/X
+ mux_bottom_ipin_12.mux_l3_in_1_/S mux_bottom_ipin_12.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_2.mux_l1_in_0_/S
+ mux_bottom_ipin_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_8.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_8.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1 mux_bottom_ipin_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_12.mux_l2_in_1_ chanx_left_in[12] mux_bottom_ipin_12.mux_l1_in_2_/X
+ mux_bottom_ipin_12.mux_l2_in_2_/S mux_bottom_ipin_12.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_15.mux_l2_in_2_/S
+ mux_bottom_ipin_15.mux_l3_in_1_/S mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_5.mux_l3_in_1_/S mux_bottom_ipin_5.mux_l4_in_0_/S
+ mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_12.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_64_ chanx_left_in[7] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S mux_bottom_ipin_15.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_12.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_bottom_ipin_12.mux_l1_in_2_/S
+ mux_bottom_ipin_12.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_7.mux_l1_in_0_/S
+ mux_bottom_ipin_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_12.mux_l1_in_2_/S
+ mux_bottom_ipin_12.mux_l2_in_2_/S mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_2.mux_l2_in_3_/S mux_bottom_ipin_2.mux_l3_in_1_/S
+ mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_47_ chanx_right_in[4] chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S mux_bottom_ipin_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S mux_bottom_ipin_14.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1 mux_bottom_ipin_10.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0 mux_bottom_ipin_1.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_8.mux_l3_in_1_/S mux_bottom_ipin_8.mux_l4_in_0_/S
+ mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S mux_bottom_ipin_13.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S mux_bottom_ipin_5.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_12.mux_l2_in_0_ mux_bottom_ipin_12.mux_l1_in_1_/X mux_bottom_ipin_12.mux_l1_in_0_/X
+ mux_bottom_ipin_12.mux_l2_in_2_/S mux_bottom_ipin_12.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_15.mux_l1_in_0_/S
+ mux_bottom_ipin_15.mux_l2_in_2_/S mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_5.mux_l2_in_3_/S mux_bottom_ipin_5.mux_l3_in_1_/S
+ mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_63_ chanx_left_in[8] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S mux_bottom_ipin_14.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S mux_bottom_ipin_12.mux_l4_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S mux_bottom_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_12.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_12.mux_l1_in_2_/S
+ mux_bottom_ipin_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_11.mux_l4_in_0_/S
+ mux_bottom_ipin_12.mux_l1_in_2_/S mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_2.mux_l1_in_0_/S mux_bottom_ipin_2.mux_l2_in_3_/S
+ mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_46_ chanx_right_in[5] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1 mux_bottom_ipin_1.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29_ _29_/HI _29_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S mux_bottom_ipin_3.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0 mux_bottom_ipin_8.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_0.mux_l4_in_0_/X top_grid_pin_16_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_bottom_ipin_12.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_12.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S mux_bottom_ipin_9.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1 mux_bottom_ipin_1.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_8.mux_l2_in_2_/S mux_bottom_ipin_8.mux_l3_in_1_/S
+ mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0 mux_bottom_ipin_8.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_14.mux_l4_in_0_/S
+ mux_bottom_ipin_15.mux_l1_in_0_/S mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_5.mux_l1_in_1_/S mux_bottom_ipin_5.mux_l2_in_3_/S
+ mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_62_ chanx_left_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0 mux_bottom_ipin_12.mux_l2_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_12.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_12.mux_l1_in_2_/S
+ mux_bottom_ipin_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_1.mux_l4_in_0_/S mux_bottom_ipin_2.mux_l1_in_0_/S
+ mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_45_ chanx_right_in[6] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_15.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_15.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_13.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S mux_bottom_ipin_11.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0 mux_bottom_ipin_12.mux_l3_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28_ _28_/HI _28_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1 mux_bottom_ipin_8.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_8.mux_l1_in_2_/S mux_bottom_ipin_8.mux_l2_in_2_/S
+ mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1 mux_bottom_ipin_14.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_3.mux_l2_in_3_ _28_/HI chanx_right_in[15] mux_bottom_ipin_3.mux_l2_in_0_/S
+ mux_bottom_ipin_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S mux_bottom_ipin_10.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0 mux_bottom_ipin_5.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1 mux_bottom_ipin_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_9.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_14.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_4.mux_l4_in_0_/S mux_bottom_ipin_5.mux_l1_in_1_/S
+ mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S mux_bottom_ipin_1.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_61_ chanx_left_in[10] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_3.mux_l4_in_0_ mux_bottom_ipin_3.mux_l3_in_1_/X mux_bottom_ipin_3.mux_l3_in_0_/X
+ mux_bottom_ipin_3.mux_l4_in_0_/S mux_bottom_ipin_3.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S mux_bottom_ipin_15.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1 mux_bottom_ipin_12.mux_l2_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_44_ chanx_right_in[7] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_8.mux_l2_in_3_ _17_/HI chanx_right_in[18] mux_bottom_ipin_8.mux_l2_in_2_/S
+ mux_bottom_ipin_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0 mux_bottom_ipin_3.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S mux_bottom_ipin_10.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S mux_bottom_ipin_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_3.mux_l3_in_1_ mux_bottom_ipin_3.mux_l2_in_3_/X mux_bottom_ipin_3.mux_l2_in_2_/X
+ mux_bottom_ipin_3.mux_l3_in_0_/S mux_bottom_ipin_3.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1 mux_bottom_ipin_12.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ _27_/HI _27_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S mux_bottom_ipin_14.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__34__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0 mux_bottom_ipin_3.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_7.mux_l4_in_0_/S mux_bottom_ipin_8.mux_l1_in_2_/S
+ mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_ipin_3.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_bottom_ipin_3.mux_l2_in_0_/S
+ mux_bottom_ipin_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_8.mux_l4_in_0_ mux_bottom_ipin_8.mux_l3_in_1_/X mux_bottom_ipin_8.mux_l3_in_0_/X
+ mux_bottom_ipin_8.mux_l4_in_0_/S mux_bottom_ipin_8.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1 mux_bottom_ipin_5.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S mux_bottom_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S mux_bottom_ipin_9.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_8.mux_l3_in_1_ mux_bottom_ipin_8.mux_l2_in_3_/X mux_bottom_ipin_8.mux_l2_in_2_/X
+ mux_bottom_ipin_8.mux_l3_in_1_/S mux_bottom_ipin_8.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__42__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_10.mux_l4_in_0_/X top_grid_pin_26_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
X_60_ chanx_left_in[11] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__37__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_43_ chanx_right_in[8] chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_8.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_bottom_ipin_8.mux_l2_in_2_/S
+ mux_bottom_ipin_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S mux_bottom_ipin_8.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1 mux_bottom_ipin_3.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_3.mux_l3_in_0_ mux_bottom_ipin_3.mux_l2_in_1_/X mux_bottom_ipin_3.mux_l2_in_0_/X
+ mux_bottom_ipin_3.mux_l3_in_0_/S mux_bottom_ipin_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_26_ _26_/HI _26_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0 _25_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__50__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1 mux_bottom_ipin_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0 mux_bottom_ipin_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_3.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_bottom_ipin_3.mux_l2_in_0_/S
+ mux_bottom_ipin_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__45__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_8.mux_l3_in_0_ mux_bottom_ipin_8.mux_l2_in_1_/X mux_bottom_ipin_8.mux_l2_in_0_/X
+ mux_bottom_ipin_8.mux_l3_in_1_/S mux_bottom_ipin_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S mux_bottom_ipin_12.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_13.mux_l2_in_3_ _24_/HI chanx_right_in[17] mux_bottom_ipin_13.mux_l2_in_3_/S
+ mux_bottom_ipin_13.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__53__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ chanx_right_in[9] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_8.mux_l2_in_1_ chanx_left_in[12] mux_bottom_ipin_8.mux_l1_in_2_/X
+ mux_bottom_ipin_8.mux_l2_in_2_/S mux_bottom_ipin_8.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S mux_bottom_ipin_11.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__48__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25_ _25_/HI _25_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S mux_bottom_ipin_7.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1 mux_bottom_ipin_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_8.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_bottom_ipin_8.mux_l1_in_2_/S
+ mux_bottom_ipin_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_ipin_13.mux_l4_in_0_ mux_bottom_ipin_13.mux_l3_in_1_/X mux_bottom_ipin_13.mux_l3_in_0_/X
+ mux_bottom_ipin_13.mux_l4_in_0_/S mux_bottom_ipin_13.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_3.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_3.mux_l1_in_0_/X
+ mux_bottom_ipin_3.mux_l2_in_0_/S mux_bottom_ipin_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S mux_bottom_ipin_10.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_3.mux_l4_in_0_/X top_grid_pin_19_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__61__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0 mux_bottom_ipin_7.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S mux_bottom_ipin_6.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__56__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_13.mux_l3_in_1_ mux_bottom_ipin_13.mux_l2_in_3_/X mux_bottom_ipin_13.mux_l2_in_2_/X
+ mux_bottom_ipin_13.mux_l3_in_1_/S mux_bottom_ipin_13.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S mux_bottom_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S mux_bottom_ipin_5.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_13.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[13] mux_bottom_ipin_13.mux_l2_in_3_/S
+ mux_bottom_ipin_13.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_41_ chanx_right_in[10] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_8.mux_l2_in_0_ mux_bottom_ipin_8.mux_l1_in_1_/X mux_bottom_ipin_8.mux_l1_in_0_/X
+ mux_bottom_ipin_8.mux_l2_in_2_/S mux_bottom_ipin_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0 mux_bottom_ipin_11.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__64__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24_ _24_/HI _24_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S mux_bottom_ipin_6.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S mux_bottom_ipin_4.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__59__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_8.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_8.mux_l1_in_2_/S
+ mux_bottom_ipin_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1 mux_bottom_ipin_7.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_13.mux_l3_in_0_ mux_bottom_ipin_13.mux_l2_in_1_/X mux_bottom_ipin_13.mux_l2_in_0_/X
+ mux_bottom_ipin_13.mux_l3_in_1_/S mux_bottom_ipin_13.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_3.mux_l1_in_0_/S
+ mux_bottom_ipin_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_12.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__67__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_13.mux_l2_in_1_ chanx_left_in[13] mux_bottom_ipin_13.mux_l1_in_2_/X
+ mux_bottom_ipin_13.mux_l2_in_3_/S mux_bottom_ipin_13.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_40_ chanx_right_in[11] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1 mux_bottom_ipin_11.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0 _19_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23_ _23_/HI _23_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0 mux_bottom_ipin_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_13.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_bottom_ipin_13.mux_l1_in_1_/S
+ mux_bottom_ipin_13.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_8.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_ipin_8.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_8.mux_l1_in_2_/S
+ mux_bottom_ipin_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_13.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S mux_bottom_ipin_13.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S mux_bottom_ipin_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S mux_bottom_ipin_12.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S mux_bottom_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S mux_bottom_ipin_8.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_13.mux_l4_in_0_/X top_grid_pin_29_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_bottom_ipin_13.mux_l2_in_0_ mux_bottom_ipin_13.mux_l1_in_1_/X mux_bottom_ipin_13.mux_l1_in_0_/X
+ mux_bottom_ipin_13.mux_l2_in_3_/S mux_bottom_ipin_13.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0 mux_bottom_ipin_9.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S mux_bottom_ipin_1.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22_ _22_/HI _22_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1 mux_bottom_ipin_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S mux_bottom_ipin_7.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_13.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_13.mux_l1_in_1_/S
+ mux_bottom_ipin_13.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0 mux_bottom_ipin_9.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S mux_bottom_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S mux_bottom_ipin_0.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S mux_bottom_ipin_6.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0 mux_bottom_ipin_13.mux_l2_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0 mux_bottom_ipin_13.mux_l3_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_5.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1 mux_bottom_ipin_9.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21_ _21_/HI _21_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_ipin_13.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_13.mux_l1_in_1_/S
+ mux_bottom_ipin_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1 mux_bottom_ipin_15.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1 mux_bottom_ipin_9.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S mux_bottom_ipin_14.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_6.mux_l4_in_0_/X top_grid_pin_22_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1 mux_bottom_ipin_13.mux_l2_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_4.mux_l2_in_3_ _29_/HI chanx_right_in[14] mux_bottom_ipin_4.mux_l2_in_0_/S
+ mux_bottom_ipin_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_11.mux_l3_in_0_/S
+ mux_bottom_ipin_11.mux_l4_in_0_/S mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S mux_bottom_ipin_13.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_1.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0 mux_bottom_ipin_4.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1 mux_bottom_ipin_13.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S mux_bottom_ipin_12.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S mux_bottom_ipin_4.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_ipin_4.mux_l4_in_0_ mux_bottom_ipin_4.mux_l3_in_1_/X mux_bottom_ipin_4.mux_l3_in_0_/X
+ mux_bottom_ipin_4.mux_l4_in_0_/S mux_bottom_ipin_4.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0 mux_bottom_ipin_4.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20_ _20_/HI _20_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_9.mux_l2_in_3_ _18_/HI chanx_right_in[19] mux_bottom_ipin_9.mux_l2_in_2_/S
+ mux_bottom_ipin_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1 mux_bottom_ipin_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S mux_bottom_ipin_13.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_4.mux_l3_in_1_ mux_bottom_ipin_4.mux_l2_in_3_/X mux_bottom_ipin_4.mux_l2_in_2_/X
+ mux_bottom_ipin_4.mux_l3_in_0_/S mux_bottom_ipin_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_14.mux_l3_in_0_/S
+ mux_bottom_ipin_14.mux_l4_in_0_/S mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S mux_bottom_ipin_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S mux_bottom_ipin_11.mux_l4_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_4.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S mux_bottom_ipin_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_bottom_ipin_4.mux_l2_in_0_/S
+ mux_bottom_ipin_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_11.mux_l2_in_3_/S
+ mux_bottom_ipin_11.mux_l3_in_0_/S mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_1.mux_l3_in_1_/S mux_bottom_ipin_1.mux_l4_in_0_/S
+ mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_bottom_ipin_9.mux_l4_in_0_ mux_bottom_ipin_9.mux_l3_in_1_/X mux_bottom_ipin_9.mux_l3_in_0_/X
+ mux_bottom_ipin_9.mux_l4_in_0_/S mux_bottom_ipin_9.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S mux_bottom_ipin_2.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1 mux_bottom_ipin_4.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S mux_bottom_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1 mux_bottom_ipin_10.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_9.mux_l3_in_1_ mux_bottom_ipin_9.mux_l2_in_3_/X mux_bottom_ipin_9.mux_l2_in_2_/X
+ mux_bottom_ipin_9.mux_l3_in_1_/S mux_bottom_ipin_9.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0 _26_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0 mux_bottom_ipin_1.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1 mux_bottom_ipin_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_7.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_7.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_9.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_bottom_ipin_9.mux_l2_in_2_/S
+ mux_bottom_ipin_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_11.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_4.mux_l3_in_0_ mux_bottom_ipin_4.mux_l2_in_1_/X mux_bottom_ipin_4.mux_l2_in_0_/X
+ mux_bottom_ipin_4.mux_l3_in_0_/S mux_bottom_ipin_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_14.mux_l2_in_1_/S
+ mux_bottom_ipin_14.mux_l3_in_0_/S mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_4.mux_l3_in_0_/S mux_bottom_ipin_4.mux_l4_in_0_/S
+ mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S mux_bottom_ipin_10.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_bottom_ipin_4.mux_l1_in_2_/X
+ mux_bottom_ipin_4.mux_l2_in_0_/S mux_bottom_ipin_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_11.mux_l1_in_0_/S
+ mux_bottom_ipin_11.mux_l2_in_3_/S mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_1.mux_l2_in_0_/S mux_bottom_ipin_1.mux_l3_in_1_/S
+ mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_4.mux_l1_in_0_/S
+ mux_bottom_ipin_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_12.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_9.mux_l3_in_0_ mux_bottom_ipin_9.mux_l2_in_1_/X mux_bottom_ipin_9.mux_l2_in_0_/X
+ mux_bottom_ipin_9.mux_l3_in_1_/S mux_bottom_ipin_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1 mux_bottom_ipin_1.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_7.mux_l3_in_0_/S mux_bottom_ipin_7.mux_l4_in_0_/S
+ mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0 _31_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_14.mux_l2_in_3_ _25_/HI chanx_right_in[18] mux_bottom_ipin_14.mux_l2_in_1_/S
+ mux_bottom_ipin_14.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S mux_bottom_ipin_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0 mux_bottom_ipin_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_9.mux_l2_in_1_ chanx_left_in[13] mux_bottom_ipin_9.mux_l1_in_2_/X
+ mux_bottom_ipin_9.mux_l2_in_2_/S mux_bottom_ipin_9.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S mux_bottom_ipin_14.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_14.mux_l1_in_0_/S
+ mux_bottom_ipin_14.mux_l2_in_1_/S mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_4.mux_l2_in_0_/S mux_bottom_ipin_4.mux_l3_in_0_/S
+ mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_ipin_9.mux_l1_in_2_ chanx_right_in[9] chanx_left_in[9] mux_bottom_ipin_9.mux_l1_in_0_/S
+ mux_bottom_ipin_9.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_14.mux_l4_in_0_ mux_bottom_ipin_14.mux_l3_in_1_/X mux_bottom_ipin_14.mux_l3_in_0_/X
+ mux_bottom_ipin_14.mux_l4_in_0_/S mux_bottom_ipin_14.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_4.mux_l2_in_0_ mux_bottom_ipin_4.mux_l1_in_1_/X mux_bottom_ipin_4.mux_l1_in_0_/X
+ mux_bottom_ipin_4.mux_l2_in_0_/S mux_bottom_ipin_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_10.mux_l4_in_0_/S
+ mux_bottom_ipin_11.mux_l1_in_0_/S mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_1.mux_l1_in_2_/S mux_bottom_ipin_1.mux_l2_in_0_/S
+ mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S mux_bottom_ipin_13.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S mux_bottom_ipin_5.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0 _21_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S mux_bottom_ipin_9.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0 mux_bottom_ipin_12.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_4.mux_l1_in_0_/S
+ mux_bottom_ipin_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_14.mux_l3_in_1_ mux_bottom_ipin_14.mux_l2_in_3_/X mux_bottom_ipin_14.mux_l2_in_2_/X
+ mux_bottom_ipin_14.mux_l3_in_0_/S mux_bottom_ipin_14.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1 mux_bottom_ipin_8.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_11.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S mux_bottom_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_7.mux_l2_in_1_/S mux_bottom_ipin_7.mux_l3_in_0_/S
+ mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S mux_bottom_ipin_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_14.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_bottom_ipin_14.mux_l2_in_1_/S
+ mux_bottom_ipin_14.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1 mux_bottom_ipin_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_9.mux_l2_in_0_ mux_bottom_ipin_9.mux_l1_in_1_/X mux_bottom_ipin_9.mux_l1_in_0_/X
+ mux_bottom_ipin_9.mux_l2_in_2_/S mux_bottom_ipin_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_13.mux_l4_in_0_/S
+ mux_bottom_ipin_14.mux_l1_in_0_/S mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_4.mux_l1_in_0_/S mux_bottom_ipin_4.mux_l2_in_0_/S
+ mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S mux_bottom_ipin_9.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S mux_bottom_ipin_7.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_9.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_9.mux_l1_in_0_/S
+ mux_bottom_ipin_9.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1 mux_bottom_ipin_12.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_9.mux_l4_in_0_/X top_grid_pin_25_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_0.mux_l4_in_0_/S mux_bottom_ipin_1.mux_l1_in_2_/S
+ mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_14.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_14.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1 mux_bottom_ipin_12.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_14.mux_l3_in_0_ mux_bottom_ipin_14.mux_l2_in_1_/X mux_bottom_ipin_14.mux_l2_in_0_/X
+ mux_bottom_ipin_14.mux_l3_in_0_/S mux_bottom_ipin_14.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0 _20_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_4.mux_l1_in_0_/S
+ mux_bottom_ipin_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0 mux_bottom_ipin_3.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_7.mux_l1_in_0_/S mux_bottom_ipin_7.mux_l2_in_1_/S
+ mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_14.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_bottom_ipin_14.mux_l2_in_1_/S
+ mux_bottom_ipin_14.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_59_ chanx_left_in[12] chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_3.mux_l4_in_0_/S mux_bottom_ipin_4.mux_l1_in_0_/S
+ mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_9.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_9.mux_l1_in_0_/S
+ mux_bottom_ipin_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S mux_bottom_ipin_10.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S mux_bottom_ipin_6.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__32__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S mux_bottom_ipin_1.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1 mux_bottom_ipin_3.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S mux_bottom_ipin_15.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S mux_bottom_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_6.mux_l4_in_0_/S mux_bottom_ipin_7.mux_l1_in_0_/S
+ mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_bottom_ipin_14.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_14.mux_l1_in_0_/X
+ mux_bottom_ipin_14.mux_l2_in_1_/S mux_bottom_ipin_14.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__40__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S mux_bottom_ipin_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_58_ chanx_left_in[13] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S mux_bottom_ipin_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__35__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0 mux_bottom_ipin_14.mux_l2_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S mux_bottom_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S mux_bottom_ipin_3.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0 mux_bottom_ipin_14.mux_l3_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S mux_bottom_ipin_9.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__43__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_10.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_2.mux_l4_in_0_/X top_grid_pin_18_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__38__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_57_ chanx_left_in[14] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_0.mux_l2_in_3_ _19_/HI chanx_right_in[16] mux_bottom_ipin_0.mux_l2_in_0_/S
+ mux_bottom_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__51__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_14.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_14.mux_l1_in_0_/S
+ mux_bottom_ipin_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1 mux_bottom_ipin_14.mux_l2_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__46__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_11.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0 mux_bottom_ipin_5.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l4_in_0_ mux_bottom_ipin_0.mux_l3_in_1_/X mux_bottom_ipin_0.mux_l3_in_0_/X
+ mux_bottom_ipin_0.mux_l4_in_0_/S mux_bottom_ipin_0.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1 mux_bottom_ipin_14.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S mux_bottom_ipin_12.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0 mux_bottom_ipin_5.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S mux_bottom_ipin_2.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_5.mux_l2_in_3_ _30_/HI chanx_right_in[15] mux_bottom_ipin_5.mux_l2_in_3_/S
+ mux_bottom_ipin_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l3_in_1_ mux_bottom_ipin_0.mux_l2_in_3_/X mux_bottom_ipin_0.mux_l2_in_2_/X
+ mux_bottom_ipin_0.mux_l3_in_0_/S mux_bottom_ipin_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__54__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1 mux_bottom_ipin_7.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S mux_bottom_ipin_11.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__49__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S mux_bottom_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_bottom_ipin_0.mux_l2_in_0_/S
+ mux_bottom_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_56_ chanx_left_in[15] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S mux_bottom_ipin_15.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_5.mux_l4_in_0_ mux_bottom_ipin_5.mux_l3_in_1_/X mux_bottom_ipin_5.mux_l3_in_0_/X
+ mux_bottom_ipin_5.mux_l4_in_0_/S mux_bottom_ipin_5.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_39_ chanx_right_in[12] chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__62__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S mux_bottom_ipin_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1 mux_bottom_ipin_5.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_5.mux_l3_in_1_ mux_bottom_ipin_5.mux_l2_in_3_/X mux_bottom_ipin_5.mux_l2_in_2_/X
+ mux_bottom_ipin_5.mux_l3_in_1_/S mux_bottom_ipin_5.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S mux_bottom_ipin_14.mux_l4_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S mux_bottom_ipin_6.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__57__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1 mux_bottom_ipin_11.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1 mux_bottom_ipin_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S mux_bottom_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_ipin_5.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_bottom_ipin_5.mux_l2_in_3_/S
+ mux_bottom_ipin_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_ipin_0.mux_l3_in_0_ mux_bottom_ipin_0.mux_l2_in_1_/X mux_bottom_ipin_0.mux_l2_in_0_/X
+ mux_bottom_ipin_0.mux_l3_in_0_/S mux_bottom_ipin_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S mux_bottom_ipin_5.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__70__A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__65__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_bottom_ipin_0.mux_l1_in_2_/X
+ mux_bottom_ipin_0.mux_l2_in_0_/S mux_bottom_ipin_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_55_ chanx_left_in[16] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0 mux_bottom_ipin_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_12.mux_l4_in_0_/X top_grid_pin_28_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_38_ chanx_right_in[13] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_0.mux_l1_in_1_/S
+ mux_bottom_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0 mux_bottom_ipin_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_5.mux_l3_in_0_ mux_bottom_ipin_5.mux_l2_in_1_/X mux_bottom_ipin_5.mux_l2_in_0_/X
+ mux_bottom_ipin_5.mux_l3_in_1_/S mux_bottom_ipin_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_7.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_13.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_10.mux_l2_in_3_ _21_/HI chanx_right_in[14] mux_bottom_ipin_10.mux_l2_in_1_/S
+ mux_bottom_ipin_10.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S mux_bottom_ipin_13.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1 mux_bottom_ipin_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__68__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_5.mux_l2_in_1_ chanx_left_in[9] mux_bottom_ipin_5.mux_l1_in_2_/X
+ mux_bottom_ipin_5.mux_l2_in_3_/S mux_bottom_ipin_5.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0 _16_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0 mux_bottom_ipin_9.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_71_ chanx_left_in[0] chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_5.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_bottom_ipin_5.mux_l1_in_1_/S
+ mux_bottom_ipin_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S mux_bottom_ipin_12.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_10.mux_l4_in_0_ mux_bottom_ipin_10.mux_l3_in_1_/X mux_bottom_ipin_10.mux_l3_in_0_/X
+ mux_bottom_ipin_10.mux_l4_in_0_/S mux_bottom_ipin_10.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_54_ chanx_left_in[17] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_0.mux_l2_in_0_ mux_bottom_ipin_0.mux_l1_in_1_/X mux_bottom_ipin_0.mux_l1_in_0_/X
+ mux_bottom_ipin_0.mux_l2_in_0_/S mux_bottom_ipin_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1 mux_bottom_ipin_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ chanx_right_in[14] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_15.mux_l2_in_3_ _26_/HI chanx_right_in[19] mux_bottom_ipin_15.mux_l2_in_2_/S
+ mux_bottom_ipin_15.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S mux_bottom_ipin_11.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_10.mux_l3_in_1_ mux_bottom_ipin_10.mux_l2_in_3_/X mux_bottom_ipin_10.mux_l2_in_2_/X
+ mux_bottom_ipin_10.mux_l3_in_1_/S mux_bottom_ipin_10.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_0.mux_l1_in_1_/S
+ mux_bottom_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0 _22_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1 mux_bottom_ipin_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0 mux_bottom_ipin_13.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1 mux_bottom_ipin_9.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_10.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_bottom_ipin_10.mux_l2_in_1_/S
+ mux_bottom_ipin_10.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S mux_bottom_ipin_12.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S mux_bottom_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S mux_bottom_ipin_10.mux_l4_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_15.mux_l4_in_0_ mux_bottom_ipin_15.mux_l3_in_1_/X mux_bottom_ipin_15.mux_l3_in_0_/X
+ ccff_tail mux_bottom_ipin_15.mux_l4_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_5.mux_l2_in_0_ mux_bottom_ipin_5.mux_l1_in_1_/X mux_bottom_ipin_5.mux_l1_in_0_/X
+ mux_bottom_ipin_5.mux_l2_in_3_/S mux_bottom_ipin_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S mux_bottom_ipin_8.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1 mux_bottom_ipin_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_5.mux_l4_in_0_/X top_grid_pin_21_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_70_ chanx_left_in[1] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_15.mux_l3_in_1_ mux_bottom_ipin_15.mux_l2_in_3_/X mux_bottom_ipin_15.mux_l2_in_2_/X
+ mux_bottom_ipin_15.mux_l3_in_1_/S mux_bottom_ipin_15.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_5.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_5.mux_l1_in_1_/S
+ mux_bottom_ipin_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S mux_bottom_ipin_1.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_53_ chanx_left_in[18] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S mux_bottom_ipin_7.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1 mux_bottom_ipin_13.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36_ chanx_right_in[15] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_15.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_bottom_ipin_15.mux_l2_in_2_/S
+ mux_bottom_ipin_15.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_10.mux_l3_in_0_ mux_bottom_ipin_10.mux_l2_in_1_/X mux_bottom_ipin_10.mux_l2_in_0_/X
+ mux_bottom_ipin_10.mux_l3_in_1_/S mux_bottom_ipin_10.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_0.mux_l1_in_1_/S
+ mux_bottom_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1 mux_bottom_ipin_13.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19_ _19_/HI _19_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0 _27_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0 mux_bottom_ipin_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_10.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_bottom_ipin_10.mux_l2_in_1_/S
+ mux_bottom_ipin_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_15.mux_l3_in_0_ mux_bottom_ipin_15.mux_l2_in_1_/X mux_bottom_ipin_15.mux_l2_in_0_/X
+ mux_bottom_ipin_15.mux_l3_in_1_/S mux_bottom_ipin_15.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_5.mux_l1_in_1_/S
+ mux_bottom_ipin_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_10.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_52_ chanx_left_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_10.mux_l3_in_1_/S
+ mux_bottom_ipin_10.mux_l4_in_0_/S mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35_ chanx_right_in[16] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_15.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_bottom_ipin_15.mux_l2_in_2_/S
+ mux_bottom_ipin_15.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1 mux_bottom_ipin_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18_ _18_/HI _18_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_15.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1 mux_bottom_ipin_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_ipin_10.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_10.mux_l1_in_0_/X
+ mux_bottom_ipin_10.mux_l2_in_1_/S mux_bottom_ipin_10.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S mux_bottom_ipin_13.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S mux_bottom_ipin_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_13.mux_l3_in_1_/S
+ mux_bottom_ipin_13.mux_l4_in_0_/S mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_3.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S mux_bottom_ipin_12.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S mux_bottom_ipin_4.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_51_ chanx_right_in[0] chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0 mux_bottom_ipin_15.mux_l2_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S mux_bottom_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_10.mux_l2_in_1_/S
+ mux_bottom_ipin_10.mux_l3_in_1_/S mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_0.mux_l3_in_0_/S mux_bottom_ipin_0.mux_l4_in_0_/S
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34_ chanx_right_in[17] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_15.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_15.mux_l1_in_0_/X
+ mux_bottom_ipin_15.mux_l2_in_2_/S mux_bottom_ipin_15.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_15.mux_l4_in_0_/X top_grid_pin_31_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S mux_bottom_ipin_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0 mux_bottom_ipin_15.mux_l3_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17_ _17_/HI _17_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S mux_bottom_ipin_7.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_6.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_6.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0 mux_bottom_ipin_8.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S mux_bottom_ipin_8.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S mux_bottom_ipin_6.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_13.mux_l2_in_3_/S
+ mux_bottom_ipin_13.mux_l3_in_1_/S mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_3.mux_l3_in_0_/S mux_bottom_ipin_3.mux_l4_in_0_/S
+ mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_bottom_ipin_10.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_10.mux_l1_in_0_/S
+ mux_bottom_ipin_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_50_ chanx_right_in[1] chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1 mux_bottom_ipin_15.mux_l2_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_6.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_10.mux_l1_in_0_/S
+ mux_bottom_ipin_10.mux_l2_in_1_/S mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_0.mux_l2_in_0_/S mux_bottom_ipin_0.mux_l3_in_0_/S
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0 mux_bottom_ipin_6.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_33_ chanx_right_in[18] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_9.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_9.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0 mux_bottom_ipin_12.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1 mux_bottom_ipin_15.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_1.mux_l2_in_3_ _20_/HI chanx_right_in[17] mux_bottom_ipin_1.mux_l2_in_0_/S
+ mux_bottom_ipin_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_16_ _16_/HI _16_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0 mux_bottom_ipin_6.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_15.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_15.mux_l1_in_0_/S
+ mux_bottom_ipin_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_6.mux_l3_in_1_/S mux_bottom_ipin_6.mux_l4_in_0_/S
+ mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1 mux_bottom_ipin_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_7.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_1.mux_l4_in_0_ mux_bottom_ipin_1.mux_l3_in_1_/X mux_bottom_ipin_1.mux_l3_in_0_/X
+ mux_bottom_ipin_1.mux_l4_in_0_/S mux_bottom_ipin_1.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0 mux_bottom_ipin_10.mux_l2_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_13.mux_l1_in_1_/S
+ mux_bottom_ipin_13.mux_l2_in_3_/S mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_3.mux_l2_in_0_/S mux_bottom_ipin_3.mux_l3_in_0_/S
+ mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_8.mux_l4_in_0_/X top_grid_pin_24_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S mux_bottom_ipin_5.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_ipin_6.mux_l2_in_3_ _31_/HI chanx_right_in[18] mux_bottom_ipin_6.mux_l2_in_3_/S
+ mux_bottom_ipin_6.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_1.mux_l3_in_1_ mux_bottom_ipin_1.mux_l2_in_3_/X mux_bottom_ipin_1.mux_l2_in_2_/X
+ mux_bottom_ipin_1.mux_l3_in_1_/S mux_bottom_ipin_1.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0 mux_bottom_ipin_10.mux_l3_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_9.mux_l4_in_0_/S mux_bottom_ipin_10.mux_l1_in_0_/S
+ mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__dfxbp_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_0.mux_l1_in_1_/S mux_bottom_ipin_0.mux_l2_in_0_/S
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S mux_bottom_ipin_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1 mux_bottom_ipin_6.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_32_ chanx_right_in[19] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_ mux_bottom_ipin_9.mux_l3_in_1_/S mux_bottom_ipin_9.mux_l4_in_0_/S
+ mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S mux_bottom_ipin_14.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S mux_bottom_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1 mux_bottom_ipin_12.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_1.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_bottom_ipin_1.mux_l2_in_0_/S
+ mux_bottom_ipin_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_6.mux_l4_in_0_ mux_bottom_ipin_6.mux_l3_in_1_/X mux_bottom_ipin_6.mux_l3_in_0_/X
+ mux_bottom_ipin_6.mux_l4_in_0_/S mux_bottom_ipin_6.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1 mux_bottom_ipin_6.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_10.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_10.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_6.mux_l2_in_3_/S mux_bottom_ipin_6.mux_l3_in_1_/S
+ mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S mux_bottom_ipin_3.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_6.mux_l3_in_1_ mux_bottom_ipin_6.mux_l2_in_3_/X mux_bottom_ipin_6.mux_l2_in_2_/X
+ mux_bottom_ipin_6.mux_l3_in_1_/S mux_bottom_ipin_6.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S mux_bottom_ipin_9.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1 mux_bottom_ipin_10.mux_l2_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_12.mux_l4_in_0_/S
+ mux_bottom_ipin_13.mux_l1_in_1_/S mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_3.mux_l1_in_0_/S mux_bottom_ipin_3.mux_l2_in_0_/S
+ mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0 mux_bottom_ipin_1.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S mux_bottom_ipin_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S mux_bottom_ipin_2.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_6.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_bottom_ipin_6.mux_l2_in_3_/S
+ mux_bottom_ipin_6.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_ipin_1.mux_l3_in_0_ mux_bottom_ipin_1.mux_l2_in_1_/X mux_bottom_ipin_1.mux_l2_in_0_/X
+ mux_bottom_ipin_1.mux_l3_in_1_/S mux_bottom_ipin_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1 mux_bottom_ipin_10.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S mux_bottom_ipin_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_bottom_ipin_0.mux_l1_in_1_/S
+ mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_13.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_31_ _31_/HI _31_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0 mux_bottom_ipin_1.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_ipin_9.mux_l2_in_2_/S mux_bottom_ipin_9.mux_l3_in_1_/S
+ mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_1.mux_l2_in_1_ chanx_left_in[11] mux_bottom_ipin_1.mux_l1_in_2_/X
+ mux_bottom_ipin_1.mux_l2_in_0_/S mux_bottom_ipin_1.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1 mux_bottom_ipin_3.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_6.mux_l1_in_0_/S mux_bottom_ipin_6.mux_l2_in_3_/S
+ mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0 _17_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_1.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_bottom_ipin_1.mux_l1_in_2_/S
+ mux_bottom_ipin_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_6.mux_l3_in_0_ mux_bottom_ipin_6.mux_l2_in_1_/X mux_bottom_ipin_6.mux_l2_in_0_/X
+ mux_bottom_ipin_6.mux_l3_in_1_/S mux_bottom_ipin_6.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_2.mux_l4_in_0_/S mux_bottom_ipin_3.mux_l1_in_0_/S
+ mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_11.mux_l2_in_3_ _22_/HI chanx_right_in[15] mux_bottom_ipin_11.mux_l2_in_3_/S
+ mux_bottom_ipin_11.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1 mux_bottom_ipin_1.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_6.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_bottom_ipin_6.mux_l2_in_3_/S
+ mux_bottom_ipin_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S mux_bottom_ipin_1.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0 _23_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30_ _30_/HI _30_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1 mux_bottom_ipin_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_ipin_9.mux_l1_in_0_/S mux_bottom_ipin_9.mux_l2_in_2_/S
+ mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0 mux_bottom_ipin_14.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S mux_bottom_ipin_15.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_1.mux_l4_in_0_/X top_grid_pin_17_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_11.mux_l4_in_0_ mux_bottom_ipin_11.mux_l3_in_1_/X mux_bottom_ipin_11.mux_l3_in_0_/X
+ mux_bottom_ipin_11.mux_l4_in_0_/S mux_bottom_ipin_11.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_1.mux_l2_in_0_ mux_bottom_ipin_1.mux_l1_in_1_/X mux_bottom_ipin_1.mux_l1_in_0_/X
+ mux_bottom_ipin_1.mux_l2_in_0_/S mux_bottom_ipin_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S mux_bottom_ipin_10.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S mux_bottom_ipin_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_5.mux_l4_in_0_/S mux_bottom_ipin_6.mux_l1_in_0_/S
+ mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_11.mux_l3_in_1_ mux_bottom_ipin_11.mux_l2_in_3_/X mux_bottom_ipin_11.mux_l2_in_2_/X
+ mux_bottom_ipin_11.mux_l3_in_0_/S mux_bottom_ipin_11.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S mux_bottom_ipin_14.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_1.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_bottom_ipin_1.mux_l1_in_2_/S
+ mux_bottom_ipin_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__33__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_11.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_bottom_ipin_11.mux_l2_in_3_/S
+ mux_bottom_ipin_11.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S mux_bottom_ipin_15.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S mux_bottom_ipin_13.mux_l4_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S mux_bottom_ipin_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_ chanx_left_in[2] mux_bottom_ipin_6.mux_l1_in_0_/X
+ mux_bottom_ipin_6.mux_l2_in_3_/S mux_bottom_ipin_6.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__41__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S mux_bottom_ipin_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_ipin_8.mux_l4_in_0_/S mux_bottom_ipin_9.mux_l1_in_0_/S
+ mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1 mux_bottom_ipin_14.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S mux_bottom_ipin_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__36__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0 mux_bottom_ipin_5.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_ipin_11.mux_l3_in_0_ mux_bottom_ipin_11.mux_l2_in_1_/X mux_bottom_ipin_11.mux_l2_in_0_/X
+ mux_bottom_ipin_11.mux_l3_in_0_/S mux_bottom_ipin_11.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_1.mux_l1_in_2_/S
+ mux_bottom_ipin_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__44__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_11.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_bottom_ipin_11.mux_l2_in_3_/S
+ mux_bottom_ipin_11.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__39__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1 mux_bottom_ipin_5.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S mux_bottom_ipin_12.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_ipin_6.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_6.mux_l1_in_0_/S
+ mux_bottom_ipin_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__52__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1 mux_bottom_ipin_5.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_6.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S mux_bottom_ipin_11.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__47__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_11.mux_l4_in_0_/X top_grid_pin_27_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S mux_bottom_ipin_10.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__60__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_11.mux_l2_in_0_ chanx_left_in[3] mux_bottom_ipin_11.mux_l1_in_0_/X
+ mux_bottom_ipin_11.mux_l2_in_3_/S mux_bottom_ipin_11.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__55__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0 mux_bottom_ipin_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S mux_bottom_ipin_11.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S mux_bottom_ipin_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S mux_bottom_ipin_15.mux_l3_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__63__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S mux_bottom_ipin_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0 mux_bottom_ipin_9.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S mux_bottom_ipin_6.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__58__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1 mux_bottom_ipin_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__71__A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0 mux_bottom_ipin_7.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S mux_bottom_ipin_9.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1 mux_bottom_ipin_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0 mux_bottom_ipin_13.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__66__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_11.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_bottom_ipin_11.mux_l1_in_0_/S
+ mux_bottom_ipin_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0 mux_bottom_ipin_7.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_4.mux_l4_in_0_/X top_grid_pin_20_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_69_ chanx_left_in[2] chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1 mux_bottom_ipin_9.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0 mux_bottom_ipin_11.mux_l2_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_2.mux_l2_in_3_ _27_/HI chanx_right_in[14] mux_bottom_ipin_2.mux_l2_in_3_/S
+ mux_bottom_ipin_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S mux_bottom_ipin_13.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__69__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0 mux_bottom_ipin_11.mux_l3_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1 mux_bottom_ipin_7.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_2.mux_l4_in_0_ mux_bottom_ipin_2.mux_l3_in_1_/X mux_bottom_ipin_2.mux_l3_in_0_/X
+ mux_bottom_ipin_2.mux_l4_in_0_/S mux_bottom_ipin_2.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S mux_bottom_ipin_12.mux_l2_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1 mux_bottom_ipin_13.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S mux_bottom_ipin_8.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_7.mux_l2_in_3_ _16_/HI chanx_right_in[19] mux_bottom_ipin_7.mux_l2_in_1_/S
+ mux_bottom_ipin_7.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1 mux_bottom_ipin_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0 mux_bottom_ipin_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1 chanx_right_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_2.mux_l3_in_1_ mux_bottom_ipin_2.mux_l2_in_3_/X mux_bottom_ipin_2.mux_l2_in_2_/X
+ mux_bottom_ipin_2.mux_l3_in_1_/S mux_bottom_ipin_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_68_ chanx_left_in[3] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S mux_bottom_ipin_11.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S mux_bottom_ipin_7.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1 mux_bottom_ipin_11.mux_l2_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_2.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_bottom_ipin_2.mux_l2_in_3_/S
+ mux_bottom_ipin_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_ipin_7.mux_l4_in_0_ mux_bottom_ipin_7.mux_l3_in_1_/X mux_bottom_ipin_7.mux_l3_in_0_/X
+ mux_bottom_ipin_7.mux_l4_in_0_/S mux_bottom_ipin_7.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0 mux_bottom_ipin_2.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S mux_bottom_ipin_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1 mux_bottom_ipin_11.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S mux_bottom_ipin_6.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_7.mux_l3_in_1_ mux_bottom_ipin_7.mux_l2_in_3_/X mux_bottom_ipin_7.mux_l2_in_2_/X
+ mux_bottom_ipin_7.mux_l3_in_0_/S mux_bottom_ipin_7.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0 mux_bottom_ipin_2.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S mux_bottom_ipin_7.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1 mux_bottom_ipin_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_7.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_bottom_ipin_7.mux_l2_in_1_/S
+ mux_bottom_ipin_7.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S mux_bottom_ipin_5.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_ipin_2.mux_l3_in_0_ mux_bottom_ipin_2.mux_l2_in_1_/X mux_bottom_ipin_2.mux_l2_in_0_/X
+ mux_bottom_ipin_2.mux_l3_in_1_/S mux_bottom_ipin_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0 _18_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_67_ chanx_left_in[4] chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_2.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_bottom_ipin_2.mux_l2_in_3_/S
+ mux_bottom_ipin_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1 mux_bottom_ipin_2.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_14.mux_l4_in_0_/X top_grid_pin_30_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_ipin_14.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_ipin_7.mux_l3_in_0_ mux_bottom_ipin_7.mux_l2_in_1_/X mux_bottom_ipin_7.mux_l2_in_0_/X
+ mux_bottom_ipin_7.mux_l3_in_0_/S mux_bottom_ipin_7.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0 _24_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1 mux_bottom_ipin_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D mux_bottom_ipin_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0 mux_bottom_ipin_15.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

