* NGSPICE file created from sb_3__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

.subckt sb_3__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ bottom_right_grid_pin_13_
+ bottom_right_grid_pin_15_ bottom_right_grid_pin_1_ bottom_right_grid_pin_3_ bottom_right_grid_pin_5_
+ bottom_right_grid_pin_7_ bottom_right_grid_pin_9_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_12_ left_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ top_right_grid_pin_13_ top_right_grid_pin_15_ top_right_grid_pin_1_ top_right_grid_pin_3_
+ top_right_grid_pin_5_ top_right_grid_pin_7_ top_right_grid_pin_9_ vpwr vgnd
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_111 vgnd vpwr scs8hd_decap_8
XFILLER_26_74 vgnd vpwr scs8hd_fill_1
XFILLER_9_137 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_1_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _26_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_76 vgnd vpwr scs8hd_decap_12
XFILLER_33_217 vgnd vpwr scs8hd_fill_1
XFILLER_5_184 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _16_/HI mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_15_217 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _43_/A vgnd vpwr scs8hd_inv_1
X_49_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_30 vgnd vpwr scs8hd_fill_1
XFILLER_34_96 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_6 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _24_/HI mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_fill_1
XFILLER_19_172 vgnd vpwr scs8hd_decap_8
XFILLER_26_109 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_10 vgnd vpwr scs8hd_decap_4
XFILLER_15_21 vgnd vpwr scs8hd_decap_12
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _16_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_3
XFILLER_26_97 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vgnd vpwr scs8hd_decap_4
XFILLER_3_57 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_204 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _18_/HI mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_66 vgnd vpwr scs8hd_fill_1
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _32_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_204 vgnd vpwr scs8hd_decap_8
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XFILLER_5_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_2_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vgnd vpwr scs8hd_decap_8
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
X_48_ _48_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _36_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_11_210 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_206 vgnd vpwr scs8hd_decap_8
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_31 vgnd vpwr scs8hd_decap_12
XFILLER_29_75 vgnd vpwr scs8hd_decap_4
XFILLER_6_46 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_15_33 vgnd vpwr scs8hd_decap_12
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_8
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_31_157 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_190 vgnd vpwr scs8hd_decap_8
XFILLER_7_9 vpwr vgnd scs8hd_fill_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_69 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _39_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_216 vgnd vpwr scs8hd_fill_1
XFILLER_8_194 vpwr vgnd scs8hd_fill_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_216 vpwr vgnd scs8hd_fill_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XFILLER_9_68 vpwr vgnd scs8hd_fill_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
X_47_ _47_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_204 vpwr vgnd scs8hd_fill_2
XFILLER_29_119 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XFILLER_29_43 vgnd vpwr scs8hd_decap_12
XFILLER_29_87 vgnd vpwr scs8hd_decap_12
XFILLER_6_58 vgnd vpwr scs8hd_fill_1
XFILLER_6_36 vgnd vpwr scs8hd_fill_1
XFILLER_15_45 vgnd vpwr scs8hd_decap_12
XFILLER_16_199 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_147 vgnd vpwr scs8hd_decap_3
XFILLER_31_169 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_90 vgnd vpwr scs8hd_decap_4
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_169 vpwr vgnd scs8hd_fill_2
XFILLER_21_180 vgnd vpwr scs8hd_decap_3
XFILLER_3_26 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_162 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_35 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_209 vgnd vpwr scs8hd_decap_8
XFILLER_5_110 vgnd vpwr scs8hd_decap_4
XFILLER_5_143 vpwr vgnd scs8hd_fill_2
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XFILLER_15_209 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_16 vgnd vpwr scs8hd_decap_4
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
X_46_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_20_201 vgnd vpwr scs8hd_decap_12
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_216 vpwr vgnd scs8hd_fill_2
X_29_ _29_/HI _29_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_55 vgnd vpwr scs8hd_decap_4
XFILLER_29_66 vgnd vpwr scs8hd_fill_1
XFILLER_29_99 vgnd vpwr scs8hd_decap_12
XFILLER_34_189 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_57 vgnd vpwr scs8hd_decap_4
XFILLER_0_200 vgnd vpwr scs8hd_fill_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_21_192 vgnd vpwr scs8hd_decap_3
XFILLER_3_38 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_130 vgnd vpwr scs8hd_decap_8
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_47 vgnd vpwr scs8hd_decap_3
XFILLER_5_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_210 vgnd vpwr scs8hd_decap_8
XFILLER_2_114 vgnd vpwr scs8hd_decap_8
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_48 vgnd vpwr scs8hd_decap_12
X_45_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_9_ mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_213 vgnd vpwr scs8hd_fill_1
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_28_ _28_/HI _28_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _19_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_124 vgnd vpwr scs8hd_decap_8
XFILLER_34_135 vgnd vpwr scs8hd_decap_12
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XFILLER_0_212 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_190 vgnd vpwr scs8hd_decap_8
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_68 vgnd vpwr scs8hd_decap_6
XFILLER_9_109 vpwr vgnd scs8hd_fill_2
XANTENNA__31__A _31_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XFILLER_12_193 vgnd vpwr scs8hd_decap_8
XFILLER_27_208 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_59 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_137 vgnd vpwr scs8hd_decap_12
XFILLER_2_126 vpwr vgnd scs8hd_fill_2
X_44_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_83 vgnd vpwr scs8hd_fill_1
X_27_ _27_/HI _27_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XANTENNA__34__A _34_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_155 vgnd vpwr scs8hd_decap_3
XFILLER_34_147 vgnd vpwr scs8hd_decap_6
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_128 vpwr vgnd scs8hd_fill_2
XFILLER_21_150 vgnd vpwr scs8hd_decap_8
XFILLER_21_172 vgnd vpwr scs8hd_decap_8
XFILLER_3_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_8
XFILLER_12_150 vgnd vpwr scs8hd_decap_3
XANTENNA__42__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__37__A _37_/A vgnd vpwr scs8hd_diode_2
X_43_ _43_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_1_193 vgnd vpwr scs8hd_decap_6
XFILLER_20_215 vgnd vpwr scs8hd_decap_3
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_208 vgnd vpwr scs8hd_decap_8
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_3
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
X_26_ _26_/HI _26_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__50__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_25_159 vgnd vpwr scs8hd_decap_12
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_192 vgnd vpwr scs8hd_fill_1
XFILLER_0_203 vgnd vpwr scs8hd_fill_1
XFILLER_16_126 vgnd vpwr scs8hd_decap_12
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__45__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_92 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_94 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_184 vgnd vpwr scs8hd_decap_8
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_188 vgnd vpwr scs8hd_decap_4
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_35_210 vgnd vpwr scs8hd_decap_8
XFILLER_12_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_147 vgnd vpwr scs8hd_decap_8
XFILLER_5_136 vgnd vpwr scs8hd_decap_4
XFILLER_4_62 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_202 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XANTENNA__53__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_7 vgnd vpwr scs8hd_decap_12
X_42_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA__48__A _48_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_25_ _25_/HI _25_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_17 vpwr vgnd scs8hd_fill_2
XFILLER_18_190 vgnd vpwr scs8hd_decap_8
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XFILLER_16_138 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _28_/HI mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/TEB
+ mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_22_108 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_119 vgnd vpwr scs8hd_decap_3
XANTENNA__56__A _56_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_178 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _38_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_162 vpwr vgnd scs8hd_fill_2
XFILLER_1_151 vpwr vgnd scs8hd_fill_2
X_41_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_9_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_20 vgnd vpwr scs8hd_decap_4
XFILLER_1_31 vgnd vpwr scs8hd_decap_4
X_24_ _24_/HI _24_/LO vgnd vpwr scs8hd_conb_1
XFILLER_34_6 vgnd vpwr scs8hd_decap_12
XFILLER_1_75 vgnd vpwr scs8hd_decap_8
XFILLER_36_180 vgnd vpwr scs8hd_decap_6
XFILLER_19_103 vpwr vgnd scs8hd_fill_2
XFILLER_19_147 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _20_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_150 vgnd vpwr scs8hd_decap_6
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_6
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _17_/HI mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_120 vpwr vgnd scs8hd_fill_2
XFILLER_12_142 vgnd vpwr scs8hd_decap_8
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_116 vgnd vpwr scs8hd_decap_4
XFILLER_27_60 vgnd vpwr scs8hd_fill_1
XFILLER_27_82 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_7_ mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_215 vgnd vpwr scs8hd_decap_3
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_13_73 vgnd vpwr scs8hd_decap_3
XFILLER_13_84 vpwr vgnd scs8hd_fill_2
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
X_40_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_13_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_54 vgnd vpwr scs8hd_fill_1
X_23_ _23_/HI _23_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_107 vgnd vpwr scs8hd_decap_12
XFILLER_33_184 vpwr vgnd scs8hd_fill_2
XFILLER_33_195 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_95 vgnd vpwr scs8hd_fill_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XFILLER_7_86 vpwr vgnd scs8hd_fill_2
XFILLER_30_198 vgnd vpwr scs8hd_decap_3
XFILLER_21_121 vgnd vpwr scs8hd_fill_1
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XFILLER_12_176 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_191 vpwr vgnd scs8hd_fill_2
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_94 vgnd vpwr scs8hd_decap_12
XFILLER_4_194 vgnd vpwr scs8hd_decap_3
XFILLER_4_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_30 vgnd vpwr scs8hd_decap_12
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_18 vgnd vpwr scs8hd_decap_12
XFILLER_1_99 vgnd vpwr scs8hd_decap_4
X_22_ _22_/HI _22_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XFILLER_3_204 vpwr vgnd scs8hd_fill_2
XFILLER_10_42 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_171 vgnd vpwr scs8hd_decap_12
XFILLER_34_108 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_119 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_141 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_130 vgnd vpwr scs8hd_decap_12
XFILLER_7_43 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_200 vgnd vpwr scs8hd_fill_1
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XFILLER_12_166 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XFILLER_17_203 vgnd vpwr scs8hd_decap_12
XFILLER_32_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_42 vgnd vpwr scs8hd_decap_4
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_9 vgnd vpwr scs8hd_fill_1
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_1_12 vgnd vpwr scs8hd_fill_1
XFILLER_27_8 vgnd vpwr scs8hd_decap_12
X_21_ _21_/HI _21_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _29_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
XFILLER_29_19 vgnd vpwr scs8hd_decap_12
XFILLER_3_216 vpwr vgnd scs8hd_fill_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_6
XFILLER_10_54 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_150 vgnd vpwr scs8hd_decap_3
XFILLER_33_131 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_86 vgnd vpwr scs8hd_decap_6
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_142 vgnd vpwr scs8hd_decap_12
XFILLER_15_175 vgnd vpwr scs8hd_decap_6
XFILLER_15_197 vgnd vpwr scs8hd_decap_4
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_3
XFILLER_17_215 vgnd vpwr scs8hd_decap_3
XFILLER_27_52 vpwr vgnd scs8hd_fill_2
XFILLER_4_130 vgnd vpwr scs8hd_decap_4
XFILLER_4_174 vgnd vpwr scs8hd_decap_12
XFILLER_4_163 vgnd vpwr scs8hd_decap_8
XFILLER_4_45 vgnd vpwr scs8hd_decap_8
XFILLER_4_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_111 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_75 vgnd vpwr scs8hd_decap_12
X_20_ _20_/HI _20_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_35 vgnd vpwr scs8hd_fill_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_66 vgnd vpwr scs8hd_decap_4
XFILLER_19_107 vgnd vpwr scs8hd_decap_12
XFILLER_19_86 vgnd vpwr scs8hd_decap_6
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _21_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XFILLER_24_198 vgnd vpwr scs8hd_decap_3
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_121 vgnd vpwr scs8hd_fill_1
XFILLER_15_154 vgnd vpwr scs8hd_decap_6
XFILLER_7_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_135 vgnd vpwr scs8hd_fill_1
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_20 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_186 vgnd vpwr scs8hd_decap_8
XFILLER_4_79 vgnd vpwr scs8hd_decap_12
XFILLER_14_208 vgnd vpwr scs8hd_decap_6
XFILLER_13_88 vgnd vpwr scs8hd_decap_4
XFILLER_13_99 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_3
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_87 vgnd vpwr scs8hd_decap_4
XFILLER_19_119 vgnd vpwr scs8hd_decap_3
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _29_/HI mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/TEB
+ mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_188 vgnd vpwr scs8hd_decap_4
XFILLER_33_199 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_90 vpwr vgnd scs8hd_fill_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_7_13 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _47_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_103 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_158 vgnd vpwr scs8hd_decap_3
XFILLER_29_203 vgnd vpwr scs8hd_decap_12
XFILLER_12_125 vgnd vpwr scs8hd_decap_8
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_35_206 vpwr vgnd scs8hd_fill_2
XFILLER_7_162 vgnd vpwr scs8hd_fill_1
XFILLER_27_32 vgnd vpwr scs8hd_decap_12
XFILLER_27_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_78 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_201 vgnd vpwr scs8hd_decap_12
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_48 vgnd vpwr scs8hd_decap_6
XFILLER_3_208 vgnd vpwr scs8hd_decap_8
XFILLER_10_79 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_8
XFILLER_33_134 vgnd vpwr scs8hd_decap_4
XFILLER_33_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_115 vgnd vpwr scs8hd_decap_6
XFILLER_29_215 vgnd vpwr scs8hd_decap_3
XFILLER_8_119 vgnd vpwr scs8hd_decap_8
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_16_78 vgnd vpwr scs8hd_decap_12
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_44 vgnd vpwr scs8hd_decap_8
XFILLER_4_15 vgnd vpwr scs8hd_decap_4
XFILLER_31_210 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_13 vgnd vpwr scs8hd_decap_6
XFILLER_13_46 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vgnd vpwr scs8hd_decap_8
XFILLER_1_147 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_3 vgnd vpwr scs8hd_decap_6
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_16 vpwr vgnd scs8hd_fill_2
XFILLER_1_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_38 vgnd vpwr scs8hd_fill_1
XFILLER_36_187 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XFILLER_18_198 vgnd vpwr scs8hd_decap_3
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _31_/A vgnd vpwr scs8hd_inv_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_26 vgnd vpwr scs8hd_decap_6
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_30_7 vgnd vpwr scs8hd_decap_12
XFILLER_21_138 vgnd vpwr scs8hd_decap_12
XFILLER_16_68 vgnd vpwr scs8hd_decap_6
XFILLER_8_109 vgnd vpwr scs8hd_fill_1
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _35_/A vgnd vpwr scs8hd_inv_1
XFILLER_7_120 vpwr vgnd scs8hd_fill_2
XFILLER_7_142 vpwr vgnd scs8hd_fill_2
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _52_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_56 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_115 vgnd vpwr scs8hd_decap_4
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_81 vgnd vpwr scs8hd_fill_1
XFILLER_24_68 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_199 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _22_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_180 vgnd vpwr scs8hd_decap_12
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_80 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_161 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_165 vgnd vpwr scs8hd_decap_12
XFILLER_7_187 vpwr vgnd scs8hd_fill_2
XFILLER_11_161 vgnd vpwr scs8hd_decap_3
XFILLER_14_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_12
XANTENNA__32__A _32_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_205 vgnd vpwr scs8hd_decap_12
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.INVTX1_2_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_156 vgnd vpwr scs8hd_decap_12
XFILLER_10_16 vgnd vpwr scs8hd_decap_12
XFILLER_10_38 vgnd vpwr scs8hd_fill_1
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_3_ mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__40__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XFILLER_2_61 vgnd vpwr scs8hd_decap_8
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_192 vgnd vpwr scs8hd_decap_4
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _22_/HI mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_126 vpwr vgnd scs8hd_fill_2
XANTENNA__35__A _35_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_7_39 vpwr vgnd scs8hd_fill_2
XFILLER_7_177 vpwr vgnd scs8hd_fill_2
XFILLER_22_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_93 vgnd vpwr scs8hd_fill_1
XFILLER_25_210 vgnd vpwr scs8hd_decap_8
XFILLER_27_69 vpwr vgnd scs8hd_fill_2
XFILLER_4_114 vgnd vpwr scs8hd_decap_3
XFILLER_17_91 vpwr vgnd scs8hd_fill_2
XFILLER_33_90 vgnd vpwr scs8hd_decap_3
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vgnd vpwr scs8hd_fill_1
XANTENNA__43__A _43_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_217 vgnd vpwr scs8hd_fill_1
XFILLER_0_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA__38__A _38_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_36_168 vgnd vpwr scs8hd_decap_12
XFILLER_10_28 vgnd vpwr scs8hd_decap_3
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_35_190 vgnd vpwr scs8hd_fill_1
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_212 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_102 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_190 vgnd vpwr scs8hd_decap_8
XFILLER_33_138 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XFILLER_15_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__51__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_11_60 vgnd vpwr scs8hd_fill_1
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_108 vgnd vpwr scs8hd_decap_12
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XANTENNA__46__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_112 vgnd vpwr scs8hd_decap_8
XFILLER_7_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_137 vgnd vpwr scs8hd_decap_12
XFILLER_4_126 vpwr vgnd scs8hd_fill_2
XFILLER_4_19 vgnd vpwr scs8hd_fill_1
XFILLER_17_70 vgnd vpwr scs8hd_fill_1
XFILLER_3_181 vpwr vgnd scs8hd_fill_2
XFILLER_1_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__54__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_36_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_147 vgnd vpwr scs8hd_decap_12
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XANTENNA__49__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_18_114 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _15_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_70 vgnd vpwr scs8hd_decap_3
X_56_ _56_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XFILLER_15_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_39_ _39_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_7_146 vgnd vpwr scs8hd_decap_12
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_73 vgnd vpwr scs8hd_decap_8
XFILLER_8_84 vgnd vpwr scs8hd_decap_8
XFILLER_4_149 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_3
XFILLER_1_119 vgnd vpwr scs8hd_fill_1
XFILLER_0_196 vgnd vpwr scs8hd_decap_4
XFILLER_28_70 vgnd vpwr scs8hd_fill_1
XFILLER_5_85 vpwr vgnd scs8hd_fill_2
XFILLER_5_200 vpwr vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_36_137 vgnd vpwr scs8hd_decap_12
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_159 vgnd vpwr scs8hd_decap_12
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_126 vgnd vpwr scs8hd_decap_12
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_33_107 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _48_/A vgnd vpwr scs8hd_inv_1
X_55_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_62 vgnd vpwr scs8hd_decap_4
XFILLER_11_84 vpwr vgnd scs8hd_fill_2
X_38_ _38_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_16_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_154 vgnd vpwr scs8hd_decap_4
XFILLER_20_165 vgnd vpwr scs8hd_decap_12
XFILLER_11_121 vgnd vpwr scs8hd_fill_1
XFILLER_7_158 vgnd vpwr scs8hd_decap_4
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _21_/HI mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_41 vgnd vpwr scs8hd_decap_8
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_60 vgnd vpwr scs8hd_fill_1
XFILLER_33_82 vgnd vpwr scs8hd_decap_8
XFILLER_13_205 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _18_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_164 vgnd vpwr scs8hd_decap_4
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_75 vgnd vpwr scs8hd_decap_6
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_42 vgnd vpwr scs8hd_decap_4
XFILLER_5_20 vpwr vgnd scs8hd_fill_2
XFILLER_6_9 vgnd vpwr scs8hd_fill_1
XFILLER_14_51 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_35_182 vgnd vpwr scs8hd_fill_1
XFILLER_2_215 vgnd vpwr scs8hd_decap_3
XFILLER_2_204 vgnd vpwr scs8hd_decap_8
XFILLER_18_138 vgnd vpwr scs8hd_decap_12
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_25_72 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_33_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_43 vgnd vpwr scs8hd_decap_12
XFILLER_2_32 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_3_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_54_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XFILLER_32_163 vgnd vpwr scs8hd_decap_8
XFILLER_32_196 vgnd vpwr scs8hd_fill_1
XFILLER_23_152 vgnd vpwr scs8hd_decap_4
XFILLER_23_163 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _15_/HI mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/TEB
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_23_196 vgnd vpwr scs8hd_decap_3
XFILLER_2_3 vgnd vpwr scs8hd_decap_6
XFILLER_11_52 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_174 vpwr vgnd scs8hd_fill_2
XFILLER_14_196 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
X_37_ _37_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_20_177 vgnd vpwr scs8hd_decap_12
XFILLER_8_97 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_8
XFILLER_17_95 vgnd vpwr scs8hd_decap_4
XFILLER_3_184 vgnd vpwr scs8hd_decap_6
XFILLER_3_173 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_217 vgnd vpwr scs8hd_fill_1
XFILLER_0_176 vgnd vpwr scs8hd_decap_8
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _33_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_62 vgnd vpwr scs8hd_decap_12
XFILLER_36_106 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_1_ mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_106 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_7_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_62 vgnd vpwr scs8hd_decap_8
XFILLER_25_95 vgnd vpwr scs8hd_decap_12
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_2_55 vpwr vgnd scs8hd_fill_2
X_53_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _37_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_175 vgnd vpwr scs8hd_decap_8
XFILLER_11_20 vgnd vpwr scs8hd_decap_6
XFILLER_11_42 vgnd vpwr scs8hd_decap_8
XFILLER_36_94 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_36_ _36_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_3
XFILLER_20_189 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_101 vgnd vpwr scs8hd_decap_12
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
XFILLER_22_96 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_3
XFILLER_8_10 vgnd vpwr scs8hd_decap_4
XFILLER_8_21 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_19_ _19_/HI _19_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_3
XFILLER_17_74 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_95 vgnd vpwr scs8hd_decap_12
XFILLER_3_152 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_207 vgnd vpwr scs8hd_decap_6
XFILLER_0_111 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_118 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_195 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vgnd vpwr scs8hd_decap_8
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XFILLER_2_78 vgnd vpwr scs8hd_decap_12
X_52_ _52_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_143 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
X_35_ _35_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
XFILLER_7_106 vgnd vpwr scs8hd_decap_4
XFILLER_11_113 vgnd vpwr scs8hd_decap_8
XFILLER_11_135 vgnd vpwr scs8hd_decap_3
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
X_18_ _18_/HI _18_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_205 vgnd vpwr scs8hd_decap_8
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_6
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
XFILLER_12_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _20_/HI mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_134 vgnd vpwr scs8hd_decap_8
XFILLER_0_145 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_52 vpwr vgnd scs8hd_fill_2
XFILLER_28_74 vgnd vpwr scs8hd_decap_12
XFILLER_5_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_204 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_86 vgnd vpwr scs8hd_decap_6
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_152 vgnd vpwr scs8hd_decap_8
XFILLER_35_163 vpwr vgnd scs8hd_fill_2
XFILLER_35_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_51_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_17_163 vpwr vgnd scs8hd_fill_2
XFILLER_17_174 vpwr vgnd scs8hd_fill_2
XFILLER_32_144 vgnd vpwr scs8hd_decap_8
XFILLER_11_66 vgnd vpwr scs8hd_fill_1
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_63 vgnd vpwr scs8hd_decap_12
XFILLER_14_166 vgnd vpwr scs8hd_decap_8
X_34_ _34_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_9_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_129 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_206 vgnd vpwr scs8hd_decap_8
XFILLER_6_162 vgnd vpwr scs8hd_decap_12
XFILLER_33_3 vpwr vgnd scs8hd_fill_2
X_17_ _17_/HI _17_/LO vgnd vpwr scs8hd_conb_1
XFILLER_33_20 vgnd vpwr scs8hd_decap_12
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_143 vpwr vgnd scs8hd_fill_2
XFILLER_3_132 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_90 vgnd vpwr scs8hd_fill_1
XFILLER_13_209 vgnd vpwr scs8hd_decap_8
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_86 vgnd vpwr scs8hd_decap_6
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _23_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_24 vgnd vpwr scs8hd_decap_3
XFILLER_14_44 vgnd vpwr scs8hd_decap_3
XFILLER_5_216 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_50_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_131 vgnd vpwr scs8hd_decap_12
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_75 vgnd vpwr scs8hd_decap_12
X_33_ _33_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_9_160 vgnd vpwr scs8hd_fill_1
XFILLER_28_215 vgnd vpwr scs8hd_decap_3
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_215 vgnd vpwr scs8hd_decap_3
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_174 vgnd vpwr scs8hd_decap_8
XFILLER_6_185 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_16_ _16_/HI _16_/LO vgnd vpwr scs8hd_conb_1
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_32 vgnd vpwr scs8hd_decap_12
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_103 vgnd vpwr scs8hd_decap_8
XFILLER_28_21 vgnd vpwr scs8hd_decap_8
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_14 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _27_/HI mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/TEB
+ mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_26_121 vgnd vpwr scs8hd_decap_12
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XFILLER_26_198 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XFILLER_17_143 vgnd vpwr scs8hd_decap_12
XFILLER_17_187 vgnd vpwr scs8hd_decap_6
XFILLER_17_198 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_135 vgnd vpwr scs8hd_decap_8
XFILLER_36_87 vgnd vpwr scs8hd_decap_6
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_135 vgnd vpwr scs8hd_decap_12
XFILLER_14_179 vgnd vpwr scs8hd_decap_8
X_32_ _32_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XFILLER_11_127 vgnd vpwr scs8hd_decap_6
XFILLER_11_149 vgnd vpwr scs8hd_decap_12
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_15_ mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_58 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_15_ _15_/HI _15_/LO vgnd vpwr scs8hd_conb_1
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_78 vpwr vgnd scs8hd_fill_2
XFILLER_33_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_167 vgnd vpwr scs8hd_decap_4
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
XFILLER_3_112 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_8
XFILLER_8_215 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_13 vgnd vpwr scs8hd_decap_12
XFILLER_14_68 vgnd vpwr scs8hd_decap_8
XFILLER_14_79 vgnd vpwr scs8hd_decap_12
XFILLER_30_56 vgnd vpwr scs8hd_decap_3
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _19_/HI mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_5_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_199 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_26_133 vgnd vpwr scs8hd_decap_12
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XFILLER_1_210 vgnd vpwr scs8hd_decap_8
XFILLER_17_155 vgnd vpwr scs8hd_decap_4
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
XFILLER_2_9 vgnd vpwr scs8hd_fill_1
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vgnd vpwr scs8hd_fill_1
XFILLER_14_147 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_31_ _31_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
XFILLER_9_184 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _24_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_56 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_205 vgnd vpwr scs8hd_decap_8
XFILLER_12_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_49 vpwr vgnd scs8hd_fill_2
XFILLER_5_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_25 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_35_167 vgnd vpwr scs8hd_decap_4
XFILLER_35_178 vgnd vpwr scs8hd_decap_4
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_26_145 vgnd vpwr scs8hd_decap_8
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XANTENNA__30__A _30_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_167 vgnd vpwr scs8hd_decap_4
XFILLER_17_178 vgnd vpwr scs8hd_decap_4
XFILLER_23_104 vgnd vpwr scs8hd_decap_12
XFILLER_23_148 vpwr vgnd scs8hd_fill_2
XFILLER_23_159 vpwr vgnd scs8hd_fill_2
XFILLER_11_26 vgnd vpwr scs8hd_fill_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_30_ _30_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_28_9 vgnd vpwr scs8hd_decap_12
XFILLER_20_129 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_207 vgnd vpwr scs8hd_decap_8
XFILLER_10_173 vgnd vpwr scs8hd_decap_8
XFILLER_10_184 vgnd vpwr scs8hd_decap_8
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_103 vgnd vpwr scs8hd_fill_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_3
XFILLER_2_191 vgnd vpwr scs8hd_decap_8
XFILLER_2_180 vgnd vpwr scs8hd_decap_8
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_81 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__33__A _33_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_5_ mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XFILLER_35_135 vgnd vpwr scs8hd_decap_6
XFILLER_6_93 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _56_/A vgnd vpwr scs8hd_inv_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_17_102 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_23_116 vgnd vpwr scs8hd_decap_6
XFILLER_31_193 vgnd vpwr scs8hd_decap_4
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XANTENNA__41__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_22_171 vgnd vpwr scs8hd_decap_12
XFILLER_9_153 vgnd vpwr scs8hd_fill_1
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA__36__A _36_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_17 vpwr vgnd scs8hd_fill_2
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XFILLER_6_123 vgnd vpwr scs8hd_decap_8
XFILLER_6_134 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _26_/HI mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_80 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _30_/A vgnd vpwr scs8hd_inv_1
XFILLER_28_58 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_111 vgnd vpwr scs8hd_decap_8
XANTENNA__44__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _34_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_2_19 vgnd vpwr scs8hd_decap_12
XANTENNA__39__A _39_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_81 vgnd vpwr scs8hd_decap_12
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_191 vgnd vpwr scs8hd_decap_8
XFILLER_31_161 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_8
XFILLER_22_183 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_165 vpwr vgnd scs8hd_fill_2
XFILLER_3_95 vgnd vpwr scs8hd_decap_8
XFILLER_3_73 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XFILLER_8_29 vpwr vgnd scs8hd_fill_2
XANTENNA__52__A _52_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_146 vgnd vpwr scs8hd_decap_6
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_15_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_116 vgnd vpwr scs8hd_fill_1
XANTENNA__47__A _47_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_204 vpwr vgnd scs8hd_fill_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_3
XFILLER_23_70 vpwr vgnd scs8hd_fill_2
XFILLER_23_92 vgnd vpwr scs8hd_decap_12
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_4
XFILLER_12_204 vgnd vpwr scs8hd_decap_8
XFILLER_12_215 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _27_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XFILLER_6_62 vgnd vpwr scs8hd_decap_8
XFILLER_6_73 vgnd vpwr scs8hd_decap_8
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XFILLER_17_159 vgnd vpwr scs8hd_fill_1
XANTENNA__55__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_93 vgnd vpwr scs8hd_decap_12
XFILLER_25_192 vgnd vpwr scs8hd_decap_3
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XFILLER_31_173 vgnd vpwr scs8hd_decap_8
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_140 vgnd vpwr scs8hd_decap_12
XFILLER_22_195 vgnd vpwr scs8hd_decap_12
XFILLER_7_3 vgnd vpwr scs8hd_decap_3
XFILLER_9_188 vpwr vgnd scs8hd_fill_2
XFILLER_13_173 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_13_ mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _25_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_158 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_213 vgnd vpwr scs8hd_decap_4
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/TEB mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_17_127 vpwr vgnd scs8hd_fill_2
XFILLER_25_171 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_9_123 vgnd vpwr scs8hd_decap_3
XFILLER_13_141 vgnd vpwr scs8hd_decap_12
XFILLER_9_156 vgnd vpwr scs8hd_decap_4
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_42 vgnd vpwr scs8hd_decap_8
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _28_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_5_192 vgnd vpwr scs8hd_fill_1
XFILLER_5_170 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/TEB mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vgnd vpwr scs8hd_decap_8
XFILLER_21_206 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _25_/HI mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_83 vgnd vpwr scs8hd_decap_8
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_71 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XFILLER_17_106 vgnd vpwr scs8hd_decap_12
XFILLER_15_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _23_/HI mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/TEB
+ mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_150 vgnd vpwr scs8hd_decap_3
XFILLER_31_153 vpwr vgnd scs8hd_fill_2
XFILLER_22_120 vgnd vpwr scs8hd_decap_12
XFILLER_9_102 vgnd vpwr scs8hd_decap_4
XFILLER_9_113 vpwr vgnd scs8hd_fill_2
XFILLER_13_153 vgnd vpwr scs8hd_decap_12
XFILLER_13_197 vgnd vpwr scs8hd_decap_4
XFILLER_3_10 vgnd vpwr scs8hd_decap_8
XFILLER_12_63 vgnd vpwr scs8hd_fill_1
XFILLER_12_96 vgnd vpwr scs8hd_decap_12
XFILLER_18_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_204 vgnd vpwr scs8hd_decap_8
XFILLER_24_215 vgnd vpwr scs8hd_decap_3
XFILLER_3_119 vgnd vpwr scs8hd_decap_3
XFILLER_3_108 vpwr vgnd scs8hd_fill_2
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_8
XFILLER_2_163 vgnd vpwr scs8hd_decap_8
XFILLER_2_130 vgnd vpwr scs8hd_decap_4
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_29 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/TEB mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_19 vgnd vpwr scs8hd_decap_12
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_29_83 vpwr vgnd scs8hd_fill_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_4
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_34_162 vpwr vgnd scs8hd_fill_2
XFILLER_34_173 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vgnd vpwr scs8hd_decap_4
XFILLER_25_184 vgnd vpwr scs8hd_decap_8
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/TEB mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_162 vgnd vpwr scs8hd_decap_3
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_132 vgnd vpwr scs8hd_decap_4
XFILLER_22_154 vgnd vpwr scs8hd_decap_8
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XFILLER_9_169 vgnd vpwr scs8hd_decap_12
XFILLER_13_165 vgnd vpwr scs8hd_fill_1
XFILLER_3_22 vgnd vpwr scs8hd_decap_4
XFILLER_3_77 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/TEB mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_106 vgnd vpwr scs8hd_decap_8
XFILLER_10_102 vgnd vpwr scs8hd_decap_8
XFILLER_10_113 vgnd vpwr scs8hd_decap_12
XFILLER_10_157 vgnd vpwr scs8hd_decap_8
XFILLER_10_168 vpwr vgnd scs8hd_fill_2
XFILLER_12_20 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_208 vgnd vpwr scs8hd_decap_6
XFILLER_23_74 vgnd vpwr scs8hd_decap_6
XFILLER_0_12 vpwr vgnd scs8hd_fill_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_78 vgnd vpwr scs8hd_decap_12
XFILLER_9_10 vpwr vgnd scs8hd_fill_2
XFILLER_9_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_84 vgnd vpwr scs8hd_decap_8
XFILLER_4_215 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_160 vgnd vpwr scs8hd_decap_12
XFILLER_34_185 vgnd vpwr scs8hd_fill_1
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_16_174 vgnd vpwr scs8hd_decap_8
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_199 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _17_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

