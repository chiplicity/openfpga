* NGSPICE file created from sb_0__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt sb_0__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_out[0]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_11_
+ top_left_grid_pin_13_ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_
+ top_left_grid_pin_5_ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_
+ vpwr vgnd
XFILLER_39_266 vgnd vpwr scs8hd_decap_8
XFILLER_39_211 vgnd vpwr scs8hd_decap_12
Xmem_right_track_12.LATCH_1_.latch data_in _115_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_166 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
XFILLER_26_85 vgnd vpwr scs8hd_decap_4
XFILLER_3_34 vgnd vpwr scs8hd_decap_12
XFILLER_36_258 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_107 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_76 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _115_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_8
XFILLER_5_173 vgnd vpwr scs8hd_decap_8
XANTENNA__124__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_4
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
X_131_ _153_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_8
XFILLER_2_132 vgnd vpwr scs8hd_decap_12
XFILLER_9_22 vgnd vpwr scs8hd_decap_4
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_20 vgnd vpwr scs8hd_decap_8
XFILLER_18_64 vgnd vpwr scs8hd_fill_1
XFILLER_18_75 vpwr vgnd scs8hd_fill_2
XFILLER_18_97 vgnd vpwr scs8hd_fill_1
XFILLER_34_85 vgnd vpwr scs8hd_decap_6
XFILLER_34_52 vpwr vgnd scs8hd_fill_2
XFILLER_7_213 vgnd vpwr scs8hd_decap_12
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
X_114_ _114_/A _114_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XANTENNA__121__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _182_/HI _119_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _187_/HI _086_/Y mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_106 vpwr vgnd scs8hd_fill_2
XFILLER_4_238 vgnd vpwr scs8hd_decap_12
XFILLER_4_227 vgnd vpwr scs8hd_decap_8
XFILLER_20_32 vgnd vpwr scs8hd_decap_8
XFILLER_20_87 vgnd vpwr scs8hd_decap_4
XFILLER_6_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_6
XFILLER_19_172 vgnd vpwr scs8hd_decap_8
Xmem_right_track_8.LATCH_1_.latch data_in _111_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_145 vgnd vpwr scs8hd_decap_8
XFILLER_31_31 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _110_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_0_274 vgnd vpwr scs8hd_decap_3
XFILLER_16_186 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _114_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_223 vgnd vpwr scs8hd_decap_12
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XFILLER_22_112 vgnd vpwr scs8hd_decap_4
Xmem_top_track_4.LATCH_0_.latch data_in _090_/A _132_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_167 vgnd vpwr scs8hd_decap_6
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XFILLER_26_75 vgnd vpwr scs8hd_decap_4
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_127 vgnd vpwr scs8hd_fill_1
XFILLER_3_46 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_99 vgnd vpwr scs8hd_fill_1
XFILLER_37_96 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XFILLER_26_270 vgnd vpwr scs8hd_decap_4
XFILLER_5_152 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_4
Xmux_top_track_6.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
X_130_ address[3] _133_/B _133_/C _175_/A _131_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_144 vgnd vpwr scs8hd_decap_8
XANTENNA__135__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_34_97 vgnd vpwr scs8hd_decap_4
XFILLER_34_64 vpwr vgnd scs8hd_fill_2
XFILLER_7_225 vgnd vpwr scs8hd_decap_12
XFILLER_11_232 vgnd vpwr scs8hd_decap_8
X_113_ _113_/A _113_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _116_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_6.tap_buf4_0_.scs8hd_inv_1 mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _210_/A vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _118_/A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_184 vgnd vpwr scs8hd_fill_1
XFILLER_1_90 vgnd vpwr scs8hd_decap_3
XFILLER_20_99 vgnd vpwr scs8hd_decap_4
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _102_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_25_165 vgnd vpwr scs8hd_decap_12
XFILLER_15_99 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_31_179 vgnd vpwr scs8hd_decap_4
XFILLER_31_168 vgnd vpwr scs8hd_decap_4
XFILLER_31_113 vgnd vpwr scs8hd_decap_3
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_198 vgnd vpwr scs8hd_decap_12
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__127__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__143__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_235 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _105_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _088_/Y mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_32 vgnd vpwr scs8hd_fill_1
XFILLER_13_102 vgnd vpwr scs8hd_fill_1
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_3_58 vgnd vpwr scs8hd_decap_3
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_8_150 vgnd vpwr scs8hd_decap_3
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_75 vpwr vgnd scs8hd_fill_2
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_6 vgnd vpwr scs8hd_decap_3
XANTENNA__140__B _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_274 vgnd vpwr scs8hd_fill_1
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_11 vpwr vgnd scs8hd_fill_2
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_79 vgnd vpwr scs8hd_decap_4
XFILLER_36_3 vgnd vpwr scs8hd_decap_6
XANTENNA__151__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _088_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_8
XFILLER_34_21 vgnd vpwr scs8hd_decap_8
XFILLER_7_237 vgnd vpwr scs8hd_decap_4
X_112_ _112_/A _112_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_4.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_152 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _107_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _105_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_20_45 vpwr vgnd scs8hd_fill_2
XFILLER_20_56 vpwr vgnd scs8hd_fill_2
XFILLER_20_78 vgnd vpwr scs8hd_decap_6
XFILLER_29_76 vgnd vpwr scs8hd_decap_3
XFILLER_28_163 vgnd vpwr scs8hd_decap_8
XFILLER_20_6 vgnd vpwr scs8hd_decap_6
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_25_177 vgnd vpwr scs8hd_decap_6
XFILLER_40_169 vgnd vpwr scs8hd_decap_12
XFILLER_31_99 vpwr vgnd scs8hd_fill_2
XFILLER_31_88 vpwr vgnd scs8hd_fill_2
XFILLER_31_44 vpwr vgnd scs8hd_fill_2
XFILLER_16_133 vgnd vpwr scs8hd_fill_1
XFILLER_31_103 vgnd vpwr scs8hd_fill_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _133_/C vgnd vpwr scs8hd_diode_2
XANTENNA__143__B _143_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _107_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_11 vgnd vpwr scs8hd_fill_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _185_/HI _109_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _090_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_68 vgnd vpwr scs8hd_fill_1
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_0_.latch data_in _085_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_fill_1
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_168 vgnd vpwr scs8hd_decap_12
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_3 vgnd vpwr scs8hd_fill_1
XANTENNA__151__B _150_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _113_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_8
XFILLER_18_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
X_111_ _111_/A _111_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XANTENNA__146__B _146_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_11 vgnd vpwr scs8hd_decap_4
XFILLER_29_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_101 vgnd vpwr scs8hd_fill_1
XANTENNA__157__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _181_/HI _117_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_104 vgnd vpwr scs8hd_fill_1
XFILLER_31_56 vpwr vgnd scs8hd_fill_2
XFILLER_31_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_123 vpwr vgnd scs8hd_fill_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_8
XFILLER_16_167 vgnd vpwr scs8hd_decap_4
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _133_/D vgnd vpwr scs8hd_diode_2
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XFILLER_38_270 vgnd vpwr scs8hd_decap_4
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_26_89 vgnd vpwr scs8hd_fill_1
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B _153_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_130 vgnd vpwr scs8hd_decap_3
XFILLER_8_163 vgnd vpwr scs8hd_decap_12
XFILLER_12_170 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _108_/A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__170__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_107 vgnd vpwr scs8hd_decap_4
XANTENNA__080__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_33 vpwr vgnd scs8hd_fill_2
XFILLER_37_22 vgnd vpwr scs8hd_decap_4
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_4
XFILLER_5_188 vgnd vpwr scs8hd_fill_1
XANTENNA__149__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_37 vgnd vpwr scs8hd_decap_12
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _112_/Y mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_79 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _110_/Y vgnd vpwr scs8hd_inv_8
XFILLER_34_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _113_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_121 vgnd vpwr scs8hd_fill_1
XFILLER_1_82 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_34 vgnd vpwr scs8hd_decap_8
XFILLER_28_143 vgnd vpwr scs8hd_decap_8
XFILLER_6_16 vgnd vpwr scs8hd_decap_12
XFILLER_3_253 vpwr vgnd scs8hd_fill_2
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_34_113 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_25_157 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A enable vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _116_/A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vpwr vgnd scs8hd_fill_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _153_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_8_142 vgnd vpwr scs8hd_decap_8
XFILLER_8_175 vgnd vpwr scs8hd_decap_12
XFILLER_12_182 vgnd vpwr scs8hd_decap_12
XANTENNA__170__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_0.LATCH_1_.latch data_in _103_/A _153_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _120_/Y mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_8.LATCH_1_.latch data_in _093_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _115_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _085_/Y mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_32_211 vgnd vpwr scs8hd_decap_3
XANTENNA__149__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_6 vpwr vgnd scs8hd_fill_2
XFILLER_14_200 vgnd vpwr scs8hd_decap_12
XFILLER_9_49 vgnd vpwr scs8hd_decap_6
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _108_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A _133_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _101_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_68 vpwr vgnd scs8hd_fill_2
XFILLER_11_258 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_169_ address[0] _169_/B _169_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_3 vpwr vgnd scs8hd_fill_2
XFILLER_37_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_28_122 vpwr vgnd scs8hd_fill_2
XFILLER_6_28 vgnd vpwr scs8hd_decap_3
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_100 vgnd vpwr scs8hd_decap_3
XFILLER_19_111 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_125 vgnd vpwr scs8hd_decap_4
XANTENNA__173__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_25_136 vpwr vgnd scs8hd_fill_2
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_180 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _103_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_60 vgnd vpwr scs8hd_fill_1
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_58 vgnd vpwr scs8hd_decap_4
Xmem_top_track_14.LATCH_0_.latch data_in _100_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_150 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _110_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_194 vgnd vpwr scs8hd_decap_12
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_187 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _152_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _087_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _198_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_79 vpwr vgnd scs8hd_fill_2
XFILLER_37_46 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_209 vgnd vpwr scs8hd_decap_4
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XANTENNA__149__D _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_17_253 vpwr vgnd scs8hd_fill_2
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _184_/HI _107_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_15 vpwr vgnd scs8hd_fill_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_182 vgnd vpwr scs8hd_fill_1
XANTENNA__176__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_260 vpwr vgnd scs8hd_fill_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_3
X_168_ _153_/A _169_/B _168_/Y vgnd vpwr scs8hd_nor2_4
X_099_ _099_/A _099_/Y vgnd vpwr scs8hd_inv_8
XFILLER_27_3 vgnd vpwr scs8hd_decap_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_3
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_95 vgnd vpwr scs8hd_decap_12
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_49 vgnd vpwr scs8hd_decap_4
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_211 vgnd vpwr scs8hd_decap_12
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_148 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _089_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__173__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_31_48 vpwr vgnd scs8hd_fill_2
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_192 vgnd vpwr scs8hd_decap_12
XFILLER_21_81 vpwr vgnd scs8hd_fill_2
XFILLER_39_207 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_15_170 vpwr vgnd scs8hd_fill_2
XFILLER_22_129 vgnd vpwr scs8hd_decap_12
XFILLER_7_72 vgnd vpwr scs8hd_decap_3
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XFILLER_26_37 vpwr vgnd scs8hd_fill_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_162 vgnd vpwr scs8hd_decap_6
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _115_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_12_140 vgnd vpwr scs8hd_decap_4
XFILLER_8_199 vgnd vpwr scs8hd_decap_12
XANTENNA__170__D _133_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_169 vpwr vgnd scs8hd_fill_2
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _106_/A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_4.LATCH_1_.latch data_in _089_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA__176__C _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_81 vpwr vgnd scs8hd_fill_2
XFILLER_40_80 vgnd vpwr scs8hd_fill_1
X_098_ _098_/A _098_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
X_167_ _145_/A _133_/B _152_/C _175_/A _169_/B vgnd vpwr scs8hd_or4_4
XFILLER_37_113 vgnd vpwr scs8hd_decap_8
XFILLER_37_157 vgnd vpwr scs8hd_decap_3
XFILLER_37_135 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_6
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _110_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_8
XFILLER_3_223 vgnd vpwr scs8hd_decap_12
XFILLER_10_83 vgnd vpwr scs8hd_decap_8
XANTENNA__173__D _173_/D vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_160 vpwr vgnd scs8hd_fill_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_127 vgnd vpwr scs8hd_decap_6
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_71 vgnd vpwr scs8hd_decap_3
XFILLER_11_7 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_182 vgnd vpwr scs8hd_fill_1
XFILLER_22_108 vpwr vgnd scs8hd_fill_2
XFILLER_7_95 vgnd vpwr scs8hd_decap_4
XFILLER_7_62 vgnd vpwr scs8hd_fill_1
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _116_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _114_/A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_26_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmem_top_track_10.LATCH_0_.latch data_in _096_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_258 vgnd vpwr scs8hd_decap_12
XFILLER_27_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _212_/A vgnd vpwr scs8hd_inv_1
XFILLER_13_94 vpwr vgnd scs8hd_fill_2
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _118_/Y mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_28 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_210 vgnd vpwr scs8hd_decap_4
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
X_097_ _097_/A _097_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ address[0] _164_/X _166_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_169 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _118_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_73 vgnd vpwr scs8hd_decap_4
XFILLER_19_82 vpwr vgnd scs8hd_fill_2
XFILLER_19_136 vgnd vpwr scs8hd_decap_12
XFILLER_34_117 vgnd vpwr scs8hd_decap_6
X_149_ address[3] address[2] _152_/C _175_/A _150_/B vgnd vpwr scs8hd_or4_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_4
XFILLER_40_109 vgnd vpwr scs8hd_decap_12
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_106 vpwr vgnd scs8hd_fill_2
XFILLER_24_150 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_94 vgnd vpwr scs8hd_decap_3
XFILLER_30_164 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_175 vgnd vpwr scs8hd_decap_12
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_120 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_6
XFILLER_32_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _107_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_8
XFILLER_27_71 vpwr vgnd scs8hd_fill_2
XFILLER_40_270 vgnd vpwr scs8hd_decap_4
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XFILLER_4_182 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_108 vgnd vpwr scs8hd_decap_12
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_14_259 vgnd vpwr scs8hd_decap_12
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_163 vgnd vpwr scs8hd_fill_1
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_241 vgnd vpwr scs8hd_decap_3
XFILLER_34_17 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _183_/HI _105_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _090_/Y vgnd vpwr
+ scs8hd_diode_2
X_165_ _153_/A _164_/X _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_3
XFILLER_34_7 vgnd vpwr scs8hd_fill_1
XFILLER_6_255 vgnd vpwr scs8hd_decap_12
X_096_ _096_/A _096_/Y vgnd vpwr scs8hd_inv_8
Xmem_top_track_0.LATCH_1_.latch data_in _086_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_104 vpwr vgnd scs8hd_fill_2
XFILLER_28_126 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _109_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_115 vgnd vpwr scs8hd_decap_4
XFILLER_19_148 vgnd vpwr scs8hd_decap_12
XFILLER_35_71 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_181 vpwr vgnd scs8hd_fill_2
X_148_ address[4] _173_/D _152_/C vgnd vpwr scs8hd_nand2_4
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XFILLER_30_187 vgnd vpwr scs8hd_decap_12
XFILLER_30_154 vgnd vpwr scs8hd_fill_1
XFILLER_30_143 vgnd vpwr scs8hd_decap_8
XFILLER_30_110 vgnd vpwr scs8hd_decap_4
XFILLER_7_20 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _096_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XFILLER_32_50 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _092_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_139 vpwr vgnd scs8hd_fill_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _179_/HI _113_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_194 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
Xmem_right_track_14.LATCH_0_.latch data_in _118_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_264 vpwr vgnd scs8hd_fill_2
XFILLER_34_29 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _104_/A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_24_51 vpwr vgnd scs8hd_fill_2
XFILLER_6_245 vgnd vpwr scs8hd_fill_1
XFILLER_6_267 vgnd vpwr scs8hd_decap_8
X_164_ _145_/A address[2] _152_/C _133_/D _164_/X vgnd vpwr scs8hd_or4_4
X_095_ _095_/A _095_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_29 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_237 vgnd vpwr scs8hd_decap_6
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XFILLER_19_105 vgnd vpwr scs8hd_decap_3
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_147_ address[0] _146_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_152 vpwr vgnd scs8hd_fill_2
XFILLER_25_108 vgnd vpwr scs8hd_decap_4
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_16_119 vpwr vgnd scs8hd_fill_2
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _101_/A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_199 vgnd vpwr scs8hd_decap_12
XFILLER_15_174 vgnd vpwr scs8hd_decap_8
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _108_/Y mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_12.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_144 vgnd vpwr scs8hd_fill_1
XFILLER_32_84 vgnd vpwr scs8hd_decap_8
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_29 vpwr vgnd scs8hd_fill_2
XFILLER_37_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_258 vgnd vpwr scs8hd_decap_12
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_4
XFILLER_27_95 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_162 vgnd vpwr scs8hd_decap_12
XFILLER_4_88 vgnd vpwr scs8hd_decap_4
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_86 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_50 vgnd vpwr scs8hd_decap_12
XFILLER_1_198 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_6
XFILLER_9_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_85 vgnd vpwr scs8hd_decap_4
XFILLER_40_84 vgnd vpwr scs8hd_decap_8
X_163_ address[0] _163_/B _163_/Y vgnd vpwr scs8hd_nor2_4
X_094_ _094_/A _094_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_242 vgnd vpwr scs8hd_decap_8
XFILLER_37_139 vpwr vgnd scs8hd_fill_2
XFILLER_28_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _115_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _116_/Y mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__212__A _212_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_35_40 vgnd vpwr scs8hd_fill_1
XFILLER_19_52 vgnd vpwr scs8hd_fill_1
XFILLER_35_84 vpwr vgnd scs8hd_fill_2
X_146_ _153_/A _146_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_33_131 vpwr vgnd scs8hd_fill_2
XFILLER_18_161 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_153 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_77 vgnd vpwr scs8hd_decap_3
X_129_ address[0] _128_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_7_182 vgnd vpwr scs8hd_fill_1
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_30 vpwr vgnd scs8hd_fill_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_4
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XFILLER_4_174 vgnd vpwr scs8hd_decap_8
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_31_240 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _117_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XFILLER_13_98 vgnd vpwr scs8hd_decap_4
XFILLER_1_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_3
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
XFILLER_38_62 vgnd vpwr scs8hd_decap_12
Xmem_top_track_14.LATCH_1_.latch data_in _099_/A _146_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _110_/Y vgnd vpwr
+ scs8hd_diode_2
X_162_ _153_/A _163_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_64 vpwr vgnd scs8hd_fill_2
XFILLER_24_97 vpwr vgnd scs8hd_fill_2
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
X_093_ _093_/A _093_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_9 vpwr vgnd scs8hd_fill_2
Xmem_right_track_10.LATCH_0_.latch data_in _114_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_35_52 vpwr vgnd scs8hd_fill_2
XFILLER_19_86 vgnd vpwr scs8hd_decap_3
XFILLER_27_162 vpwr vgnd scs8hd_fill_2
XFILLER_27_173 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _178_/HI _103_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _145_/A _133_/B _133_/C _133_/D _146_/B vgnd vpwr scs8hd_or4_4
XFILLER_32_7 vgnd vpwr scs8hd_fill_1
XANTENNA__122__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
XFILLER_18_173 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_132 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_32 vpwr vgnd scs8hd_fill_2
XFILLER_21_76 vgnd vpwr scs8hd_decap_3
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
X_128_ _153_/A _128_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_168 vgnd vpwr scs8hd_decap_4
XFILLER_7_56 vpwr vgnd scs8hd_fill_2
XFILLER_7_12 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.tap_buf4_0_.scs8hd_inv_1 mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _208_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_168 vgnd vpwr scs8hd_fill_1
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_12_124 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _112_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _089_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_75 vpwr vgnd scs8hd_fill_2
XFILLER_40_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA__130__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_11 vgnd vpwr scs8hd_decap_12
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_178 vgnd vpwr scs8hd_decap_4
XFILLER_38_96 vgnd vpwr scs8hd_decap_12
XFILLER_38_74 vgnd vpwr scs8hd_fill_1
Xmem_right_track_6.LATCH_0_.latch data_in _110_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_4
XANTENNA__141__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_182 vgnd vpwr scs8hd_fill_1
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_161_ _145_/A address[2] _152_/C _175_/A _163_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_32 vgnd vpwr scs8hd_decap_6
X_092_ _092_/A _092_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__136__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_163 vgnd vpwr scs8hd_decap_12
XFILLER_28_108 vgnd vpwr scs8hd_decap_3
XFILLER_10_56 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _095_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_119 vgnd vpwr scs8hd_fill_1
XFILLER_35_97 vpwr vgnd scs8hd_fill_2
XFILLER_35_20 vpwr vgnd scs8hd_fill_2
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ address[0] _143_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _213_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_33_100 vpwr vgnd scs8hd_fill_2
XFILLER_18_141 vpwr vgnd scs8hd_fill_2
XFILLER_18_185 vgnd vpwr scs8hd_decap_12
XFILLER_33_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _091_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_11 vpwr vgnd scs8hd_fill_2
XFILLER_21_99 vgnd vpwr scs8hd_decap_3
XFILLER_30_125 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_7_24 vgnd vpwr scs8hd_decap_12
X_127_ address[3] address[2] _133_/C _133_/D _128_/B vgnd vpwr scs8hd_or4_4
XANTENNA__133__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_32_21 vpwr vgnd scs8hd_fill_2
XFILLER_32_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_107 vpwr vgnd scs8hd_fill_2
XFILLER_8_118 vgnd vpwr scs8hd_decap_12
XFILLER_12_103 vpwr vgnd scs8hd_fill_2
XFILLER_12_147 vgnd vpwr scs8hd_decap_6
XFILLER_12_158 vgnd vpwr scs8hd_decap_12
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_3
XANTENNA__128__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_decap_3
XANTENNA__144__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_162 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _099_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _106_/Y mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_4_198 vgnd vpwr scs8hd_decap_12
XANTENNA__130__C _133_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_23 vgnd vpwr scs8hd_decap_12
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_268 vgnd vpwr scs8hd_decap_8
XANTENNA__141__B _139_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_172 vpwr vgnd scs8hd_fill_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_091_ _091_/A _091_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_10_201 vgnd vpwr scs8hd_decap_12
X_160_ address[0] _160_/B _160_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_98 vgnd vpwr scs8hd_decap_6
XFILLER_40_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_109 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_271 vgnd vpwr scs8hd_decap_6
XANTENNA__152__A address[3] vgnd vpwr scs8hd_diode_2
Xmem_top_track_10.LATCH_1_.latch data_in _095_/A _140_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_175 vgnd vpwr scs8hd_decap_12
XFILLER_10_79 vpwr vgnd scs8hd_fill_2
XFILLER_19_44 vgnd vpwr scs8hd_decap_8
XFILLER_19_55 vgnd vpwr scs8hd_decap_4
XFILLER_19_66 vgnd vpwr scs8hd_fill_1
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
X_212_ _212_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_35_32 vpwr vgnd scs8hd_fill_2
X_143_ _153_/A _143_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_7 vgnd vpwr scs8hd_decap_8
XFILLER_18_197 vgnd vpwr scs8hd_decap_12
XFILLER_33_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__147__A address[0] vgnd vpwr scs8hd_diode_2
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_101 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _114_/Y mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_7_36 vgnd vpwr scs8hd_decap_12
XANTENNA__133__C _133_/C vgnd vpwr scs8hd_diode_2
X_126_ address[1] enable _133_/D vgnd vpwr scs8hd_nand2_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_21_115 vpwr vgnd scs8hd_fill_2
XFILLER_21_126 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _118_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _143_/B vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _109_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__160__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_22 vpwr vgnd scs8hd_fill_2
XFILLER_27_88 vgnd vpwr scs8hd_decap_4
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_122 vgnd vpwr scs8hd_fill_1
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA__130__D _175_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_13_35 vgnd vpwr scs8hd_decap_12
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_4
XFILLER_38_21 vgnd vpwr scs8hd_decap_8
XFILLER_13_232 vgnd vpwr scs8hd_decap_8
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XFILLER_13_265 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_39_162 vgnd vpwr scs8hd_decap_4
XFILLER_39_151 vgnd vpwr scs8hd_decap_4
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
X_090_ _090_/A _090_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_239 vgnd vpwr scs8hd_decap_6
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_24_89 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _102_/A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA__136__C _133_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__152__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_187 vgnd vpwr scs8hd_decap_12
XFILLER_36_121 vgnd vpwr scs8hd_decap_4
Xmem_right_track_2.LATCH_0_.latch data_in _106_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_12 vpwr vgnd scs8hd_fill_2
XFILLER_19_78 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_88 vgnd vpwr scs8hd_decap_4
XFILLER_35_66 vgnd vpwr scs8hd_decap_3
X_211_ _211_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_142_ _145_/A _133_/B _133_/C _175_/A _143_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _120_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_146 vgnd vpwr scs8hd_decap_4
XFILLER_33_113 vgnd vpwr scs8hd_decap_8
XFILLER_18_154 vgnd vpwr scs8hd_decap_4
XANTENNA__147__B _146_/B vgnd vpwr scs8hd_diode_2
XANTENNA__163__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_157 vgnd vpwr scs8hd_decap_8
XFILLER_24_168 vgnd vpwr scs8hd_decap_12
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_157 vpwr vgnd scs8hd_fill_2
X_125_ address[0] _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_138 vgnd vpwr scs8hd_decap_3
XFILLER_7_48 vgnd vpwr scs8hd_decap_6
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__133__D _133_/D vgnd vpwr scs8hd_diode_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_21_138 vgnd vpwr scs8hd_decap_12
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_67 vpwr vgnd scs8hd_fill_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_7_142 vgnd vpwr scs8hd_decap_3
X_108_ _108_/A _108_/Y vgnd vpwr scs8hd_inv_8
XFILLER_21_3 vgnd vpwr scs8hd_decap_3
XANTENNA__160__B _160_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _109_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_4_145 vgnd vpwr scs8hd_decap_8
XFILLER_4_134 vgnd vpwr scs8hd_decap_8
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XANTENNA__139__C _133_/C vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__155__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_47 vgnd vpwr scs8hd_decap_12
XFILLER_38_11 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_4
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__166__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _096_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_70 vgnd vpwr scs8hd_fill_1
XFILLER_39_196 vgnd vpwr scs8hd_decap_8
XFILLER_24_68 vpwr vgnd scs8hd_fill_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XANTENNA__136__D _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XANTENNA__152__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_36_111 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _092_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_56 vgnd vpwr scs8hd_decap_3
XFILLER_27_166 vpwr vgnd scs8hd_fill_2
XFILLER_27_177 vpwr vgnd scs8hd_fill_2
X_210_ _210_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_141_ address[0] _139_/X _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _093_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_111 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _117_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _111_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_136 vgnd vpwr scs8hd_decap_12
XFILLER_21_36 vpwr vgnd scs8hd_fill_2
XFILLER_30_117 vgnd vpwr scs8hd_decap_6
XFILLER_30_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_136 vgnd vpwr scs8hd_decap_4
XFILLER_7_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
X_124_ _153_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _175_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_128 vgnd vpwr scs8hd_decap_12
X_107_ _107_/A _107_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _098_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__169__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XFILLER_4_157 vgnd vpwr scs8hd_decap_3
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XANTENNA__139__D _133_/D vgnd vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _094_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__155__C _152_/C vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _170_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _097_/A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _104_/Y mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_9_238 vgnd vpwr scs8hd_fill_1
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_260 vgnd vpwr scs8hd_decap_4
XFILLER_5_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_8
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XANTENNA__152__D _133_/D vgnd vpwr scs8hd_diode_2
XFILLER_36_145 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _133_/D vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_24 vpwr vgnd scs8hd_fill_2
XFILLER_27_145 vpwr vgnd scs8hd_fill_2
X_140_ _153_/A _139_/X _140_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_200 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _101_/Y mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_33_126 vgnd vpwr scs8hd_decap_3
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_115 vpwr vgnd scs8hd_fill_2
XFILLER_21_15 vpwr vgnd scs8hd_fill_2
Xmem_top_track_6.LATCH_0_.latch data_in _092_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_123_ address[3] address[2] _133_/C _175_/A _125_/B vgnd vpwr scs8hd_or4_4
XANTENNA__158__C _152_/C vgnd vpwr scs8hd_diode_2
XANTENNA__174__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_240 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_107 vgnd vpwr scs8hd_decap_4
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_25 vgnd vpwr scs8hd_decap_6
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XFILLER_7_166 vgnd vpwr scs8hd_decap_12
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
X_106_ _106_/A _106_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
XANTENNA__169__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_71 vpwr vgnd scs8hd_fill_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_232 vgnd vpwr scs8hd_decap_12
XFILLER_27_47 vpwr vgnd scs8hd_fill_2
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_91 vgnd vpwr scs8hd_decap_3
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__155__D _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_5_50 vgnd vpwr scs8hd_decap_8
XFILLER_39_176 vgnd vpwr scs8hd_decap_6
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_36_102 vgnd vpwr scs8hd_decap_3
XANTENNA__177__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_35_36 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _117_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_212 vpwr vgnd scs8hd_fill_2
XFILLER_18_124 vgnd vpwr scs8hd_decap_3
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _100_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_199_ _199_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_84 vgnd vpwr scs8hd_decap_8
XFILLER_24_105 vgnd vpwr scs8hd_fill_1
XFILLER_32_182 vgnd vpwr scs8hd_decap_8
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
X_122_ address[1] _122_/B _175_/A vgnd vpwr scs8hd_or2_4
XFILLER_11_71 vgnd vpwr scs8hd_decap_4
XANTENNA__158__D _133_/D vgnd vpwr scs8hd_diode_2
XFILLER_21_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__C _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_32_37 vgnd vpwr scs8hd_decap_4
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
Xmem_right_track_10.LATCH_1_.latch data_in _113_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_7_101 vpwr vgnd scs8hd_fill_2
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
X_105_ _105_/A _105_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_70 vgnd vpwr scs8hd_decap_4
XFILLER_7_178 vgnd vpwr scs8hd_decap_4
XFILLER_7_189 vgnd vpwr scs8hd_decap_12
XFILLER_27_26 vpwr vgnd scs8hd_fill_2
XFILLER_40_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_70 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_107 vgnd vpwr scs8hd_decap_12
XFILLER_38_36 vgnd vpwr scs8hd_fill_1
XFILLER_13_258 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _119_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_140 vgnd vpwr scs8hd_fill_1
XFILLER_0_184 vpwr vgnd scs8hd_fill_2
XFILLER_5_73 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_8
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_70 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _112_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_125 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__177__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_16 vpwr vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_18_158 vgnd vpwr scs8hd_fill_1
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_96 vgnd vpwr scs8hd_decap_12
XFILLER_17_180 vgnd vpwr scs8hd_decap_3
Xmem_right_track_6.LATCH_1_.latch data_in _109_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_121_ address[4] address[5] _133_/C vgnd vpwr scs8hd_or2_4
Xmux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _091_/A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
X_104_ _104_/A _104_/Y vgnd vpwr scs8hd_inv_8
Xmem_top_track_2.LATCH_0_.latch data_in _088_/A _129_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_34_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _095_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_204 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _091_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_92 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_119 vgnd vpwr scs8hd_decap_3
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_30_93 vgnd vpwr scs8hd_decap_4
XFILLER_5_200 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _095_/A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_91 vgnd vpwr scs8hd_decap_3
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_19_39 vgnd vpwr scs8hd_decap_3
XFILLER_27_115 vpwr vgnd scs8hd_fill_2
XFILLER_27_126 vgnd vpwr scs8hd_decap_4
XFILLER_35_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _197_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _104_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
X_197_ _197_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _097_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_93 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
X_120_ _120_/A _120_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_3
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _093_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _099_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_154 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _103_/A _103_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_158 vpwr vgnd scs8hd_fill_2
XFILLER_22_83 vpwr vgnd scs8hd_fill_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_40_205 vgnd vpwr scs8hd_decap_8
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_106 vgnd vpwr scs8hd_decap_12
XFILLER_17_50 vgnd vpwr scs8hd_decap_8
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_216 vgnd vpwr scs8hd_decap_12
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _094_/A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_164 vgnd vpwr scs8hd_decap_12
XFILLER_28_82 vpwr vgnd scs8hd_fill_2
XFILLER_28_71 vgnd vpwr scs8hd_decap_3
XFILLER_12_260 vgnd vpwr scs8hd_decap_12
XFILLER_5_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_168 vgnd vpwr scs8hd_fill_1
XFILLER_39_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _200_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_83 vgnd vpwr scs8hd_decap_8
XFILLER_5_245 vgnd vpwr scs8hd_decap_3
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_149 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_119 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vpwr vgnd scs8hd_fill_2
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _098_/A mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _105_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
X_102_ _102_/A _102_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_51 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _120_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_118 vgnd vpwr scs8hd_decap_4
XFILLER_17_62 vgnd vpwr scs8hd_decap_8
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_228 vgnd vpwr scs8hd_decap_12
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_195 vpwr vgnd scs8hd_fill_2
XFILLER_3_184 vpwr vgnd scs8hd_fill_2
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
XFILLER_38_39 vpwr vgnd scs8hd_fill_2
XFILLER_38_17 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _102_/Y mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_110 vgnd vpwr scs8hd_decap_12
XFILLER_0_132 vgnd vpwr scs8hd_decap_8
XFILLER_0_154 vgnd vpwr scs8hd_fill_1
XFILLER_0_176 vgnd vpwr scs8hd_decap_8
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_12_272 vgnd vpwr scs8hd_decap_3
XFILLER_39_158 vpwr vgnd scs8hd_fill_2
XFILLER_39_147 vpwr vgnd scs8hd_fill_2
XFILLER_40_18 vgnd vpwr scs8hd_decap_12
XFILLER_39_60 vgnd vpwr scs8hd_fill_1
XFILLER_36_128 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_26_150 vgnd vpwr scs8hd_decap_3
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in _102_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_164 vgnd vpwr scs8hd_fill_1
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XFILLER_36_72 vgnd vpwr scs8hd_fill_1
Xmux_top_track_4.tap_buf4_0_.scs8hd_inv_1 mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _211_/A vgnd vpwr scs8hd_inv_1
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_112 vgnd vpwr scs8hd_decap_4
XFILLER_20_123 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_212 vpwr vgnd scs8hd_fill_2
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
X_101_ _101_/A _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_123 vgnd vpwr scs8hd_decap_3
XFILLER_11_156 vgnd vpwr scs8hd_decap_12
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_204 vgnd vpwr scs8hd_decap_8
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _089_/A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__210__A _210_/A vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _111_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_74 vgnd vpwr scs8hd_decap_6
XFILLER_17_96 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_38_29 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_122 vpwr vgnd scs8hd_fill_2
XFILLER_0_144 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_40 vgnd vpwr scs8hd_fill_1
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_8_211 vgnd vpwr scs8hd_decap_3
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_77 vgnd vpwr scs8hd_decap_3
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _098_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_41 vgnd vpwr scs8hd_decap_3
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _093_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_107 vgnd vpwr scs8hd_decap_4
XFILLER_29_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _094_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_107 vpwr vgnd scs8hd_fill_2
XFILLER_18_129 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_52 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_165 vgnd vpwr scs8hd_decap_8
XFILLER_17_140 vpwr vgnd scs8hd_fill_2
XFILLER_17_151 vgnd vpwr scs8hd_decap_6
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_110 vpwr vgnd scs8hd_fill_2
XFILLER_23_132 vgnd vpwr scs8hd_decap_12
XFILLER_11_98 vpwr vgnd scs8hd_fill_2
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_84 vpwr vgnd scs8hd_fill_2
XFILLER_36_62 vgnd vpwr scs8hd_fill_1
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
XFILLER_14_165 vgnd vpwr scs8hd_decap_8
XFILLER_14_176 vgnd vpwr scs8hd_decap_12
X_177_ _133_/D _175_/B address[0] _177_/Y vgnd vpwr scs8hd_nor3_4
Xmux_top_track_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__123__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_135 vgnd vpwr scs8hd_decap_12
XFILLER_9_180 vgnd vpwr scs8hd_decap_3
X_100_ _100_/A _100_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_102 vgnd vpwr scs8hd_decap_4
XFILLER_11_168 vgnd vpwr scs8hd_decap_12
XANTENNA__208__A _208_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _100_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _189_/HI _097_/Y mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_12.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_52 vpwr vgnd scs8hd_fill_2
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_96 vpwr vgnd scs8hd_fill_2
Xmem_top_track_6.LATCH_1_.latch data_in _091_/A _134_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_153 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _103_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_52 vgnd vpwr scs8hd_decap_4
XFILLER_8_256 vpwr vgnd scs8hd_fill_2
XFILLER_8_267 vgnd vpwr scs8hd_decap_8
XFILLER_39_105 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _153_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_259 vgnd vpwr scs8hd_decap_12
XFILLER_5_204 vgnd vpwr scs8hd_decap_12
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _092_/A mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_270 vgnd vpwr scs8hd_decap_4
XFILLER_27_119 vgnd vpwr scs8hd_decap_3
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XFILLER_35_174 vgnd vpwr scs8hd_decap_8
XFILLER_35_163 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_25_31 vpwr vgnd scs8hd_fill_2
XFILLER_26_163 vgnd vpwr scs8hd_decap_12
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XFILLER_25_97 vpwr vgnd scs8hd_fill_2
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_199 vgnd vpwr scs8hd_decap_12
XFILLER_32_133 vpwr vgnd scs8hd_fill_2
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _085_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_144 vgnd vpwr scs8hd_decap_12
XFILLER_11_11 vgnd vpwr scs8hd_decap_12
XFILLER_36_30 vgnd vpwr scs8hd_fill_1
XFILLER_14_188 vgnd vpwr scs8hd_decap_12
X_176_ _133_/D _175_/B _153_/A _176_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_147 vgnd vpwr scs8hd_decap_6
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_4
XFILLER_22_87 vgnd vpwr scs8hd_decap_4
Xmem_top_track_12.LATCH_0_.latch data_in _098_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vpwr vgnd scs8hd_fill_2
XFILLER_8_67 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _153_/A vgnd vpwr scs8hd_diode_2
X_159_ _153_/A _160_/B _159_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_10 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_75 vgnd vpwr scs8hd_decap_4
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _096_/A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_121 vgnd vpwr scs8hd_fill_1
XANTENNA__129__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_209 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_86 vgnd vpwr scs8hd_decap_6
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_54 vgnd vpwr scs8hd_fill_1
XFILLER_5_216 vgnd vpwr scs8hd_decap_12
XFILLER_39_74 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _100_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__B enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_109 vgnd vpwr scs8hd_decap_4
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_10 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_26_142 vgnd vpwr scs8hd_decap_8
XFILLER_26_175 vgnd vpwr scs8hd_decap_12
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_145 vgnd vpwr scs8hd_decap_8
XFILLER_32_112 vgnd vpwr scs8hd_decap_8
XANTENNA__137__A _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _119_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_156 vgnd vpwr scs8hd_decap_8
XFILLER_11_23 vgnd vpwr scs8hd_decap_12
XFILLER_23_167 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_67 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
X_175_ _175_/A _175_/B address[0] _175_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__C _133_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_204 vgnd vpwr scs8hd_decap_12
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XFILLER_28_6 vpwr vgnd scs8hd_fill_2
XFILLER_9_160 vgnd vpwr scs8hd_decap_12
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_28_204 vgnd vpwr scs8hd_decap_8
XFILLER_36_270 vgnd vpwr scs8hd_decap_4
XFILLER_11_115 vpwr vgnd scs8hd_fill_2
XFILLER_11_137 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_11 vgnd vpwr scs8hd_decap_3
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_13 vgnd vpwr scs8hd_decap_12
X_089_ _089_/A _089_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__134__B _135_/B vgnd vpwr scs8hd_diode_2
X_158_ address[3] _133_/B _152_/C _133_/D _160_/B vgnd vpwr scs8hd_or4_4
XANTENNA__150__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_8
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_10 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_199 vgnd vpwr scs8hd_decap_12
XFILLER_3_188 vgnd vpwr scs8hd_decap_4
XANTENNA__129__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
XFILLER_28_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_76 vgnd vpwr scs8hd_decap_3
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _087_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_58 vgnd vpwr scs8hd_decap_3
XFILLER_5_14 vgnd vpwr scs8hd_decap_12
Xmem_top_track_2.LATCH_1_.latch data_in _087_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_162 vpwr vgnd scs8hd_fill_2
XFILLER_30_22 vpwr vgnd scs8hd_fill_2
XFILLER_5_228 vgnd vpwr scs8hd_decap_12
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_39_31 vpwr vgnd scs8hd_fill_2
XFILLER_30_66 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_29_173 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_132 vgnd vpwr scs8hd_decap_4
XFILLER_26_121 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_88 vgnd vpwr scs8hd_decap_3
XFILLER_26_187 vgnd vpwr scs8hd_decap_12
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_242 vpwr vgnd scs8hd_fill_2
XFILLER_17_121 vgnd vpwr scs8hd_fill_1
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XANTENNA__137__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _091_/Y mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_179 vgnd vpwr scs8hd_decap_4
XFILLER_11_35 vgnd vpwr scs8hd_decap_12
XFILLER_36_54 vgnd vpwr scs8hd_decap_8
XFILLER_36_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_124 vpwr vgnd scs8hd_fill_2
XANTENNA__123__D _175_/A vgnd vpwr scs8hd_diode_2
X_174_ _175_/A _175_/B _153_/A _174_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_37_216 vgnd vpwr scs8hd_decap_12
XANTENNA__148__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_8_25 vgnd vpwr scs8hd_decap_6
X_157_ address[0] _157_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_6 vgnd vpwr scs8hd_decap_12
X_088_ _088_/A _088_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__150__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _104_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _097_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_33 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in _120_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_156 vgnd vpwr scs8hd_decap_12
XFILLER_3_123 vpwr vgnd scs8hd_fill_2
XFILLER_30_211 vgnd vpwr scs8hd_decap_3
XFILLER_15_263 vgnd vpwr scs8hd_decap_12
X_209_ _209_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__161__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _093_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_148 vgnd vpwr scs8hd_decap_6
XFILLER_5_26 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _188_/HI _095_/Y mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__156__A _153_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _199_/A vgnd vpwr scs8hd_inv_1
XFILLER_38_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_10 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.tap_buf4_0_.scs8hd_inv_1 mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XFILLER_39_87 vpwr vgnd scs8hd_fill_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XFILLER_29_152 vpwr vgnd scs8hd_fill_2
XANTENNA__142__C _133_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_25_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_199 vgnd vpwr scs8hd_decap_12
XFILLER_1_210 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_100 vpwr vgnd scs8hd_fill_2
XFILLER_17_111 vgnd vpwr scs8hd_decap_4
XANTENNA__153__B _153_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _106_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _090_/A mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _099_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_47 vgnd vpwr scs8hd_decap_12
XFILLER_36_88 vgnd vpwr scs8hd_decap_4
XFILLER_36_66 vgnd vpwr scs8hd_decap_6
X_173_ address[3] address[2] address[4] _173_/D _175_/B vgnd vpwr scs8hd_or4_4
XFILLER_37_228 vgnd vpwr scs8hd_decap_12
XANTENNA__148__B _173_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_087_ _087_/A _087_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_165 vgnd vpwr scs8hd_decap_12
X_156_ _153_/A _157_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XFILLER_6_198 vgnd vpwr scs8hd_decap_12
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _153_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_56 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _094_/Y mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_168 vgnd vpwr scs8hd_decap_12
XFILLER_3_135 vgnd vpwr scs8hd_fill_1
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XFILLER_15_253 vpwr vgnd scs8hd_fill_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
XANTENNA__145__C _133_/C vgnd vpwr scs8hd_diode_2
X_139_ _145_/A address[2] _133_/C _133_/D _139_/X vgnd vpwr scs8hd_or4_4
X_208_ _208_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__161__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_fill_1
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_12_256 vpwr vgnd scs8hd_fill_2
XFILLER_5_38 vgnd vpwr scs8hd_decap_12
XFILLER_39_109 vgnd vpwr scs8hd_decap_12
XANTENNA__172__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _086_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_46 vgnd vpwr scs8hd_decap_8
XANTENNA__082__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XFILLER_4_252 vgnd vpwr scs8hd_decap_3
XANTENNA__142__D _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_101 vpwr vgnd scs8hd_fill_2
XANTENNA__167__A _145_/A vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_35 vpwr vgnd scs8hd_fill_2
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_1_222 vgnd vpwr scs8hd_decap_12
XFILLER_32_137 vgnd vpwr scs8hd_decap_3
XFILLER_40_181 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _098_/Y mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_192 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _111_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_172_ address[0] _170_/X _172_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_130 vpwr vgnd scs8hd_fill_2
XANTENNA__164__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_118 vpwr vgnd scs8hd_fill_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_82 vpwr vgnd scs8hd_fill_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_4
XFILLER_22_47 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_111 vpwr vgnd scs8hd_fill_2
XFILLER_6_177 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
X_155_ address[3] _133_/B _152_/C _175_/A _157_/B vgnd vpwr scs8hd_or4_4
X_086_ _086_/A _086_/Y vgnd vpwr scs8hd_inv_8
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _160_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_14 vgnd vpwr scs8hd_decap_12
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_58 vgnd vpwr scs8hd_decap_3
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_103 vgnd vpwr scs8hd_decap_12
XFILLER_3_147 vgnd vpwr scs8hd_decap_6
Xmem_top_track_16.LATCH_1_.latch data_in _101_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
XANTENNA__145__D _133_/D vgnd vpwr scs8hd_diode_2
X_207_ _207_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_138_ address[0] _138_/B _138_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_180 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_8
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XFILLER_0_106 vpwr vgnd scs8hd_fill_2
XFILLER_0_128 vpwr vgnd scs8hd_fill_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_235 vgnd vpwr scs8hd_fill_1
Xmem_right_track_12.LATCH_0_.latch data_in _116_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__172__B _170_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_fill_1
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_110 vgnd vpwr scs8hd_decap_4
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XFILLER_35_146 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _119_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__167__B _133_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _086_/A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_14 vpwr vgnd scs8hd_fill_2
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_234 vgnd vpwr scs8hd_decap_8
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_168 vgnd vpwr scs8hd_decap_12
XFILLER_40_193 vgnd vpwr scs8hd_decap_12
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vpwr vgnd scs8hd_fill_2
XFILLER_14_149 vgnd vpwr scs8hd_decap_4
X_171_ _153_/A _170_/X _171_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_153 vgnd vpwr scs8hd_fill_1
XANTENNA__164__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_36_274 vgnd vpwr scs8hd_fill_1
XFILLER_11_119 vgnd vpwr scs8hd_decap_3
Xmux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _089_/Y mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_263 vgnd vpwr scs8hd_decap_12
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_130 vpwr vgnd scs8hd_fill_2
XFILLER_10_141 vpwr vgnd scs8hd_fill_2
X_085_ _085_/A _085_/Y vgnd vpwr scs8hd_inv_8
X_154_ address[0] _153_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XANTENNA__175__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_26 vgnd vpwr scs8hd_decap_12
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_25 vgnd vpwr scs8hd_decap_6
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_115 vgnd vpwr scs8hd_decap_6
Xmem_right_track_8.LATCH_0_.latch data_in _112_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
X_137_ _153_/A _138_/B _137_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_192 vgnd vpwr scs8hd_decap_4
XANTENNA__161__D _175_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_36 vgnd vpwr scs8hd_decap_4
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _114_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr scs8hd_diode_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_7_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_38_144 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_26 vgnd vpwr scs8hd_decap_4
XFILLER_39_35 vpwr vgnd scs8hd_fill_2
XFILLER_29_133 vpwr vgnd scs8hd_fill_2
XFILLER_4_210 vgnd vpwr scs8hd_decap_4
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _100_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__167__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_180 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_48 vpwr vgnd scs8hd_fill_2
XFILLER_26_125 vpwr vgnd scs8hd_fill_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_15_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _103_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_106 vpwr vgnd scs8hd_fill_2
XFILLER_31_172 vgnd vpwr scs8hd_fill_1
XFILLER_14_128 vgnd vpwr scs8hd_decap_4
X_170_ _145_/A _133_/B _152_/C _133_/D _170_/X vgnd vpwr scs8hd_or4_4
XFILLER_9_143 vpwr vgnd scs8hd_fill_2
XANTENNA__164__D _133_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_275 vpwr vgnd scs8hd_fill_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
X_153_ _153_/A _153_/B _153_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _088_/A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_102 vgnd vpwr scs8hd_decap_3
X_084_ address[0] _153_/A vgnd vpwr scs8hd_inv_8
XFILLER_12_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_7 vgnd vpwr scs8hd_decap_3
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA__175__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_17_38 vgnd vpwr scs8hd_decap_12
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_37 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_127 vgnd vpwr scs8hd_decap_8
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _085_/Y vgnd vpwr
+ scs8hd_diode_2
X_205_ _205_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _102_/A vgnd vpwr
+ scs8hd_diode_2
X_136_ _145_/A address[2] _133_/C _175_/A _138_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_92 vgnd vpwr scs8hd_fill_1
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_83 vgnd vpwr scs8hd_fill_1
XFILLER_28_59 vgnd vpwr scs8hd_fill_1
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
Xmux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _092_/Y mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _105_/A vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_12.LATCH_1_.latch data_in _097_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_241 vgnd vpwr scs8hd_fill_1
XFILLER_7_274 vgnd vpwr scs8hd_decap_3
X_119_ _119_/A _119_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_14 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_156 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vgnd vpwr scs8hd_fill_1
XFILLER_20_60 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_4
XFILLER_35_159 vpwr vgnd scs8hd_fill_2
XANTENNA__167__D _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_6_73 vpwr vgnd scs8hd_fill_2
XFILLER_6_62 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XFILLER_34_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XFILLER_32_129 vpwr vgnd scs8hd_fill_2
XFILLER_31_92 vgnd vpwr scs8hd_decap_4
XFILLER_31_151 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_6
XFILLER_39_262 vpwr vgnd scs8hd_fill_2
XFILLER_36_37 vgnd vpwr scs8hd_decap_6
XFILLER_22_173 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _088_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_140 vgnd vpwr scs8hd_decap_12
XFILLER_26_81 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_8
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _096_/Y mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_125 vgnd vpwr scs8hd_fill_1
X_083_ enable _122_/B vgnd vpwr scs8hd_inv_8
XFILLER_10_165 vgnd vpwr scs8hd_decap_12
X_152_ address[3] address[2] _152_/C _133_/D _153_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _109_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ address[0] _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_7 vgnd vpwr scs8hd_decap_3
XFILLER_24_6 vgnd vpwr scs8hd_decap_6
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XFILLER_9_95 vgnd vpwr scs8hd_decap_4
XFILLER_12_227 vgnd vpwr scs8hd_decap_8
XFILLER_18_71 vgnd vpwr scs8hd_fill_1
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XFILLER_34_81 vpwr vgnd scs8hd_fill_2
X_118_ _118_/A _118_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_3 vgnd vpwr scs8hd_decap_8
Xmem_right_track_4.LATCH_0_.latch data_in _108_/A _160_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_48 vgnd vpwr scs8hd_decap_12
XFILLER_39_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_92 vgnd vpwr scs8hd_decap_3
XFILLER_35_138 vgnd vpwr scs8hd_decap_6
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_138 vpwr vgnd scs8hd_fill_2
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_60 vgnd vpwr scs8hd_fill_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _117_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_141 vgnd vpwr scs8hd_decap_12
XFILLER_22_185 vgnd vpwr scs8hd_decap_12
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_4
XFILLER_13_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_9_156 vpwr vgnd scs8hd_fill_2
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
XFILLER_6_137 vgnd vpwr scs8hd_decap_6
XFILLER_6_115 vgnd vpwr scs8hd_decap_8
X_151_ address[0] _150_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_122 vgnd vpwr scs8hd_decap_6
XFILLER_10_177 vgnd vpwr scs8hd_decap_12
X_082_ address[2] _133_/B vgnd vpwr scs8hd_inv_8
XFILLER_37_92 vpwr vgnd scs8hd_fill_2
XFILLER_37_70 vpwr vgnd scs8hd_fill_2
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _087_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
X_203_ _203_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_134_ _153_/A _135_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_162 vpwr vgnd scs8hd_fill_2
XFILLER_17_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vgnd vpwr scs8hd_decap_8
XFILLER_12_239 vgnd vpwr scs8hd_decap_8
XFILLER_34_93 vpwr vgnd scs8hd_fill_2
X_117_ _117_/A _117_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_158 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_18 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _112_/A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_40 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vgnd vpwr scs8hd_fill_1
XFILLER_29_71 vgnd vpwr scs8hd_decap_3
XFILLER_28_180 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_1_.latch data_in _119_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_17_117 vpwr vgnd scs8hd_fill_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_161 vpwr vgnd scs8hd_fill_2
XFILLER_15_95 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_14_109 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_197 vgnd vpwr scs8hd_decap_12
XFILLER_13_175 vgnd vpwr scs8hd_decap_8
XFILLER_3_10 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _113_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
X_150_ _153_/A _150_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_149 vgnd vpwr scs8hd_decap_4
XFILLER_10_145 vgnd vpwr scs8hd_decap_8
XFILLER_10_189 vgnd vpwr scs8hd_decap_12
X_081_ address[3] _145_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_204 vgnd vpwr scs8hd_decap_8
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _106_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
X_133_ address[3] _133_/B _133_/C _133_/D _135_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
XFILLER_23_84 vgnd vpwr scs8hd_decap_8
X_202_ _202_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _099_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _120_/A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _085_/A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
XFILLER_7_266 vgnd vpwr scs8hd_decap_8
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XFILLER_11_262 vgnd vpwr scs8hd_decap_12
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _116_/A _116_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_148 vgnd vpwr scs8hd_decap_4
XFILLER_29_137 vpwr vgnd scs8hd_fill_2
XFILLER_37_192 vgnd vpwr scs8hd_decap_12
XFILLER_37_181 vpwr vgnd scs8hd_fill_2
XFILLER_4_258 vgnd vpwr scs8hd_decap_12
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_28_192 vgnd vpwr scs8hd_decap_12
XFILLER_6_65 vgnd vpwr scs8hd_decap_8
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _090_/Y mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_34_140 vgnd vpwr scs8hd_decap_8
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch data_in _104_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_0_.latch data_in _094_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_40_121 vgnd vpwr scs8hd_decap_12
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_25_140 vgnd vpwr scs8hd_decap_6
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_132 vgnd vpwr scs8hd_decap_6
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_36_18 vgnd vpwr scs8hd_decap_12
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _108_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _101_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _086_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_147 vgnd vpwr scs8hd_decap_6
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_3_22 vgnd vpwr scs8hd_decap_12
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_99 vpwr vgnd scs8hd_fill_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ address[5] _173_/D vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_50 vgnd vpwr scs8hd_decap_8
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_132_ address[0] _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
X_201_ _201_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_23_30 vgnd vpwr scs8hd_decap_4
XFILLER_2_120 vgnd vpwr scs8hd_decap_12
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _196_/A vgnd vpwr scs8hd_inv_1
XFILLER_9_10 vgnd vpwr scs8hd_decap_12
XFILLER_14_271 vgnd vpwr scs8hd_decap_4
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _107_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XANTENNA__211__A _211_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_40 vgnd vpwr scs8hd_fill_1
XFILLER_7_201 vgnd vpwr scs8hd_decap_12
XFILLER_7_245 vpwr vgnd scs8hd_fill_2
XFILLER_11_274 vgnd vpwr scs8hd_decap_3
X_115_ _115_/A _115_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_116 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _087_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_64 vgnd vpwr scs8hd_decap_3
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vgnd vpwr scs8hd_decap_4
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_26_108 vpwr vgnd scs8hd_fill_2
XFILLER_34_163 vgnd vpwr scs8hd_decap_8
XFILLER_34_152 vgnd vpwr scs8hd_fill_1
XFILLER_19_160 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _186_/HI _111_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_133 vgnd vpwr scs8hd_decap_12
XFILLER_15_86 vgnd vpwr scs8hd_decap_6
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_96 vgnd vpwr scs8hd_fill_1
XFILLER_31_52 vpwr vgnd scs8hd_fill_2
XFILLER_0_262 vgnd vpwr scs8hd_decap_12
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XFILLER_16_174 vgnd vpwr scs8hd_decap_12
XFILLER_31_155 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

